netcdf ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-1.clm2.h0.0001-01-02-00000 {
dimensions:
	lndgrid = 338 ;
	gridcell = 338 ;
	landunit = 1352 ;
	column = 5408 ;
	pft = 10816 ;
	levgrnd = 15 ;
	levurb = 5 ;
	levlak = 10 ;
	numrad = 2 ;
	string_length = 8 ;
	levdcmp = 15 ;
	hist_interval = 2 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float levgrnd(levgrnd) ;
		levgrnd:long_name = "coordinate soil levels" ;
		levgrnd:units = "m" ;
	float levlak(levlak) ;
		levlak:long_name = "coordinate lake levels" ;
		levlak:units = "m" ;
	float levdcmp(levdcmp) ;
		levdcmp:long_name = "coordinate soil levels" ;
		levdcmp:units = "m" ;
	float time(time) ;
		time:long_name = "time" ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bounds" ;
	int mcdate(time) ;
		mcdate:long_name = "current date (YYYYMMDD)" ;
	int mcsec(time) ;
		mcsec:long_name = "current seconds of current date" ;
		mcsec:units = "s" ;
	int mdcur(time) ;
		mdcur:long_name = "current day (from base day)" ;
	int mscur(time) ;
		mscur:long_name = "current seconds of current day" ;
	int nstep(time) ;
		nstep:long_name = "time step" ;
	double time_bounds(time, hist_interval) ;
		time_bounds:long_name = "history time interval endpoints" ;
	char date_written(time, string_length) ;
	char time_written(time, string_length) ;
	float lon(lndgrid) ;
		lon:long_name = "coordinate longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = 1.e+36f ;
		lon:missing_value = 1.e+36f ;
	float lat(lndgrid) ;
		lat:long_name = "coordinate latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = 1.e+36f ;
		lat:missing_value = 1.e+36f ;
	float area(lndgrid) ;
		area:long_name = "grid cell areas" ;
		area:units = "km^2" ;
		area:_FillValue = 1.e+36f ;
		area:missing_value = 1.e+36f ;
	float topo(lndgrid) ;
		topo:long_name = "grid cell topography" ;
		topo:units = "m" ;
		topo:_FillValue = 1.e+36f ;
		topo:missing_value = 1.e+36f ;
	float landfrac(lndgrid) ;
		landfrac:long_name = "land fraction" ;
		landfrac:_FillValue = 1.e+36f ;
		landfrac:missing_value = 1.e+36f ;
	int landmask(lndgrid) ;
		landmask:long_name = "land/ocean mask (0.=ocean and 1.=land)" ;
		landmask:_FillValue = -9999 ;
		landmask:missing_value = -9999 ;
	int pftmask(lndgrid) ;
		pftmask:long_name = "pft real/fake mask (0.=fake and 1.=real)" ;
		pftmask:_FillValue = -9999 ;
		pftmask:missing_value = -9999 ;
	float ACTUAL_IMMOB(time, lndgrid) ;
		ACTUAL_IMMOB:long_name = "actual N immobilization" ;
		ACTUAL_IMMOB:units = "gN/m^2/s" ;
		ACTUAL_IMMOB:cell_methods = "time: mean" ;
		ACTUAL_IMMOB:_FillValue = 1.e+36f ;
		ACTUAL_IMMOB:missing_value = 1.e+36f ;
	float AGNPP(time, lndgrid) ;
		AGNPP:long_name = "aboveground NPP" ;
		AGNPP:units = "gC/m^2/s" ;
		AGNPP:cell_methods = "time: mean" ;
		AGNPP:_FillValue = 1.e+36f ;
		AGNPP:missing_value = 1.e+36f ;
	float ALT(time, lndgrid) ;
		ALT:long_name = "current active layer thickness" ;
		ALT:units = "m" ;
		ALT:cell_methods = "time: mean" ;
		ALT:_FillValue = 1.e+36f ;
		ALT:missing_value = 1.e+36f ;
	float ALTMAX(time, lndgrid) ;
		ALTMAX:long_name = "maximum annual active layer thickness" ;
		ALTMAX:units = "m" ;
		ALTMAX:cell_methods = "time: mean" ;
		ALTMAX:_FillValue = 1.e+36f ;
		ALTMAX:missing_value = 1.e+36f ;
	float ALTMAX_LASTYEAR(time, lndgrid) ;
		ALTMAX_LASTYEAR:long_name = "maximum prior year active layer thickness" ;
		ALTMAX_LASTYEAR:units = "m" ;
		ALTMAX_LASTYEAR:cell_methods = "time: mean" ;
		ALTMAX_LASTYEAR:_FillValue = 1.e+36f ;
		ALTMAX_LASTYEAR:missing_value = 1.e+36f ;
	float AR(time, lndgrid) ;
		AR:long_name = "autotrophic respiration (MR + GR)" ;
		AR:units = "gC/m^2/s" ;
		AR:cell_methods = "time: mean" ;
		AR:_FillValue = 1.e+36f ;
		AR:missing_value = 1.e+36f ;
	float BAF_CROP(time, lndgrid) ;
		BAF_CROP:long_name = "timestep fractional area burned for crop" ;
		BAF_CROP:units = "proportion" ;
		BAF_CROP:cell_methods = "time: mean" ;
		BAF_CROP:_FillValue = 1.e+36f ;
		BAF_CROP:missing_value = 1.e+36f ;
	float BAF_PEATF(time, lndgrid) ;
		BAF_PEATF:long_name = "timestep fractional area burned in peatland" ;
		BAF_PEATF:units = "proportion" ;
		BAF_PEATF:cell_methods = "time: mean" ;
		BAF_PEATF:_FillValue = 1.e+36f ;
		BAF_PEATF:missing_value = 1.e+36f ;
	float BCDEP(time, lndgrid) ;
		BCDEP:long_name = "total BC deposition (dry+wet) from atmosphere" ;
		BCDEP:units = "kg/m^2/s" ;
		BCDEP:cell_methods = "time: mean" ;
		BCDEP:_FillValue = 1.e+36f ;
		BCDEP:missing_value = 1.e+36f ;
	float BGNPP(time, lndgrid) ;
		BGNPP:long_name = "belowground NPP" ;
		BGNPP:units = "gC/m^2/s" ;
		BGNPP:cell_methods = "time: mean" ;
		BGNPP:_FillValue = 1.e+36f ;
		BGNPP:missing_value = 1.e+36f ;
	float BTRAN(time, lndgrid) ;
		BTRAN:long_name = "transpiration beta factor" ;
		BTRAN:units = "unitless" ;
		BTRAN:cell_methods = "time: mean" ;
		BTRAN:_FillValue = 1.e+36f ;
		BTRAN:missing_value = 1.e+36f ;
	float BUILDHEAT(time, lndgrid) ;
		BUILDHEAT:long_name = "heat flux from urban building interior to walls and roof" ;
		BUILDHEAT:units = "W/m^2" ;
		BUILDHEAT:cell_methods = "time: mean" ;
		BUILDHEAT:_FillValue = 1.e+36f ;
		BUILDHEAT:missing_value = 1.e+36f ;
	float CH4PROD(time, lndgrid) ;
		CH4PROD:long_name = "Gridcell total production of CH4" ;
		CH4PROD:units = "gC/m2/s" ;
		CH4PROD:cell_methods = "time: mean" ;
		CH4PROD:_FillValue = 1.e+36f ;
		CH4PROD:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_SAT(time, lndgrid) ;
		CH4_SURF_AERE_SAT:long_name = "aerenchyma surface CH4 flux for inundated area; (+ to atm)" ;
		CH4_SURF_AERE_SAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_SAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_UNSAT(time, lndgrid) ;
		CH4_SURF_AERE_UNSAT:long_name = "aerenchyma surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_AERE_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_SAT(time, lndgrid) ;
		CH4_SURF_DIFF_SAT:long_name = "diffusive surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_DIFF_SAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_SAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_UNSAT(time, lndgrid) ;
		CH4_SURF_DIFF_UNSAT:long_name = "diffusive surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_DIFF_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_SAT(time, lndgrid) ;
		CH4_SURF_EBUL_SAT:long_name = "ebullition surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_EBUL_SAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_SAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_UNSAT(time, lndgrid) ;
		CH4_SURF_EBUL_UNSAT:long_name = "ebullition surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_EBUL_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_UNSAT:missing_value = 1.e+36f ;
	float COL_CTRUNC(time, lndgrid) ;
		COL_CTRUNC:long_name = "column-level sink for C truncation" ;
		COL_CTRUNC:units = "gC/m^2" ;
		COL_CTRUNC:cell_methods = "time: mean" ;
		COL_CTRUNC:_FillValue = 1.e+36f ;
		COL_CTRUNC:missing_value = 1.e+36f ;
	float COL_FIRE_CLOSS(time, lndgrid) ;
		COL_FIRE_CLOSS:long_name = "total column-level fire C loss for non-peat fires outside land-type converted region" ;
		COL_FIRE_CLOSS:units = "gC/m^2/s" ;
		COL_FIRE_CLOSS:cell_methods = "time: mean" ;
		COL_FIRE_CLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_CLOSS:missing_value = 1.e+36f ;
	float COL_FIRE_NLOSS(time, lndgrid) ;
		COL_FIRE_NLOSS:long_name = "total column-level fire N loss" ;
		COL_FIRE_NLOSS:units = "gN/m^2/s" ;
		COL_FIRE_NLOSS:cell_methods = "time: mean" ;
		COL_FIRE_NLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_NLOSS:missing_value = 1.e+36f ;
	float COL_NTRUNC(time, lndgrid) ;
		COL_NTRUNC:long_name = "column-level sink for N truncation" ;
		COL_NTRUNC:units = "gN/m^2" ;
		COL_NTRUNC:cell_methods = "time: mean" ;
		COL_NTRUNC:_FillValue = 1.e+36f ;
		COL_NTRUNC:missing_value = 1.e+36f ;
	float CONC_CH4_SAT(time, levgrnd, lndgrid) ;
		CONC_CH4_SAT:long_name = "CH4 soil Concentration for inundated / lake area" ;
		CONC_CH4_SAT:units = "mol/m3" ;
		CONC_CH4_SAT:cell_methods = "time: mean" ;
		CONC_CH4_SAT:_FillValue = 1.e+36f ;
		CONC_CH4_SAT:missing_value = 1.e+36f ;
	float CONC_CH4_UNSAT(time, levgrnd, lndgrid) ;
		CONC_CH4_UNSAT:long_name = "CH4 soil Concentration for non-inundated area" ;
		CONC_CH4_UNSAT:units = "mol/m3" ;
		CONC_CH4_UNSAT:cell_methods = "time: mean" ;
		CONC_CH4_UNSAT:_FillValue = 1.e+36f ;
		CONC_CH4_UNSAT:missing_value = 1.e+36f ;
	float CONC_O2_SAT(time, levgrnd, lndgrid) ;
		CONC_O2_SAT:long_name = "O2 soil Concentration for inundated / lake area" ;
		CONC_O2_SAT:units = "mol/m3" ;
		CONC_O2_SAT:cell_methods = "time: mean" ;
		CONC_O2_SAT:_FillValue = 1.e+36f ;
		CONC_O2_SAT:missing_value = 1.e+36f ;
	float CONC_O2_UNSAT(time, levgrnd, lndgrid) ;
		CONC_O2_UNSAT:long_name = "O2 soil Concentration for non-inundated area" ;
		CONC_O2_UNSAT:units = "mol/m3" ;
		CONC_O2_UNSAT:cell_methods = "time: mean" ;
		CONC_O2_UNSAT:_FillValue = 1.e+36f ;
		CONC_O2_UNSAT:missing_value = 1.e+36f ;
	float CPOOL(time, lndgrid) ;
		CPOOL:long_name = "temporary photosynthate C pool" ;
		CPOOL:units = "gC/m^2" ;
		CPOOL:cell_methods = "time: mean" ;
		CPOOL:_FillValue = 1.e+36f ;
		CPOOL:missing_value = 1.e+36f ;
	float CWDC(time, lndgrid) ;
		CWDC:long_name = "CWD C" ;
		CWDC:units = "gC/m^2" ;
		CWDC:cell_methods = "time: mean" ;
		CWDC:_FillValue = 1.e+36f ;
		CWDC:missing_value = 1.e+36f ;
	float CWDC_HR(time, lndgrid) ;
		CWDC_HR:long_name = "coarse woody debris C heterotrophic respiration" ;
		CWDC_HR:units = "gC/m^2/s" ;
		CWDC_HR:cell_methods = "time: mean" ;
		CWDC_HR:_FillValue = 1.e+36f ;
		CWDC_HR:missing_value = 1.e+36f ;
	float CWDC_LOSS(time, lndgrid) ;
		CWDC_LOSS:long_name = "coarse woody debris C loss" ;
		CWDC_LOSS:units = "gC/m^2/s" ;
		CWDC_LOSS:cell_methods = "time: mean" ;
		CWDC_LOSS:_FillValue = 1.e+36f ;
		CWDC_LOSS:missing_value = 1.e+36f ;
	float CWDC_TO_LITR2C(time, lndgrid) ;
		CWDC_TO_LITR2C:long_name = "decomp. of coarse woody debris C to litter 2 C" ;
		CWDC_TO_LITR2C:units = "gC/m^2/s" ;
		CWDC_TO_LITR2C:cell_methods = "time: mean" ;
		CWDC_TO_LITR2C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR2C:missing_value = 1.e+36f ;
	float CWDC_TO_LITR3C(time, lndgrid) ;
		CWDC_TO_LITR3C:long_name = "decomp. of coarse woody debris C to litter 3 C" ;
		CWDC_TO_LITR3C:units = "gC/m^2/s" ;
		CWDC_TO_LITR3C:cell_methods = "time: mean" ;
		CWDC_TO_LITR3C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR3C:missing_value = 1.e+36f ;
	float CWDC_vr(time, levdcmp, lndgrid) ;
		CWDC_vr:long_name = "CWD C (vertically resolved)" ;
		CWDC_vr:units = "gC/m^3" ;
		CWDC_vr:cell_methods = "time: mean" ;
		CWDC_vr:_FillValue = 1.e+36f ;
		CWDC_vr:missing_value = 1.e+36f ;
	float CWDN(time, lndgrid) ;
		CWDN:long_name = "CWD N" ;
		CWDN:units = "gN/m^2" ;
		CWDN:cell_methods = "time: mean" ;
		CWDN:_FillValue = 1.e+36f ;
		CWDN:missing_value = 1.e+36f ;
	float CWDN_TO_LITR2N(time, lndgrid) ;
		CWDN_TO_LITR2N:long_name = "decomp. of coarse woody debris N to litter 2 N" ;
		CWDN_TO_LITR2N:units = "gN/m^2" ;
		CWDN_TO_LITR2N:cell_methods = "time: mean" ;
		CWDN_TO_LITR2N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR2N:missing_value = 1.e+36f ;
	float CWDN_TO_LITR3N(time, lndgrid) ;
		CWDN_TO_LITR3N:long_name = "decomp. of coarse woody debris N to litter 3 N" ;
		CWDN_TO_LITR3N:units = "gN/m^2" ;
		CWDN_TO_LITR3N:cell_methods = "time: mean" ;
		CWDN_TO_LITR3N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR3N:missing_value = 1.e+36f ;
	float CWDN_vr(time, levdcmp, lndgrid) ;
		CWDN_vr:long_name = "CWD N (vertically resolved)" ;
		CWDN_vr:units = "gN/m^3" ;
		CWDN_vr:cell_methods = "time: mean" ;
		CWDN_vr:_FillValue = 1.e+36f ;
		CWDN_vr:missing_value = 1.e+36f ;
	float DEADCROOTC(time, lndgrid) ;
		DEADCROOTC:long_name = "dead coarse root C" ;
		DEADCROOTC:units = "gC/m^2" ;
		DEADCROOTC:cell_methods = "time: mean" ;
		DEADCROOTC:_FillValue = 1.e+36f ;
		DEADCROOTC:missing_value = 1.e+36f ;
	float DEADCROOTN(time, lndgrid) ;
		DEADCROOTN:long_name = "dead coarse root N" ;
		DEADCROOTN:units = "gN/m^2" ;
		DEADCROOTN:cell_methods = "time: mean" ;
		DEADCROOTN:_FillValue = 1.e+36f ;
		DEADCROOTN:missing_value = 1.e+36f ;
	float DEADSTEMC(time, lndgrid) ;
		DEADSTEMC:long_name = "dead stem C" ;
		DEADSTEMC:units = "gC/m^2" ;
		DEADSTEMC:cell_methods = "time: mean" ;
		DEADSTEMC:_FillValue = 1.e+36f ;
		DEADSTEMC:missing_value = 1.e+36f ;
	float DEADSTEMN(time, lndgrid) ;
		DEADSTEMN:long_name = "dead stem N" ;
		DEADSTEMN:units = "gN/m^2" ;
		DEADSTEMN:cell_methods = "time: mean" ;
		DEADSTEMN:_FillValue = 1.e+36f ;
		DEADSTEMN:missing_value = 1.e+36f ;
	float DENIT(time, lndgrid) ;
		DENIT:long_name = "total rate of denitrification" ;
		DENIT:units = "gN/m^2/s" ;
		DENIT:cell_methods = "time: mean" ;
		DENIT:_FillValue = 1.e+36f ;
		DENIT:missing_value = 1.e+36f ;
	float DISPVEGC(time, lndgrid) ;
		DISPVEGC:long_name = "displayed veg carbon, excluding storage and cpool" ;
		DISPVEGC:units = "gC/m^2" ;
		DISPVEGC:cell_methods = "time: mean" ;
		DISPVEGC:_FillValue = 1.e+36f ;
		DISPVEGC:missing_value = 1.e+36f ;
	float DISPVEGN(time, lndgrid) ;
		DISPVEGN:long_name = "displayed vegetation nitrogen" ;
		DISPVEGN:units = "gN/m^2" ;
		DISPVEGN:cell_methods = "time: mean" ;
		DISPVEGN:_FillValue = 1.e+36f ;
		DISPVEGN:missing_value = 1.e+36f ;
	float DSTDEP(time, lndgrid) ;
		DSTDEP:long_name = "total dust deposition (dry+wet) from atmosphere" ;
		DSTDEP:units = "kg/m^2/s" ;
		DSTDEP:cell_methods = "time: mean" ;
		DSTDEP:_FillValue = 1.e+36f ;
		DSTDEP:missing_value = 1.e+36f ;
	float DSTFLXT(time, lndgrid) ;
		DSTFLXT:long_name = "total surface dust emission" ;
		DSTFLXT:units = "kg/m2/s" ;
		DSTFLXT:cell_methods = "time: mean" ;
		DSTFLXT:_FillValue = 1.e+36f ;
		DSTFLXT:missing_value = 1.e+36f ;
	float DWT_CLOSS(time, lndgrid) ;
		DWT_CLOSS:long_name = "total carbon loss from land cover conversion" ;
		DWT_CLOSS:units = "gC/m^2/s" ;
		DWT_CLOSS:cell_methods = "time: mean" ;
		DWT_CLOSS:_FillValue = 1.e+36f ;
		DWT_CLOSS:missing_value = 1.e+36f ;
	float DWT_CONV_CFLUX(time, lndgrid) ;
		DWT_CONV_CFLUX:long_name = "conversion C flux (immediate loss to atm)" ;
		DWT_CONV_CFLUX:units = "gC/m^2/s" ;
		DWT_CONV_CFLUX:cell_methods = "time: mean" ;
		DWT_CONV_CFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_CFLUX:missing_value = 1.e+36f ;
	float DWT_CONV_NFLUX(time, lndgrid) ;
		DWT_CONV_NFLUX:long_name = "conversion N flux (immediate loss to atm)" ;
		DWT_CONV_NFLUX:units = "gN/m^2/s" ;
		DWT_CONV_NFLUX:cell_methods = "time: mean" ;
		DWT_CONV_NFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_NFLUX:missing_value = 1.e+36f ;
	float DWT_NLOSS(time, lndgrid) ;
		DWT_NLOSS:long_name = "total nitrogen loss from landcover conversion" ;
		DWT_NLOSS:units = "gN/m^2/s" ;
		DWT_NLOSS:cell_methods = "time: mean" ;
		DWT_NLOSS:_FillValue = 1.e+36f ;
		DWT_NLOSS:missing_value = 1.e+36f ;
	float DWT_PROD100C_GAIN(time, lndgrid) ;
		DWT_PROD100C_GAIN:long_name = "landcover change-driven addition to 100-yr wood product pool" ;
		DWT_PROD100C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD100C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD100N_GAIN(time, lndgrid) ;
		DWT_PROD100N_GAIN:long_name = "addition to 100-yr wood product pool" ;
		DWT_PROD100N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD100N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100N_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10C_GAIN(time, lndgrid) ;
		DWT_PROD10C_GAIN:long_name = "landcover change-driven addition to 10-yr wood product pool" ;
		DWT_PROD10C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD10C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10N_GAIN(time, lndgrid) ;
		DWT_PROD10N_GAIN:long_name = "addition to 10-yr wood product pool" ;
		DWT_PROD10N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD10N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10N_GAIN:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDC_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDC_TO_DEADSTEM:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_LEAF(time, lndgrid) ;
		DWT_SEEDC_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDC_TO_LEAF:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_LEAF:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDN_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDN_TO_DEADSTEM:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_LEAF(time, lndgrid) ;
		DWT_SEEDN_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDN_TO_LEAF:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_LEAF:missing_value = 1.e+36f ;
	float EFLX_DYNBAL(time, lndgrid) ;
		EFLX_DYNBAL:long_name = "dynamic land cover change conversion energy flux" ;
		EFLX_DYNBAL:units = "W/m^2" ;
		EFLX_DYNBAL:cell_methods = "time: mean" ;
		EFLX_DYNBAL:_FillValue = 1.e+36f ;
		EFLX_DYNBAL:missing_value = 1.e+36f ;
	float EFLX_GRND_LAKE(time, lndgrid) ;
		EFLX_GRND_LAKE:long_name = "net heat flux into lake/snow surface, excluding light transmission" ;
		EFLX_GRND_LAKE:units = "W/m^2" ;
		EFLX_GRND_LAKE:cell_methods = "time: mean" ;
		EFLX_GRND_LAKE:_FillValue = 1.e+36f ;
		EFLX_GRND_LAKE:missing_value = 1.e+36f ;
	float EFLX_LH_TOT(time, lndgrid) ;
		EFLX_LH_TOT:long_name = "total latent heat flux [+ to atm]" ;
		EFLX_LH_TOT:units = "W/m^2" ;
		EFLX_LH_TOT:cell_methods = "time: mean" ;
		EFLX_LH_TOT:_FillValue = 1.e+36f ;
		EFLX_LH_TOT:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_R(time, lndgrid) ;
		EFLX_LH_TOT_R:long_name = "Rural total evaporation" ;
		EFLX_LH_TOT_R:units = "W/m^2" ;
		EFLX_LH_TOT_R:cell_methods = "time: mean" ;
		EFLX_LH_TOT_R:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_R:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_U(time, lndgrid) ;
		EFLX_LH_TOT_U:long_name = "Urban total evaporation" ;
		EFLX_LH_TOT_U:units = "W/m^2" ;
		EFLX_LH_TOT_U:cell_methods = "time: mean" ;
		EFLX_LH_TOT_U:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_U:missing_value = 1.e+36f ;
	float ELAI(time, lndgrid) ;
		ELAI:long_name = "exposed one-sided leaf area index" ;
		ELAI:units = "m^2/m^2" ;
		ELAI:cell_methods = "time: mean" ;
		ELAI:_FillValue = 1.e+36f ;
		ELAI:missing_value = 1.e+36f ;
	float ER(time, lndgrid) ;
		ER:long_name = "total ecosystem respiration, autotrophic + heterotrophic" ;
		ER:units = "gC/m^2/s" ;
		ER:cell_methods = "time: mean" ;
		ER:_FillValue = 1.e+36f ;
		ER:missing_value = 1.e+36f ;
	float ERRH2O(time, lndgrid) ;
		ERRH2O:long_name = "total water conservation error" ;
		ERRH2O:units = "mm" ;
		ERRH2O:cell_methods = "time: mean" ;
		ERRH2O:_FillValue = 1.e+36f ;
		ERRH2O:missing_value = 1.e+36f ;
	float ERRH2OSNO(time, lndgrid) ;
		ERRH2OSNO:long_name = "imbalance in snow depth (liquid water)" ;
		ERRH2OSNO:units = "mm" ;
		ERRH2OSNO:cell_methods = "time: mean" ;
		ERRH2OSNO:_FillValue = 1.e+36f ;
		ERRH2OSNO:missing_value = 1.e+36f ;
	float ERRSEB(time, lndgrid) ;
		ERRSEB:long_name = "surface energy conservation error" ;
		ERRSEB:units = "W/m^2" ;
		ERRSEB:cell_methods = "time: mean" ;
		ERRSEB:_FillValue = 1.e+36f ;
		ERRSEB:missing_value = 1.e+36f ;
	float ERRSOI(time, lndgrid) ;
		ERRSOI:long_name = "soil/lake energy conservation error" ;
		ERRSOI:units = "W/m^2" ;
		ERRSOI:cell_methods = "time: mean" ;
		ERRSOI:_FillValue = 1.e+36f ;
		ERRSOI:missing_value = 1.e+36f ;
	float ERRSOL(time, lndgrid) ;
		ERRSOL:long_name = "solar radiation conservation error" ;
		ERRSOL:units = "W/m^2" ;
		ERRSOL:cell_methods = "time: mean" ;
		ERRSOL:_FillValue = 1.e+36f ;
		ERRSOL:missing_value = 1.e+36f ;
	float ESAI(time, lndgrid) ;
		ESAI:long_name = "exposed one-sided stem area index" ;
		ESAI:units = "m^2/m^2" ;
		ESAI:cell_methods = "time: mean" ;
		ESAI:_FillValue = 1.e+36f ;
		ESAI:missing_value = 1.e+36f ;
	float FAREA_BURNED(time, lndgrid) ;
		FAREA_BURNED:long_name = "timestep fractional area burned" ;
		FAREA_BURNED:units = "proportion" ;
		FAREA_BURNED:cell_methods = "time: mean" ;
		FAREA_BURNED:_FillValue = 1.e+36f ;
		FAREA_BURNED:missing_value = 1.e+36f ;
	float FCEV(time, lndgrid) ;
		FCEV:long_name = "canopy evaporation" ;
		FCEV:units = "W/m^2" ;
		FCEV:cell_methods = "time: mean" ;
		FCEV:_FillValue = 1.e+36f ;
		FCEV:missing_value = 1.e+36f ;
	float FCH4(time, lndgrid) ;
		FCH4:long_name = "Gridcell surface CH4 flux to atmosphere (+ to atm)" ;
		FCH4:units = "kgC/m2/s" ;
		FCH4:cell_methods = "time: mean" ;
		FCH4:_FillValue = 1.e+36f ;
		FCH4:missing_value = 1.e+36f ;
	float FCH4TOCO2(time, lndgrid) ;
		FCH4TOCO2:long_name = "Gridcell oxidation of CH4 to CO2" ;
		FCH4TOCO2:units = "gC/m2/s" ;
		FCH4TOCO2:cell_methods = "time: mean" ;
		FCH4TOCO2:_FillValue = 1.e+36f ;
		FCH4TOCO2:missing_value = 1.e+36f ;
	float FCH4_DFSAT(time, lndgrid) ;
		FCH4_DFSAT:long_name = "CH4 additional flux due to changing fsat, vegetated landunits only" ;
		FCH4_DFSAT:units = "kgC/m2/s" ;
		FCH4_DFSAT:cell_methods = "time: mean" ;
		FCH4_DFSAT:_FillValue = 1.e+36f ;
		FCH4_DFSAT:missing_value = 1.e+36f ;
	float FCOV(time, lndgrid) ;
		FCOV:long_name = "fractional impermeable area" ;
		FCOV:units = "unitless" ;
		FCOV:cell_methods = "time: mean" ;
		FCOV:_FillValue = 1.e+36f ;
		FCOV:missing_value = 1.e+36f ;
	float FCTR(time, lndgrid) ;
		FCTR:long_name = "canopy transpiration" ;
		FCTR:units = "W/m^2" ;
		FCTR:cell_methods = "time: mean" ;
		FCTR:_FillValue = 1.e+36f ;
		FCTR:missing_value = 1.e+36f ;
	float FGEV(time, lndgrid) ;
		FGEV:long_name = "ground evaporation" ;
		FGEV:units = "W/m^2" ;
		FGEV:cell_methods = "time: mean" ;
		FGEV:_FillValue = 1.e+36f ;
		FGEV:missing_value = 1.e+36f ;
	float FGR(time, lndgrid) ;
		FGR:long_name = "heat flux into soil/snow including snow melt and lake / snow light transmission" ;
		FGR:units = "W/m^2" ;
		FGR:cell_methods = "time: mean" ;
		FGR:_FillValue = 1.e+36f ;
		FGR:missing_value = 1.e+36f ;
	float FGR12(time, lndgrid) ;
		FGR12:long_name = "heat flux between soil layers 1 and 2" ;
		FGR12:units = "W/m^2" ;
		FGR12:cell_methods = "time: mean" ;
		FGR12:_FillValue = 1.e+36f ;
		FGR12:missing_value = 1.e+36f ;
	float FGR_R(time, lndgrid) ;
		FGR_R:long_name = "Rural heat flux into soil/snow including snow melt and snow light transmission" ;
		FGR_R:units = "W/m^2" ;
		FGR_R:cell_methods = "time: mean" ;
		FGR_R:_FillValue = 1.e+36f ;
		FGR_R:missing_value = 1.e+36f ;
	float FGR_U(time, lndgrid) ;
		FGR_U:long_name = "Urban heat flux into soil/snow including snow melt" ;
		FGR_U:units = "W/m^2" ;
		FGR_U:cell_methods = "time: mean" ;
		FGR_U:_FillValue = 1.e+36f ;
		FGR_U:missing_value = 1.e+36f ;
	float FH2OSFC(time, lndgrid) ;
		FH2OSFC:long_name = "fraction of ground covered by surface water" ;
		FH2OSFC:units = "unitless" ;
		FH2OSFC:cell_methods = "time: mean" ;
		FH2OSFC:_FillValue = 1.e+36f ;
		FH2OSFC:missing_value = 1.e+36f ;
	float FINUNDATED(time, lndgrid) ;
		FINUNDATED:long_name = "fractional inundated area of vegetated columns" ;
		FINUNDATED:units = "unitless" ;
		FINUNDATED:cell_methods = "time: mean" ;
		FINUNDATED:_FillValue = 1.e+36f ;
		FINUNDATED:missing_value = 1.e+36f ;
	float FINUNDATED_LAG(time, lndgrid) ;
		FINUNDATED_LAG:long_name = "time-lagged inundated fraction of vegetated columns" ;
		FINUNDATED_LAG:units = "unitless" ;
		FINUNDATED_LAG:cell_methods = "time: mean" ;
		FINUNDATED_LAG:_FillValue = 1.e+36f ;
		FINUNDATED_LAG:missing_value = 1.e+36f ;
	float FIRA(time, lndgrid) ;
		FIRA:long_name = "net infrared (longwave) radiation" ;
		FIRA:units = "W/m^2" ;
		FIRA:cell_methods = "time: mean" ;
		FIRA:_FillValue = 1.e+36f ;
		FIRA:missing_value = 1.e+36f ;
	float FIRA_R(time, lndgrid) ;
		FIRA_R:long_name = "Rural net infrared (longwave) radiation" ;
		FIRA_R:units = "W/m^2" ;
		FIRA_R:cell_methods = "time: mean" ;
		FIRA_R:_FillValue = 1.e+36f ;
		FIRA_R:missing_value = 1.e+36f ;
	float FIRA_U(time, lndgrid) ;
		FIRA_U:long_name = "Urban net infrared (longwave) radiation" ;
		FIRA_U:units = "W/m^2" ;
		FIRA_U:cell_methods = "time: mean" ;
		FIRA_U:_FillValue = 1.e+36f ;
		FIRA_U:missing_value = 1.e+36f ;
	float FIRE(time, lndgrid) ;
		FIRE:long_name = "emitted infrared (longwave) radiation" ;
		FIRE:units = "W/m^2" ;
		FIRE:cell_methods = "time: mean" ;
		FIRE:_FillValue = 1.e+36f ;
		FIRE:missing_value = 1.e+36f ;
	float FIRE_R(time, lndgrid) ;
		FIRE_R:long_name = "Rural emitted infrared (longwave) radiation" ;
		FIRE_R:units = "W/m^2" ;
		FIRE_R:cell_methods = "time: mean" ;
		FIRE_R:_FillValue = 1.e+36f ;
		FIRE_R:missing_value = 1.e+36f ;
	float FIRE_U(time, lndgrid) ;
		FIRE_U:long_name = "Urban emitted infrared (longwave) radiation" ;
		FIRE_U:units = "W/m^2" ;
		FIRE_U:cell_methods = "time: mean" ;
		FIRE_U:_FillValue = 1.e+36f ;
		FIRE_U:missing_value = 1.e+36f ;
	float FLDS(time, lndgrid) ;
		FLDS:long_name = "atmospheric longwave radiation" ;
		FLDS:units = "W/m^2" ;
		FLDS:cell_methods = "time: mean" ;
		FLDS:_FillValue = 1.e+36f ;
		FLDS:missing_value = 1.e+36f ;
	float FPG(time, lndgrid) ;
		FPG:long_name = "fraction of potential gpp" ;
		FPG:units = "proportion" ;
		FPG:cell_methods = "time: mean" ;
		FPG:_FillValue = 1.e+36f ;
		FPG:missing_value = 1.e+36f ;
	float FPI(time, lndgrid) ;
		FPI:long_name = "fraction of potential immobilization" ;
		FPI:units = "proportion" ;
		FPI:cell_methods = "time: mean" ;
		FPI:_FillValue = 1.e+36f ;
		FPI:missing_value = 1.e+36f ;
	float FPI_vr(time, levdcmp, lndgrid) ;
		FPI_vr:long_name = "fraction of potential immobilization" ;
		FPI_vr:units = "proportion" ;
		FPI_vr:cell_methods = "time: mean" ;
		FPI_vr:_FillValue = 1.e+36f ;
		FPI_vr:missing_value = 1.e+36f ;
	float FPSN(time, lndgrid) ;
		FPSN:long_name = "photosynthesis" ;
		FPSN:units = "umol/m2s" ;
		FPSN:cell_methods = "time: mean" ;
		FPSN:_FillValue = 1.e+36f ;
		FPSN:missing_value = 1.e+36f ;
	float FPSN_WC(time, lndgrid) ;
		FPSN_WC:long_name = "Rubisco-limited photosynthesis" ;
		FPSN_WC:units = "umol/m2s" ;
		FPSN_WC:cell_methods = "time: mean" ;
		FPSN_WC:_FillValue = 1.e+36f ;
		FPSN_WC:missing_value = 1.e+36f ;
	float FPSN_WJ(time, lndgrid) ;
		FPSN_WJ:long_name = "RuBP-limited photosynthesis" ;
		FPSN_WJ:units = "umol/m2s" ;
		FPSN_WJ:cell_methods = "time: mean" ;
		FPSN_WJ:_FillValue = 1.e+36f ;
		FPSN_WJ:missing_value = 1.e+36f ;
	float FPSN_WP(time, lndgrid) ;
		FPSN_WP:long_name = "Product-limited photosynthesis" ;
		FPSN_WP:units = "umol/m2s" ;
		FPSN_WP:cell_methods = "time: mean" ;
		FPSN_WP:_FillValue = 1.e+36f ;
		FPSN_WP:missing_value = 1.e+36f ;
	float FROOTC(time, lndgrid) ;
		FROOTC:long_name = "fine root C" ;
		FROOTC:units = "gC/m^2" ;
		FROOTC:cell_methods = "time: mean" ;
		FROOTC:_FillValue = 1.e+36f ;
		FROOTC:missing_value = 1.e+36f ;
	float FROOTC_ALLOC(time, lndgrid) ;
		FROOTC_ALLOC:long_name = "fine root C allocation" ;
		FROOTC_ALLOC:units = "gC/m^2/s" ;
		FROOTC_ALLOC:cell_methods = "time: mean" ;
		FROOTC_ALLOC:_FillValue = 1.e+36f ;
		FROOTC_ALLOC:missing_value = 1.e+36f ;
	float FROOTC_LOSS(time, lndgrid) ;
		FROOTC_LOSS:long_name = "fine root C loss" ;
		FROOTC_LOSS:units = "gC/m^2/s" ;
		FROOTC_LOSS:cell_methods = "time: mean" ;
		FROOTC_LOSS:_FillValue = 1.e+36f ;
		FROOTC_LOSS:missing_value = 1.e+36f ;
	float FROOTN(time, lndgrid) ;
		FROOTN:long_name = "fine root N" ;
		FROOTN:units = "gN/m^2" ;
		FROOTN:cell_methods = "time: mean" ;
		FROOTN:_FillValue = 1.e+36f ;
		FROOTN:missing_value = 1.e+36f ;
	float FROST_TABLE(time, lndgrid) ;
		FROST_TABLE:long_name = "frost table depth (vegetated landunits only)" ;
		FROST_TABLE:units = "m" ;
		FROST_TABLE:cell_methods = "time: mean" ;
		FROST_TABLE:_FillValue = 1.e+36f ;
		FROST_TABLE:missing_value = 1.e+36f ;
	float FSA(time, lndgrid) ;
		FSA:long_name = "absorbed solar radiation" ;
		FSA:units = "W/m^2" ;
		FSA:cell_methods = "time: mean" ;
		FSA:_FillValue = 1.e+36f ;
		FSA:missing_value = 1.e+36f ;
	float FSAT(time, lndgrid) ;
		FSAT:long_name = "fractional area with water table at surface" ;
		FSAT:units = "unitless" ;
		FSAT:cell_methods = "time: mean" ;
		FSAT:_FillValue = 1.e+36f ;
		FSAT:missing_value = 1.e+36f ;
	float FSA_R(time, lndgrid) ;
		FSA_R:long_name = "Rural absorbed solar radiation" ;
		FSA_R:units = "W/m^2" ;
		FSA_R:cell_methods = "time: mean" ;
		FSA_R:_FillValue = 1.e+36f ;
		FSA_R:missing_value = 1.e+36f ;
	float FSA_U(time, lndgrid) ;
		FSA_U:long_name = "Urban absorbed solar radiation" ;
		FSA_U:units = "W/m^2" ;
		FSA_U:cell_methods = "time: mean" ;
		FSA_U:_FillValue = 1.e+36f ;
		FSA_U:missing_value = 1.e+36f ;
	float FSDS(time, lndgrid) ;
		FSDS:long_name = "atmospheric incident solar radiation" ;
		FSDS:units = "W/m^2" ;
		FSDS:cell_methods = "time: mean" ;
		FSDS:_FillValue = 1.e+36f ;
		FSDS:missing_value = 1.e+36f ;
	float FSDSND(time, lndgrid) ;
		FSDSND:long_name = "direct nir incident solar radiation" ;
		FSDSND:units = "W/m^2" ;
		FSDSND:cell_methods = "time: mean" ;
		FSDSND:_FillValue = 1.e+36f ;
		FSDSND:missing_value = 1.e+36f ;
	float FSDSNDLN(time, lndgrid) ;
		FSDSNDLN:long_name = "direct nir incident solar radiation at local noon" ;
		FSDSNDLN:units = "W/m^2" ;
		FSDSNDLN:cell_methods = "time: mean" ;
		FSDSNDLN:_FillValue = 1.e+36f ;
		FSDSNDLN:missing_value = 1.e+36f ;
	float FSDSNI(time, lndgrid) ;
		FSDSNI:long_name = "diffuse nir incident solar radiation" ;
		FSDSNI:units = "W/m^2" ;
		FSDSNI:cell_methods = "time: mean" ;
		FSDSNI:_FillValue = 1.e+36f ;
		FSDSNI:missing_value = 1.e+36f ;
	float FSDSVD(time, lndgrid) ;
		FSDSVD:long_name = "direct vis incident solar radiation" ;
		FSDSVD:units = "W/m^2" ;
		FSDSVD:cell_methods = "time: mean" ;
		FSDSVD:_FillValue = 1.e+36f ;
		FSDSVD:missing_value = 1.e+36f ;
	float FSDSVDLN(time, lndgrid) ;
		FSDSVDLN:long_name = "direct vis incident solar radiation at local noon" ;
		FSDSVDLN:units = "W/m^2" ;
		FSDSVDLN:cell_methods = "time: mean" ;
		FSDSVDLN:_FillValue = 1.e+36f ;
		FSDSVDLN:missing_value = 1.e+36f ;
	float FSDSVI(time, lndgrid) ;
		FSDSVI:long_name = "diffuse vis incident solar radiation" ;
		FSDSVI:units = "W/m^2" ;
		FSDSVI:cell_methods = "time: mean" ;
		FSDSVI:_FillValue = 1.e+36f ;
		FSDSVI:missing_value = 1.e+36f ;
	float FSDSVILN(time, lndgrid) ;
		FSDSVILN:long_name = "diffuse vis incident solar radiation at local noon" ;
		FSDSVILN:units = "W/m^2" ;
		FSDSVILN:cell_methods = "time: mean" ;
		FSDSVILN:_FillValue = 1.e+36f ;
		FSDSVILN:missing_value = 1.e+36f ;
	float FSH(time, lndgrid) ;
		FSH:long_name = "sensible heat" ;
		FSH:units = "W/m^2" ;
		FSH:cell_methods = "time: mean" ;
		FSH:_FillValue = 1.e+36f ;
		FSH:missing_value = 1.e+36f ;
	float FSH_G(time, lndgrid) ;
		FSH_G:long_name = "sensible heat from ground" ;
		FSH_G:units = "W/m^2" ;
		FSH_G:cell_methods = "time: mean" ;
		FSH_G:_FillValue = 1.e+36f ;
		FSH_G:missing_value = 1.e+36f ;
	float FSH_NODYNLNDUSE(time, lndgrid) ;
		FSH_NODYNLNDUSE:long_name = "sensible heat not including correction for land use change" ;
		FSH_NODYNLNDUSE:units = "W/m^2" ;
		FSH_NODYNLNDUSE:cell_methods = "time: mean" ;
		FSH_NODYNLNDUSE:_FillValue = 1.e+36f ;
		FSH_NODYNLNDUSE:missing_value = 1.e+36f ;
	float FSH_R(time, lndgrid) ;
		FSH_R:long_name = "Rural sensible heat" ;
		FSH_R:units = "W/m^2" ;
		FSH_R:cell_methods = "time: mean" ;
		FSH_R:_FillValue = 1.e+36f ;
		FSH_R:missing_value = 1.e+36f ;
	float FSH_U(time, lndgrid) ;
		FSH_U:long_name = "Urban sensible heat" ;
		FSH_U:units = "W/m^2" ;
		FSH_U:cell_methods = "time: mean" ;
		FSH_U:_FillValue = 1.e+36f ;
		FSH_U:missing_value = 1.e+36f ;
	float FSH_V(time, lndgrid) ;
		FSH_V:long_name = "sensible heat from veg" ;
		FSH_V:units = "W/m^2" ;
		FSH_V:cell_methods = "time: mean" ;
		FSH_V:_FillValue = 1.e+36f ;
		FSH_V:missing_value = 1.e+36f ;
	float FSM(time, lndgrid) ;
		FSM:long_name = "snow melt heat flux" ;
		FSM:units = "W/m^2" ;
		FSM:cell_methods = "time: mean" ;
		FSM:_FillValue = 1.e+36f ;
		FSM:missing_value = 1.e+36f ;
	float FSM_R(time, lndgrid) ;
		FSM_R:long_name = "Rural snow melt heat flux" ;
		FSM_R:units = "W/m^2" ;
		FSM_R:cell_methods = "time: mean" ;
		FSM_R:_FillValue = 1.e+36f ;
		FSM_R:missing_value = 1.e+36f ;
	float FSM_U(time, lndgrid) ;
		FSM_U:long_name = "Urban snow melt heat flux" ;
		FSM_U:units = "W/m^2" ;
		FSM_U:cell_methods = "time: mean" ;
		FSM_U:_FillValue = 1.e+36f ;
		FSM_U:missing_value = 1.e+36f ;
	float FSNO(time, lndgrid) ;
		FSNO:long_name = "fraction of ground covered by snow" ;
		FSNO:units = "unitless" ;
		FSNO:cell_methods = "time: mean" ;
		FSNO:_FillValue = 1.e+36f ;
		FSNO:missing_value = 1.e+36f ;
	float FSNO_EFF(time, lndgrid) ;
		FSNO_EFF:long_name = "effective fraction of ground covered by snow" ;
		FSNO_EFF:units = "unitless" ;
		FSNO_EFF:cell_methods = "time: mean" ;
		FSNO_EFF:_FillValue = 1.e+36f ;
		FSNO_EFF:missing_value = 1.e+36f ;
	float FSR(time, lndgrid) ;
		FSR:long_name = "reflected solar radiation" ;
		FSR:units = "W/m^2" ;
		FSR:cell_methods = "time: mean" ;
		FSR:_FillValue = 1.e+36f ;
		FSR:missing_value = 1.e+36f ;
	float FSRND(time, lndgrid) ;
		FSRND:long_name = "direct nir reflected solar radiation" ;
		FSRND:units = "W/m^2" ;
		FSRND:cell_methods = "time: mean" ;
		FSRND:_FillValue = 1.e+36f ;
		FSRND:missing_value = 1.e+36f ;
	float FSRNDLN(time, lndgrid) ;
		FSRNDLN:long_name = "direct nir reflected solar radiation at local noon" ;
		FSRNDLN:units = "W/m^2" ;
		FSRNDLN:cell_methods = "time: mean" ;
		FSRNDLN:_FillValue = 1.e+36f ;
		FSRNDLN:missing_value = 1.e+36f ;
	float FSRNI(time, lndgrid) ;
		FSRNI:long_name = "diffuse nir reflected solar radiation" ;
		FSRNI:units = "W/m^2" ;
		FSRNI:cell_methods = "time: mean" ;
		FSRNI:_FillValue = 1.e+36f ;
		FSRNI:missing_value = 1.e+36f ;
	float FSRVD(time, lndgrid) ;
		FSRVD:long_name = "direct vis reflected solar radiation" ;
		FSRVD:units = "W/m^2" ;
		FSRVD:cell_methods = "time: mean" ;
		FSRVD:_FillValue = 1.e+36f ;
		FSRVD:missing_value = 1.e+36f ;
	float FSRVDLN(time, lndgrid) ;
		FSRVDLN:long_name = "direct vis reflected solar radiation at local noon" ;
		FSRVDLN:units = "W/m^2" ;
		FSRVDLN:cell_methods = "time: mean" ;
		FSRVDLN:_FillValue = 1.e+36f ;
		FSRVDLN:missing_value = 1.e+36f ;
	float FSRVI(time, lndgrid) ;
		FSRVI:long_name = "diffuse vis reflected solar radiation" ;
		FSRVI:units = "W/m^2" ;
		FSRVI:cell_methods = "time: mean" ;
		FSRVI:_FillValue = 1.e+36f ;
		FSRVI:missing_value = 1.e+36f ;
	float FUELC(time, lndgrid) ;
		FUELC:long_name = "fuel load" ;
		FUELC:units = "gC/m^2" ;
		FUELC:cell_methods = "time: mean" ;
		FUELC:_FillValue = 1.e+36f ;
		FUELC:missing_value = 1.e+36f ;
	float F_DENIT(time, lndgrid) ;
		F_DENIT:long_name = "denitrification flux" ;
		F_DENIT:units = "gN/m^2/s" ;
		F_DENIT:cell_methods = "time: mean" ;
		F_DENIT:_FillValue = 1.e+36f ;
		F_DENIT:missing_value = 1.e+36f ;
	float F_DENIT_vr(time, levdcmp, lndgrid) ;
		F_DENIT_vr:long_name = "denitrification flux" ;
		F_DENIT_vr:units = "gN/m^3/s" ;
		F_DENIT_vr:cell_methods = "time: mean" ;
		F_DENIT_vr:_FillValue = 1.e+36f ;
		F_DENIT_vr:missing_value = 1.e+36f ;
	float F_N2O_DENIT(time, lndgrid) ;
		F_N2O_DENIT:long_name = "denitrification N2O flux" ;
		F_N2O_DENIT:units = "gN/m^2/s" ;
		F_N2O_DENIT:cell_methods = "time: mean" ;
		F_N2O_DENIT:_FillValue = 1.e+36f ;
		F_N2O_DENIT:missing_value = 1.e+36f ;
	float F_N2O_NIT(time, lndgrid) ;
		F_N2O_NIT:long_name = "nitrification N2O flux" ;
		F_N2O_NIT:units = "gN/m^2/s" ;
		F_N2O_NIT:cell_methods = "time: mean" ;
		F_N2O_NIT:_FillValue = 1.e+36f ;
		F_N2O_NIT:missing_value = 1.e+36f ;
	float F_NIT(time, lndgrid) ;
		F_NIT:long_name = "nitrification flux" ;
		F_NIT:units = "gN/m^2/s" ;
		F_NIT:cell_methods = "time: mean" ;
		F_NIT:_FillValue = 1.e+36f ;
		F_NIT:missing_value = 1.e+36f ;
	float F_NIT_vr(time, levdcmp, lndgrid) ;
		F_NIT_vr:long_name = "nitrification flux" ;
		F_NIT_vr:units = "gN/m^3/s" ;
		F_NIT_vr:cell_methods = "time: mean" ;
		F_NIT_vr:_FillValue = 1.e+36f ;
		F_NIT_vr:missing_value = 1.e+36f ;
	float GC_HEAT1(time, lndgrid) ;
		GC_HEAT1:long_name = "initial gridcell total heat content" ;
		GC_HEAT1:units = "J/m^2" ;
		GC_HEAT1:cell_methods = "time: mean" ;
		GC_HEAT1:_FillValue = 1.e+36f ;
		GC_HEAT1:missing_value = 1.e+36f ;
	float GC_ICE1(time, lndgrid) ;
		GC_ICE1:long_name = "initial gridcell total ice content" ;
		GC_ICE1:units = "mm" ;
		GC_ICE1:cell_methods = "time: mean" ;
		GC_ICE1:_FillValue = 1.e+36f ;
		GC_ICE1:missing_value = 1.e+36f ;
	float GC_LIQ1(time, lndgrid) ;
		GC_LIQ1:long_name = "initial gridcell total liq content" ;
		GC_LIQ1:units = "mm" ;
		GC_LIQ1:cell_methods = "time: mean" ;
		GC_LIQ1:_FillValue = 1.e+36f ;
		GC_LIQ1:missing_value = 1.e+36f ;
	float GPP(time, lndgrid) ;
		GPP:long_name = "gross primary production" ;
		GPP:units = "gC/m^2/s" ;
		GPP:cell_methods = "time: mean" ;
		GPP:_FillValue = 1.e+36f ;
		GPP:missing_value = 1.e+36f ;
	float GR(time, lndgrid) ;
		GR:long_name = "total growth respiration" ;
		GR:units = "gC/m^2/s" ;
		GR:cell_methods = "time: mean" ;
		GR:_FillValue = 1.e+36f ;
		GR:missing_value = 1.e+36f ;
	float GROSS_NMIN(time, lndgrid) ;
		GROSS_NMIN:long_name = "gross rate of N mineralization" ;
		GROSS_NMIN:units = "gN/m^2/s" ;
		GROSS_NMIN:cell_methods = "time: mean" ;
		GROSS_NMIN:_FillValue = 1.e+36f ;
		GROSS_NMIN:missing_value = 1.e+36f ;
	float H2OCAN(time, lndgrid) ;
		H2OCAN:long_name = "intercepted water" ;
		H2OCAN:units = "mm" ;
		H2OCAN:cell_methods = "time: mean" ;
		H2OCAN:_FillValue = 1.e+36f ;
		H2OCAN:missing_value = 1.e+36f ;
	float H2OSFC(time, lndgrid) ;
		H2OSFC:long_name = "surface water depth" ;
		H2OSFC:units = "mm" ;
		H2OSFC:cell_methods = "time: mean" ;
		H2OSFC:_FillValue = 1.e+36f ;
		H2OSFC:missing_value = 1.e+36f ;
	float H2OSNO(time, lndgrid) ;
		H2OSNO:long_name = "snow depth (liquid water)" ;
		H2OSNO:units = "mm" ;
		H2OSNO:cell_methods = "time: mean" ;
		H2OSNO:_FillValue = 1.e+36f ;
		H2OSNO:missing_value = 1.e+36f ;
	float H2OSNO_TOP(time, lndgrid) ;
		H2OSNO_TOP:long_name = "mass of snow in top snow layer" ;
		H2OSNO_TOP:units = "kg/m2" ;
		H2OSNO_TOP:cell_methods = "time: mean" ;
		H2OSNO_TOP:_FillValue = 1.e+36f ;
		H2OSNO_TOP:missing_value = 1.e+36f ;
	float H2OSOI(time, levgrnd, lndgrid) ;
		H2OSOI:long_name = "volumetric soil water (vegetated landunits only)" ;
		H2OSOI:units = "mm3/mm3" ;
		H2OSOI:cell_methods = "time: mean" ;
		H2OSOI:_FillValue = 1.e+36f ;
		H2OSOI:missing_value = 1.e+36f ;
	float HC(time, lndgrid) ;
		HC:long_name = "heat content of soil/snow/lake" ;
		HC:units = "MJ/m2" ;
		HC:cell_methods = "time: mean" ;
		HC:_FillValue = 1.e+36f ;
		HC:missing_value = 1.e+36f ;
	float HCSOI(time, lndgrid) ;
		HCSOI:long_name = "soil heat content" ;
		HCSOI:units = "MJ/m2" ;
		HCSOI:cell_methods = "time: mean" ;
		HCSOI:_FillValue = 1.e+36f ;
		HCSOI:missing_value = 1.e+36f ;
	float HEAT_FROM_AC(time, lndgrid) ;
		HEAT_FROM_AC:long_name = "sensible heat flux put into canyon due to heat removed from air conditioning" ;
		HEAT_FROM_AC:units = "W/m^2" ;
		HEAT_FROM_AC:cell_methods = "time: mean" ;
		HEAT_FROM_AC:_FillValue = 1.e+36f ;
		HEAT_FROM_AC:missing_value = 1.e+36f ;
	float HR(time, lndgrid) ;
		HR:long_name = "total heterotrophic respiration" ;
		HR:units = "gC/m^2/s" ;
		HR:cell_methods = "time: mean" ;
		HR:_FillValue = 1.e+36f ;
		HR:missing_value = 1.e+36f ;
	float HR_vr(time, levdcmp, lndgrid) ;
		HR_vr:long_name = "total vertically resolved heterotrophic respiration" ;
		HR_vr:units = "gC/m^3/s" ;
		HR_vr:cell_methods = "time: mean" ;
		HR_vr:_FillValue = 1.e+36f ;
		HR_vr:missing_value = 1.e+36f ;
	float HTOP(time, lndgrid) ;
		HTOP:long_name = "canopy top" ;
		HTOP:units = "m" ;
		HTOP:cell_methods = "time: mean" ;
		HTOP:_FillValue = 1.e+36f ;
		HTOP:missing_value = 1.e+36f ;
	float INT_SNOW(time, lndgrid) ;
		INT_SNOW:long_name = "accumulated swe (vegetated landunits only)" ;
		INT_SNOW:units = "mm" ;
		INT_SNOW:cell_methods = "time: mean" ;
		INT_SNOW:_FillValue = 1.e+36f ;
		INT_SNOW:missing_value = 1.e+36f ;
	float LAISHA(time, lndgrid) ;
		LAISHA:long_name = "shaded projected leaf area index" ;
		LAISHA:units = "none" ;
		LAISHA:cell_methods = "time: mean" ;
		LAISHA:_FillValue = 1.e+36f ;
		LAISHA:missing_value = 1.e+36f ;
	float LAISUN(time, lndgrid) ;
		LAISUN:long_name = "sunlit projected leaf area index" ;
		LAISUN:units = "none" ;
		LAISUN:cell_methods = "time: mean" ;
		LAISUN:_FillValue = 1.e+36f ;
		LAISUN:missing_value = 1.e+36f ;
	float LAKEICEFRAC(time, levlak, lndgrid) ;
		LAKEICEFRAC:long_name = "lake layer ice mass fraction" ;
		LAKEICEFRAC:units = "unitless" ;
		LAKEICEFRAC:cell_methods = "time: mean" ;
		LAKEICEFRAC:_FillValue = 1.e+36f ;
		LAKEICEFRAC:missing_value = 1.e+36f ;
	float LAKEICETHICK(time, lndgrid) ;
		LAKEICETHICK:long_name = "thickness of lake ice (including physical expansion on freezing)" ;
		LAKEICETHICK:units = "m" ;
		LAKEICETHICK:cell_methods = "time: mean" ;
		LAKEICETHICK:_FillValue = 1.e+36f ;
		LAKEICETHICK:missing_value = 1.e+36f ;
	float LAND_UPTAKE(time, lndgrid) ;
		LAND_UPTAKE:long_name = "NEE minus LAND_USE_FLUX, negative for update" ;
		LAND_UPTAKE:units = "gC/m^2/s" ;
		LAND_UPTAKE:cell_methods = "time: mean" ;
		LAND_UPTAKE:_FillValue = 1.e+36f ;
		LAND_UPTAKE:missing_value = 1.e+36f ;
	float LAND_USE_FLUX(time, lndgrid) ;
		LAND_USE_FLUX:long_name = "total C emitted from land cover conversion and wood product pools" ;
		LAND_USE_FLUX:units = "gC/m^2/s" ;
		LAND_USE_FLUX:cell_methods = "time: mean" ;
		LAND_USE_FLUX:_FillValue = 1.e+36f ;
		LAND_USE_FLUX:missing_value = 1.e+36f ;
	float LEAFC(time, lndgrid) ;
		LEAFC:long_name = "leaf C" ;
		LEAFC:units = "gC/m^2" ;
		LEAFC:cell_methods = "time: mean" ;
		LEAFC:_FillValue = 1.e+36f ;
		LEAFC:missing_value = 1.e+36f ;
	float LEAFC_ALLOC(time, lndgrid) ;
		LEAFC_ALLOC:long_name = "leaf C allocation" ;
		LEAFC_ALLOC:units = "gC/m^2/s" ;
		LEAFC_ALLOC:cell_methods = "time: mean" ;
		LEAFC_ALLOC:_FillValue = 1.e+36f ;
		LEAFC_ALLOC:missing_value = 1.e+36f ;
	float LEAFC_LOSS(time, lndgrid) ;
		LEAFC_LOSS:long_name = "leaf C loss" ;
		LEAFC_LOSS:units = "gC/m^2/s" ;
		LEAFC_LOSS:cell_methods = "time: mean" ;
		LEAFC_LOSS:_FillValue = 1.e+36f ;
		LEAFC_LOSS:missing_value = 1.e+36f ;
	float LEAFN(time, lndgrid) ;
		LEAFN:long_name = "leaf N" ;
		LEAFN:units = "gN/m^2" ;
		LEAFN:cell_methods = "time: mean" ;
		LEAFN:_FillValue = 1.e+36f ;
		LEAFN:missing_value = 1.e+36f ;
	float LEAF_MR(time, lndgrid) ;
		LEAF_MR:long_name = "leaf maintenance respiration" ;
		LEAF_MR:units = "gC/m^2/s" ;
		LEAF_MR:cell_methods = "time: mean" ;
		LEAF_MR:_FillValue = 1.e+36f ;
		LEAF_MR:missing_value = 1.e+36f ;
	float LFC2(time, lndgrid) ;
		LFC2:long_name = "conversion area fraction of BET and BDT that burned in this timestep" ;
		LFC2:units = "per timestep" ;
		LFC2:cell_methods = "time: mean" ;
		LFC2:_FillValue = 1.e+36f ;
		LFC2:missing_value = 1.e+36f ;
	float LF_CONV_CFLUX(time, lndgrid) ;
		LF_CONV_CFLUX:long_name = "conversion carbon due to BET and BDT area decreasing" ;
		LF_CONV_CFLUX:units = "gC/m^2/s" ;
		LF_CONV_CFLUX:cell_methods = "time: mean" ;
		LF_CONV_CFLUX:_FillValue = 1.e+36f ;
		LF_CONV_CFLUX:missing_value = 1.e+36f ;
	float LITFALL(time, lndgrid) ;
		LITFALL:long_name = "litterfall (leaves and fine roots)" ;
		LITFALL:units = "gC/m^2/s" ;
		LITFALL:cell_methods = "time: mean" ;
		LITFALL:_FillValue = 1.e+36f ;
		LITFALL:missing_value = 1.e+36f ;
	float LITHR(time, lndgrid) ;
		LITHR:long_name = "litter heterotrophic respiration" ;
		LITHR:units = "gC/m^2/s" ;
		LITHR:cell_methods = "time: mean" ;
		LITHR:_FillValue = 1.e+36f ;
		LITHR:missing_value = 1.e+36f ;
	float LITR1C(time, lndgrid) ;
		LITR1C:long_name = "LITR1 C" ;
		LITR1C:units = "gC/m^2" ;
		LITR1C:cell_methods = "time: mean" ;
		LITR1C:_FillValue = 1.e+36f ;
		LITR1C:missing_value = 1.e+36f ;
	float LITR1C_TO_SOIL1C(time, lndgrid) ;
		LITR1C_TO_SOIL1C:long_name = "decomp. of litter 1 C to soil 1 C" ;
		LITR1C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR1C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR1C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR1C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR1C_vr(time, levdcmp, lndgrid) ;
		LITR1C_vr:long_name = "LITR1 C (vertically resolved)" ;
		LITR1C_vr:units = "gC/m^3" ;
		LITR1C_vr:cell_methods = "time: mean" ;
		LITR1C_vr:_FillValue = 1.e+36f ;
		LITR1C_vr:missing_value = 1.e+36f ;
	float LITR1N(time, lndgrid) ;
		LITR1N:long_name = "LITR1 N" ;
		LITR1N:units = "gN/m^2" ;
		LITR1N:cell_methods = "time: mean" ;
		LITR1N:_FillValue = 1.e+36f ;
		LITR1N:missing_value = 1.e+36f ;
	float LITR1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR1N_TNDNCY_VERT_TRANS:long_name = "litter 1 N tendency due to vertical transport" ;
		LITR1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR1N_TO_SOIL1N(time, lndgrid) ;
		LITR1N_TO_SOIL1N:long_name = "decomp. of litter 1 N to soil 1 N" ;
		LITR1N_TO_SOIL1N:units = "gN/m^2" ;
		LITR1N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR1N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR1N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR1N_vr(time, levdcmp, lndgrid) ;
		LITR1N_vr:long_name = "LITR1 N (vertically resolved)" ;
		LITR1N_vr:units = "gN/m^3" ;
		LITR1N_vr:cell_methods = "time: mean" ;
		LITR1N_vr:_FillValue = 1.e+36f ;
		LITR1N_vr:missing_value = 1.e+36f ;
	float LITR1_HR(time, lndgrid) ;
		LITR1_HR:long_name = "Het. Resp. from litter 1" ;
		LITR1_HR:units = "gC/m^2/s" ;
		LITR1_HR:cell_methods = "time: mean" ;
		LITR1_HR:_FillValue = 1.e+36f ;
		LITR1_HR:missing_value = 1.e+36f ;
	float LITR2C(time, lndgrid) ;
		LITR2C:long_name = "LITR2 C" ;
		LITR2C:units = "gC/m^2" ;
		LITR2C:cell_methods = "time: mean" ;
		LITR2C:_FillValue = 1.e+36f ;
		LITR2C:missing_value = 1.e+36f ;
	float LITR2C_TO_SOIL1C(time, lndgrid) ;
		LITR2C_TO_SOIL1C:long_name = "decomp. of litter 2 C to soil 1 C" ;
		LITR2C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR2C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR2C_vr(time, levdcmp, lndgrid) ;
		LITR2C_vr:long_name = "LITR2 C (vertically resolved)" ;
		LITR2C_vr:units = "gC/m^3" ;
		LITR2C_vr:cell_methods = "time: mean" ;
		LITR2C_vr:_FillValue = 1.e+36f ;
		LITR2C_vr:missing_value = 1.e+36f ;
	float LITR2N(time, lndgrid) ;
		LITR2N:long_name = "LITR2 N" ;
		LITR2N:units = "gN/m^2" ;
		LITR2N:cell_methods = "time: mean" ;
		LITR2N:_FillValue = 1.e+36f ;
		LITR2N:missing_value = 1.e+36f ;
	float LITR2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR2N_TNDNCY_VERT_TRANS:long_name = "litter 2 N tendency due to vertical transport" ;
		LITR2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR2N_TO_SOIL1N(time, lndgrid) ;
		LITR2N_TO_SOIL1N:long_name = "decomp. of litter 2 N to soil 1 N" ;
		LITR2N_TO_SOIL1N:units = "gN/m^2" ;
		LITR2N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR2N_vr(time, levdcmp, lndgrid) ;
		LITR2N_vr:long_name = "LITR2 N (vertically resolved)" ;
		LITR2N_vr:units = "gN/m^3" ;
		LITR2N_vr:cell_methods = "time: mean" ;
		LITR2N_vr:_FillValue = 1.e+36f ;
		LITR2N_vr:missing_value = 1.e+36f ;
	float LITR2_HR(time, lndgrid) ;
		LITR2_HR:long_name = "Het. Resp. from litter 2" ;
		LITR2_HR:units = "gC/m^2/s" ;
		LITR2_HR:cell_methods = "time: mean" ;
		LITR2_HR:_FillValue = 1.e+36f ;
		LITR2_HR:missing_value = 1.e+36f ;
	float LITR3C(time, lndgrid) ;
		LITR3C:long_name = "LITR3 C" ;
		LITR3C:units = "gC/m^2" ;
		LITR3C:cell_methods = "time: mean" ;
		LITR3C:_FillValue = 1.e+36f ;
		LITR3C:missing_value = 1.e+36f ;
	float LITR3C_TO_SOIL2C(time, lndgrid) ;
		LITR3C_TO_SOIL2C:long_name = "decomp. of litter 3 C to soil 2 C" ;
		LITR3C_TO_SOIL2C:units = "gC/m^2/s" ;
		LITR3C_TO_SOIL2C:cell_methods = "time: mean" ;
		LITR3C_TO_SOIL2C:_FillValue = 1.e+36f ;
		LITR3C_TO_SOIL2C:missing_value = 1.e+36f ;
	float LITR3C_vr(time, levdcmp, lndgrid) ;
		LITR3C_vr:long_name = "LITR3 C (vertically resolved)" ;
		LITR3C_vr:units = "gC/m^3" ;
		LITR3C_vr:cell_methods = "time: mean" ;
		LITR3C_vr:_FillValue = 1.e+36f ;
		LITR3C_vr:missing_value = 1.e+36f ;
	float LITR3N(time, lndgrid) ;
		LITR3N:long_name = "LITR3 N" ;
		LITR3N:units = "gN/m^2" ;
		LITR3N:cell_methods = "time: mean" ;
		LITR3N:_FillValue = 1.e+36f ;
		LITR3N:missing_value = 1.e+36f ;
	float LITR3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR3N_TNDNCY_VERT_TRANS:long_name = "litter 3 N tendency due to vertical transport" ;
		LITR3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR3N_TO_SOIL2N(time, lndgrid) ;
		LITR3N_TO_SOIL2N:long_name = "decomp. of litter 3 N to soil 2 N" ;
		LITR3N_TO_SOIL2N:units = "gN/m^2" ;
		LITR3N_TO_SOIL2N:cell_methods = "time: mean" ;
		LITR3N_TO_SOIL2N:_FillValue = 1.e+36f ;
		LITR3N_TO_SOIL2N:missing_value = 1.e+36f ;
	float LITR3N_vr(time, levdcmp, lndgrid) ;
		LITR3N_vr:long_name = "LITR3 N (vertically resolved)" ;
		LITR3N_vr:units = "gN/m^3" ;
		LITR3N_vr:cell_methods = "time: mean" ;
		LITR3N_vr:_FillValue = 1.e+36f ;
		LITR3N_vr:missing_value = 1.e+36f ;
	float LITR3_HR(time, lndgrid) ;
		LITR3_HR:long_name = "Het. Resp. from litter 3" ;
		LITR3_HR:units = "gC/m^2/s" ;
		LITR3_HR:cell_methods = "time: mean" ;
		LITR3_HR:_FillValue = 1.e+36f ;
		LITR3_HR:missing_value = 1.e+36f ;
	float LITTERC(time, lndgrid) ;
		LITTERC:long_name = "litter C" ;
		LITTERC:units = "gC/m^2" ;
		LITTERC:cell_methods = "time: mean" ;
		LITTERC:_FillValue = 1.e+36f ;
		LITTERC:missing_value = 1.e+36f ;
	float LITTERC_HR(time, lndgrid) ;
		LITTERC_HR:long_name = "litter C heterotrophic respiration" ;
		LITTERC_HR:units = "gC/m^2/s" ;
		LITTERC_HR:cell_methods = "time: mean" ;
		LITTERC_HR:_FillValue = 1.e+36f ;
		LITTERC_HR:missing_value = 1.e+36f ;
	float LITTERC_LOSS(time, lndgrid) ;
		LITTERC_LOSS:long_name = "litter C loss" ;
		LITTERC_LOSS:units = "gC/m^2/s" ;
		LITTERC_LOSS:cell_methods = "time: mean" ;
		LITTERC_LOSS:_FillValue = 1.e+36f ;
		LITTERC_LOSS:missing_value = 1.e+36f ;
	float LIVECROOTC(time, lndgrid) ;
		LIVECROOTC:long_name = "live coarse root C" ;
		LIVECROOTC:units = "gC/m^2" ;
		LIVECROOTC:cell_methods = "time: mean" ;
		LIVECROOTC:_FillValue = 1.e+36f ;
		LIVECROOTC:missing_value = 1.e+36f ;
	float LIVECROOTN(time, lndgrid) ;
		LIVECROOTN:long_name = "live coarse root N" ;
		LIVECROOTN:units = "gN/m^2" ;
		LIVECROOTN:cell_methods = "time: mean" ;
		LIVECROOTN:_FillValue = 1.e+36f ;
		LIVECROOTN:missing_value = 1.e+36f ;
	float LIVESTEMC(time, lndgrid) ;
		LIVESTEMC:long_name = "live stem C" ;
		LIVESTEMC:units = "gC/m^2" ;
		LIVESTEMC:cell_methods = "time: mean" ;
		LIVESTEMC:_FillValue = 1.e+36f ;
		LIVESTEMC:missing_value = 1.e+36f ;
	float LIVESTEMN(time, lndgrid) ;
		LIVESTEMN:long_name = "live stem N" ;
		LIVESTEMN:units = "gN/m^2" ;
		LIVESTEMN:cell_methods = "time: mean" ;
		LIVESTEMN:_FillValue = 1.e+36f ;
		LIVESTEMN:missing_value = 1.e+36f ;
	float MEG_acetaldehyde(time, lndgrid) ;
		MEG_acetaldehyde:long_name = "MEGAN flux" ;
		MEG_acetaldehyde:units = "kg/m2/sec" ;
		MEG_acetaldehyde:cell_methods = "time: mean" ;
		MEG_acetaldehyde:_FillValue = 1.e+36f ;
		MEG_acetaldehyde:missing_value = 1.e+36f ;
	float MEG_acetic_acid(time, lndgrid) ;
		MEG_acetic_acid:long_name = "MEGAN flux" ;
		MEG_acetic_acid:units = "kg/m2/sec" ;
		MEG_acetic_acid:cell_methods = "time: mean" ;
		MEG_acetic_acid:_FillValue = 1.e+36f ;
		MEG_acetic_acid:missing_value = 1.e+36f ;
	float MEG_acetone(time, lndgrid) ;
		MEG_acetone:long_name = "MEGAN flux" ;
		MEG_acetone:units = "kg/m2/sec" ;
		MEG_acetone:cell_methods = "time: mean" ;
		MEG_acetone:_FillValue = 1.e+36f ;
		MEG_acetone:missing_value = 1.e+36f ;
	float MEG_carene_3(time, lndgrid) ;
		MEG_carene_3:long_name = "MEGAN flux" ;
		MEG_carene_3:units = "kg/m2/sec" ;
		MEG_carene_3:cell_methods = "time: mean" ;
		MEG_carene_3:_FillValue = 1.e+36f ;
		MEG_carene_3:missing_value = 1.e+36f ;
	float MEG_ethanol(time, lndgrid) ;
		MEG_ethanol:long_name = "MEGAN flux" ;
		MEG_ethanol:units = "kg/m2/sec" ;
		MEG_ethanol:cell_methods = "time: mean" ;
		MEG_ethanol:_FillValue = 1.e+36f ;
		MEG_ethanol:missing_value = 1.e+36f ;
	float MEG_formaldehyde(time, lndgrid) ;
		MEG_formaldehyde:long_name = "MEGAN flux" ;
		MEG_formaldehyde:units = "kg/m2/sec" ;
		MEG_formaldehyde:cell_methods = "time: mean" ;
		MEG_formaldehyde:_FillValue = 1.e+36f ;
		MEG_formaldehyde:missing_value = 1.e+36f ;
	float MEG_isoprene(time, lndgrid) ;
		MEG_isoprene:long_name = "MEGAN flux" ;
		MEG_isoprene:units = "kg/m2/sec" ;
		MEG_isoprene:cell_methods = "time: mean" ;
		MEG_isoprene:_FillValue = 1.e+36f ;
		MEG_isoprene:missing_value = 1.e+36f ;
	float MEG_methanol(time, lndgrid) ;
		MEG_methanol:long_name = "MEGAN flux" ;
		MEG_methanol:units = "kg/m2/sec" ;
		MEG_methanol:cell_methods = "time: mean" ;
		MEG_methanol:_FillValue = 1.e+36f ;
		MEG_methanol:missing_value = 1.e+36f ;
	float MEG_pinene_a(time, lndgrid) ;
		MEG_pinene_a:long_name = "MEGAN flux" ;
		MEG_pinene_a:units = "kg/m2/sec" ;
		MEG_pinene_a:cell_methods = "time: mean" ;
		MEG_pinene_a:_FillValue = 1.e+36f ;
		MEG_pinene_a:missing_value = 1.e+36f ;
	float MEG_thujene_a(time, lndgrid) ;
		MEG_thujene_a:long_name = "MEGAN flux" ;
		MEG_thujene_a:units = "kg/m2/sec" ;
		MEG_thujene_a:cell_methods = "time: mean" ;
		MEG_thujene_a:_FillValue = 1.e+36f ;
		MEG_thujene_a:missing_value = 1.e+36f ;
	float MR(time, lndgrid) ;
		MR:long_name = "maintenance respiration" ;
		MR:units = "gC/m^2/s" ;
		MR:cell_methods = "time: mean" ;
		MR:_FillValue = 1.e+36f ;
		MR:missing_value = 1.e+36f ;
	float M_LITR1C_TO_LEACHING(time, lndgrid) ;
		M_LITR1C_TO_LEACHING:long_name = "litter 1 C leaching loss" ;
		M_LITR1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR2C_TO_LEACHING(time, lndgrid) ;
		M_LITR2C_TO_LEACHING:long_name = "litter 2 C leaching loss" ;
		M_LITR2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR3C_TO_LEACHING(time, lndgrid) ;
		M_LITR3C_TO_LEACHING:long_name = "litter 3 C leaching loss" ;
		M_LITR3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR3C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL1C_TO_LEACHING(time, lndgrid) ;
		M_SOIL1C_TO_LEACHING:long_name = "soil 1 C leaching loss" ;
		M_SOIL1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL2C_TO_LEACHING(time, lndgrid) ;
		M_SOIL2C_TO_LEACHING:long_name = "soil 2 C leaching loss" ;
		M_SOIL2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL3C_TO_LEACHING(time, lndgrid) ;
		M_SOIL3C_TO_LEACHING:long_name = "soil 3 C leaching loss" ;
		M_SOIL3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL3C_TO_LEACHING:missing_value = 1.e+36f ;
	float NBP(time, lndgrid) ;
		NBP:long_name = "net biome production, includes fire, landuse, and harvest flux, positive for sink" ;
		NBP:units = "gC/m^2/s" ;
		NBP:cell_methods = "time: mean" ;
		NBP:_FillValue = 1.e+36f ;
		NBP:missing_value = 1.e+36f ;
	float NDEPLOY(time, lndgrid) ;
		NDEPLOY:long_name = "total N deployed in new growth" ;
		NDEPLOY:units = "gN/m^2/s" ;
		NDEPLOY:cell_methods = "time: mean" ;
		NDEPLOY:_FillValue = 1.e+36f ;
		NDEPLOY:missing_value = 1.e+36f ;
	float NDEP_TO_SMINN(time, lndgrid) ;
		NDEP_TO_SMINN:long_name = "atmospheric N deposition to soil mineral N" ;
		NDEP_TO_SMINN:units = "gN/m^2/s" ;
		NDEP_TO_SMINN:cell_methods = "time: mean" ;
		NDEP_TO_SMINN:_FillValue = 1.e+36f ;
		NDEP_TO_SMINN:missing_value = 1.e+36f ;
	float NEE(time, lndgrid) ;
		NEE:long_name = "net ecosystem exchange of carbon, includes fire, landuse, harvest, and hrv_xsmrpool flux, positive for source" ;
		NEE:units = "gC/m^2/s" ;
		NEE:cell_methods = "time: mean" ;
		NEE:_FillValue = 1.e+36f ;
		NEE:missing_value = 1.e+36f ;
	float NEM(time, lndgrid) ;
		NEM:long_name = "Gridcell net adjustment to NEE passed to atm. for methane production" ;
		NEM:units = "gC/m2/s" ;
		NEM:cell_methods = "time: mean" ;
		NEM:_FillValue = 1.e+36f ;
		NEM:missing_value = 1.e+36f ;
	float NEP(time, lndgrid) ;
		NEP:long_name = "net ecosystem production, excludes fire, landuse, and harvest flux, positive for sink" ;
		NEP:units = "gC/m^2/s" ;
		NEP:cell_methods = "time: mean" ;
		NEP:_FillValue = 1.e+36f ;
		NEP:missing_value = 1.e+36f ;
	float NET_NMIN(time, lndgrid) ;
		NET_NMIN:long_name = "net rate of N mineralization" ;
		NET_NMIN:units = "gN/m^2/s" ;
		NET_NMIN:cell_methods = "time: mean" ;
		NET_NMIN:_FillValue = 1.e+36f ;
		NET_NMIN:missing_value = 1.e+36f ;
	float NFIRE(time, lndgrid) ;
		NFIRE:long_name = "timestep fire counts valid only in Reg.C" ;
		NFIRE:units = "counts/km2/timestep" ;
		NFIRE:cell_methods = "time: mean" ;
		NFIRE:_FillValue = 1.e+36f ;
		NFIRE:missing_value = 1.e+36f ;
	float NFIX_TO_SMINN(time, lndgrid) ;
		NFIX_TO_SMINN:long_name = "symbiotic/asymbiotic N fixation to soil mineral N" ;
		NFIX_TO_SMINN:units = "gN/m^2/s" ;
		NFIX_TO_SMINN:cell_methods = "time: mean" ;
		NFIX_TO_SMINN:_FillValue = 1.e+36f ;
		NFIX_TO_SMINN:missing_value = 1.e+36f ;
	float NPP(time, lndgrid) ;
		NPP:long_name = "net primary production" ;
		NPP:units = "gC/m^2/s" ;
		NPP:cell_methods = "time: mean" ;
		NPP:_FillValue = 1.e+36f ;
		NPP:missing_value = 1.e+36f ;
	float OCDEP(time, lndgrid) ;
		OCDEP:long_name = "total OC deposition (dry+wet) from atmosphere" ;
		OCDEP:units = "kg/m^2/s" ;
		OCDEP:cell_methods = "time: mean" ;
		OCDEP:_FillValue = 1.e+36f ;
		OCDEP:missing_value = 1.e+36f ;
	float O_SCALAR(time, levdcmp, lndgrid) ;
		O_SCALAR:long_name = "fraction by which decomposition is reduced due to anoxia" ;
		O_SCALAR:units = "unitless" ;
		O_SCALAR:cell_methods = "time: mean" ;
		O_SCALAR:_FillValue = 1.e+36f ;
		O_SCALAR:missing_value = 1.e+36f ;
	float PARVEGLN(time, lndgrid) ;
		PARVEGLN:long_name = "absorbed par by vegetation at local noon" ;
		PARVEGLN:units = "W/m^2" ;
		PARVEGLN:cell_methods = "time: mean" ;
		PARVEGLN:_FillValue = 1.e+36f ;
		PARVEGLN:missing_value = 1.e+36f ;
	float PBOT(time, lndgrid) ;
		PBOT:long_name = "atmospheric pressure" ;
		PBOT:units = "Pa" ;
		PBOT:cell_methods = "time: mean" ;
		PBOT:_FillValue = 1.e+36f ;
		PBOT:missing_value = 1.e+36f ;
	float PCH4(time, lndgrid) ;
		PCH4:long_name = "atmospheric partial pressure of CH4" ;
		PCH4:units = "Pa" ;
		PCH4:cell_methods = "time: mean" ;
		PCH4:_FillValue = 1.e+36f ;
		PCH4:missing_value = 1.e+36f ;
	float PCO2(time, lndgrid) ;
		PCO2:long_name = "atmospheric partial pressure of CO2" ;
		PCO2:units = "Pa" ;
		PCO2:cell_methods = "time: mean" ;
		PCO2:_FillValue = 1.e+36f ;
		PCO2:missing_value = 1.e+36f ;
	float PFT_CTRUNC(time, lndgrid) ;
		PFT_CTRUNC:long_name = "pft-level sink for C truncation" ;
		PFT_CTRUNC:units = "gC/m^2" ;
		PFT_CTRUNC:cell_methods = "time: mean" ;
		PFT_CTRUNC:_FillValue = 1.e+36f ;
		PFT_CTRUNC:missing_value = 1.e+36f ;
	float PFT_FIRE_CLOSS(time, lndgrid) ;
		PFT_FIRE_CLOSS:long_name = "total pft-level fire C loss for non-peat fires outside land-type converted region" ;
		PFT_FIRE_CLOSS:units = "gC/m^2/s" ;
		PFT_FIRE_CLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_CLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_CLOSS:missing_value = 1.e+36f ;
	float PFT_FIRE_NLOSS(time, lndgrid) ;
		PFT_FIRE_NLOSS:long_name = "total pft-level fire N loss" ;
		PFT_FIRE_NLOSS:units = "gN/m^2/s" ;
		PFT_FIRE_NLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_NLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_NLOSS:missing_value = 1.e+36f ;
	float PFT_NTRUNC(time, lndgrid) ;
		PFT_NTRUNC:long_name = "pft-level sink for N truncation" ;
		PFT_NTRUNC:units = "gN/m^2" ;
		PFT_NTRUNC:cell_methods = "time: mean" ;
		PFT_NTRUNC:_FillValue = 1.e+36f ;
		PFT_NTRUNC:missing_value = 1.e+36f ;
	float PLANT_NDEMAND(time, lndgrid) ;
		PLANT_NDEMAND:long_name = "N flux required to support initial GPP" ;
		PLANT_NDEMAND:units = "gN/m^2/s" ;
		PLANT_NDEMAND:cell_methods = "time: mean" ;
		PLANT_NDEMAND:_FillValue = 1.e+36f ;
		PLANT_NDEMAND:missing_value = 1.e+36f ;
	float POTENTIAL_IMMOB(time, lndgrid) ;
		POTENTIAL_IMMOB:long_name = "potential N immobilization" ;
		POTENTIAL_IMMOB:units = "gN/m^2/s" ;
		POTENTIAL_IMMOB:cell_methods = "time: mean" ;
		POTENTIAL_IMMOB:_FillValue = 1.e+36f ;
		POTENTIAL_IMMOB:missing_value = 1.e+36f ;
	float POT_F_DENIT(time, lndgrid) ;
		POT_F_DENIT:long_name = "potential denitrification flux" ;
		POT_F_DENIT:units = "gN/m^2/s" ;
		POT_F_DENIT:cell_methods = "time: mean" ;
		POT_F_DENIT:_FillValue = 1.e+36f ;
		POT_F_DENIT:missing_value = 1.e+36f ;
	float POT_F_NIT(time, lndgrid) ;
		POT_F_NIT:long_name = "potential nitrification flux" ;
		POT_F_NIT:units = "gN/m^2/s" ;
		POT_F_NIT:cell_methods = "time: mean" ;
		POT_F_NIT:_FillValue = 1.e+36f ;
		POT_F_NIT:missing_value = 1.e+36f ;
	float PROD100C(time, lndgrid) ;
		PROD100C:long_name = "100-yr wood product C" ;
		PROD100C:units = "gC/m^2" ;
		PROD100C:cell_methods = "time: mean" ;
		PROD100C:_FillValue = 1.e+36f ;
		PROD100C:missing_value = 1.e+36f ;
	float PROD100C_LOSS(time, lndgrid) ;
		PROD100C_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100C_LOSS:units = "gC/m^2/s" ;
		PROD100C_LOSS:cell_methods = "time: mean" ;
		PROD100C_LOSS:_FillValue = 1.e+36f ;
		PROD100C_LOSS:missing_value = 1.e+36f ;
	float PROD100N(time, lndgrid) ;
		PROD100N:long_name = "100-yr wood product N" ;
		PROD100N:units = "gN/m^2" ;
		PROD100N:cell_methods = "time: mean" ;
		PROD100N:_FillValue = 1.e+36f ;
		PROD100N:missing_value = 1.e+36f ;
	float PROD100N_LOSS(time, lndgrid) ;
		PROD100N_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100N_LOSS:units = "gN/m^2/s" ;
		PROD100N_LOSS:cell_methods = "time: mean" ;
		PROD100N_LOSS:_FillValue = 1.e+36f ;
		PROD100N_LOSS:missing_value = 1.e+36f ;
	float PROD10C(time, lndgrid) ;
		PROD10C:long_name = "10-yr wood product C" ;
		PROD10C:units = "gC/m^2" ;
		PROD10C:cell_methods = "time: mean" ;
		PROD10C:_FillValue = 1.e+36f ;
		PROD10C:missing_value = 1.e+36f ;
	float PROD10C_LOSS(time, lndgrid) ;
		PROD10C_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10C_LOSS:units = "gC/m^2/s" ;
		PROD10C_LOSS:cell_methods = "time: mean" ;
		PROD10C_LOSS:_FillValue = 1.e+36f ;
		PROD10C_LOSS:missing_value = 1.e+36f ;
	float PROD10N(time, lndgrid) ;
		PROD10N:long_name = "10-yr wood product N" ;
		PROD10N:units = "gN/m^2" ;
		PROD10N:cell_methods = "time: mean" ;
		PROD10N:_FillValue = 1.e+36f ;
		PROD10N:missing_value = 1.e+36f ;
	float PROD10N_LOSS(time, lndgrid) ;
		PROD10N_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10N_LOSS:units = "gN/m^2/s" ;
		PROD10N_LOSS:cell_methods = "time: mean" ;
		PROD10N_LOSS:_FillValue = 1.e+36f ;
		PROD10N_LOSS:missing_value = 1.e+36f ;
	float PRODUCT_CLOSS(time, lndgrid) ;
		PRODUCT_CLOSS:long_name = "total carbon loss from wood product pools" ;
		PRODUCT_CLOSS:units = "gC/m^2/s" ;
		PRODUCT_CLOSS:cell_methods = "time: mean" ;
		PRODUCT_CLOSS:_FillValue = 1.e+36f ;
		PRODUCT_CLOSS:missing_value = 1.e+36f ;
	float PRODUCT_NLOSS(time, lndgrid) ;
		PRODUCT_NLOSS:long_name = "total N loss from wood product pools" ;
		PRODUCT_NLOSS:units = "gN/m^2/s" ;
		PRODUCT_NLOSS:cell_methods = "time: mean" ;
		PRODUCT_NLOSS:_FillValue = 1.e+36f ;
		PRODUCT_NLOSS:missing_value = 1.e+36f ;
	float PSNSHA(time, lndgrid) ;
		PSNSHA:long_name = "shaded leaf photosynthesis" ;
		PSNSHA:units = "umolCO2/m^2/s" ;
		PSNSHA:cell_methods = "time: mean" ;
		PSNSHA:_FillValue = 1.e+36f ;
		PSNSHA:missing_value = 1.e+36f ;
	float PSNSHADE_TO_CPOOL(time, lndgrid) ;
		PSNSHADE_TO_CPOOL:long_name = "C fixation from shaded canopy" ;
		PSNSHADE_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSHADE_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSHADE_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSHADE_TO_CPOOL:missing_value = 1.e+36f ;
	float PSNSUN(time, lndgrid) ;
		PSNSUN:long_name = "sunlit leaf photosynthesis" ;
		PSNSUN:units = "umolCO2/m^2/s" ;
		PSNSUN:cell_methods = "time: mean" ;
		PSNSUN:_FillValue = 1.e+36f ;
		PSNSUN:missing_value = 1.e+36f ;
	float PSNSUN_TO_CPOOL(time, lndgrid) ;
		PSNSUN_TO_CPOOL:long_name = "C fixation from sunlit canopy" ;
		PSNSUN_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSUN_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSUN_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSUN_TO_CPOOL:missing_value = 1.e+36f ;
	float Q2M(time, lndgrid) ;
		Q2M:long_name = "2m specific humidity" ;
		Q2M:units = "kg/kg" ;
		Q2M:cell_methods = "time: mean" ;
		Q2M:_FillValue = 1.e+36f ;
		Q2M:missing_value = 1.e+36f ;
	float QBOT(time, lndgrid) ;
		QBOT:long_name = "atmospheric specific humidity" ;
		QBOT:units = "kg/kg" ;
		QBOT:cell_methods = "time: mean" ;
		QBOT:_FillValue = 1.e+36f ;
		QBOT:missing_value = 1.e+36f ;
	float QCHARGE(time, lndgrid) ;
		QCHARGE:long_name = "aquifer recharge rate (vegetated landunits only)" ;
		QCHARGE:units = "mm/s" ;
		QCHARGE:cell_methods = "time: mean" ;
		QCHARGE:_FillValue = 1.e+36f ;
		QCHARGE:missing_value = 1.e+36f ;
	float QDRAI(time, lndgrid) ;
		QDRAI:long_name = "sub-surface drainage" ;
		QDRAI:units = "mm/s" ;
		QDRAI:cell_methods = "time: mean" ;
		QDRAI:_FillValue = 1.e+36f ;
		QDRAI:missing_value = 1.e+36f ;
	float QDRAI_PERCH(time, lndgrid) ;
		QDRAI_PERCH:long_name = "perched wt drainage" ;
		QDRAI_PERCH:units = "mm/s" ;
		QDRAI_PERCH:cell_methods = "time: mean" ;
		QDRAI_PERCH:_FillValue = 1.e+36f ;
		QDRAI_PERCH:missing_value = 1.e+36f ;
	float QDRAI_XS(time, lndgrid) ;
		QDRAI_XS:long_name = "saturation excess drainage" ;
		QDRAI_XS:units = "mm/s" ;
		QDRAI_XS:cell_methods = "time: mean" ;
		QDRAI_XS:_FillValue = 1.e+36f ;
		QDRAI_XS:missing_value = 1.e+36f ;
	float QDRIP(time, lndgrid) ;
		QDRIP:long_name = "throughfall" ;
		QDRIP:units = "mm/s" ;
		QDRIP:cell_methods = "time: mean" ;
		QDRIP:_FillValue = 1.e+36f ;
		QDRIP:missing_value = 1.e+36f ;
	float QFLOOD(time, lndgrid) ;
		QFLOOD:long_name = "runoff from river flooding" ;
		QFLOOD:units = "mm/s" ;
		QFLOOD:cell_methods = "time: mean" ;
		QFLOOD:_FillValue = 1.e+36f ;
		QFLOOD:missing_value = 1.e+36f ;
	float QFLX_ICE_DYNBAL(time, lndgrid) ;
		QFLX_ICE_DYNBAL:long_name = "ice dynamic land cover change conversion runoff flux" ;
		QFLX_ICE_DYNBAL:units = "mm/s" ;
		QFLX_ICE_DYNBAL:cell_methods = "time: mean" ;
		QFLX_ICE_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_ICE_DYNBAL:missing_value = 1.e+36f ;
	float QFLX_LIQ_DYNBAL(time, lndgrid) ;
		QFLX_LIQ_DYNBAL:long_name = "liq dynamic land cover change conversion runoff flux" ;
		QFLX_LIQ_DYNBAL:units = "mm/s" ;
		QFLX_LIQ_DYNBAL:cell_methods = "time: mean" ;
		QFLX_LIQ_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_LIQ_DYNBAL:missing_value = 1.e+36f ;
	float QH2OSFC(time, lndgrid) ;
		QH2OSFC:long_name = "surface water runoff" ;
		QH2OSFC:units = "mm/s" ;
		QH2OSFC:cell_methods = "time: mean" ;
		QH2OSFC:_FillValue = 1.e+36f ;
		QH2OSFC:missing_value = 1.e+36f ;
	float QINFL(time, lndgrid) ;
		QINFL:long_name = "infiltration" ;
		QINFL:units = "mm/s" ;
		QINFL:cell_methods = "time: mean" ;
		QINFL:_FillValue = 1.e+36f ;
		QINFL:missing_value = 1.e+36f ;
	float QINTR(time, lndgrid) ;
		QINTR:long_name = "interception" ;
		QINTR:units = "mm/s" ;
		QINTR:cell_methods = "time: mean" ;
		QINTR:_FillValue = 1.e+36f ;
		QINTR:missing_value = 1.e+36f ;
	float QIRRIG(time, lndgrid) ;
		QIRRIG:long_name = "water added through irrigation" ;
		QIRRIG:units = "mm/s" ;
		QIRRIG:cell_methods = "time: mean" ;
		QIRRIG:_FillValue = 1.e+36f ;
		QIRRIG:missing_value = 1.e+36f ;
	float QOVER(time, lndgrid) ;
		QOVER:long_name = "surface runoff" ;
		QOVER:units = "mm/s" ;
		QOVER:cell_methods = "time: mean" ;
		QOVER:_FillValue = 1.e+36f ;
		QOVER:missing_value = 1.e+36f ;
	float QOVER_LAG(time, lndgrid) ;
		QOVER_LAG:long_name = "time-lagged surface runoff for soil columns" ;
		QOVER_LAG:units = "mm/s" ;
		QOVER_LAG:cell_methods = "time: mean" ;
		QOVER_LAG:_FillValue = 1.e+36f ;
		QOVER_LAG:missing_value = 1.e+36f ;
	float QRGWL(time, lndgrid) ;
		QRGWL:long_name = "surface runoff at glaciers (liquid only), wetlands, lakes" ;
		QRGWL:units = "mm/s" ;
		QRGWL:cell_methods = "time: mean" ;
		QRGWL:_FillValue = 1.e+36f ;
		QRGWL:missing_value = 1.e+36f ;
	float QRUNOFF(time, lndgrid) ;
		QRUNOFF:long_name = "total liquid runoff (does not include QSNWCPICE)" ;
		QRUNOFF:units = "mm/s" ;
		QRUNOFF:cell_methods = "time: mean" ;
		QRUNOFF:_FillValue = 1.e+36f ;
		QRUNOFF:missing_value = 1.e+36f ;
	float QRUNOFF_NODYNLNDUSE(time, lndgrid) ;
		QRUNOFF_NODYNLNDUSE:long_name = "total liquid runoff (does not include QSNWCPICE) not including correction for land use change" ;
		QRUNOFF_NODYNLNDUSE:units = "mm/s" ;
		QRUNOFF_NODYNLNDUSE:cell_methods = "time: mean" ;
		QRUNOFF_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QRUNOFF_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QRUNOFF_R(time, lndgrid) ;
		QRUNOFF_R:long_name = "Rural total runoff" ;
		QRUNOFF_R:units = "mm/s" ;
		QRUNOFF_R:cell_methods = "time: mean" ;
		QRUNOFF_R:_FillValue = 1.e+36f ;
		QRUNOFF_R:missing_value = 1.e+36f ;
	float QRUNOFF_U(time, lndgrid) ;
		QRUNOFF_U:long_name = "Urban total runoff" ;
		QRUNOFF_U:units = "mm/s" ;
		QRUNOFF_U:cell_methods = "time: mean" ;
		QRUNOFF_U:_FillValue = 1.e+36f ;
		QRUNOFF_U:missing_value = 1.e+36f ;
	float QSNOMELT(time, lndgrid) ;
		QSNOMELT:long_name = "snow melt" ;
		QSNOMELT:units = "mm/s" ;
		QSNOMELT:cell_methods = "time: mean" ;
		QSNOMELT:_FillValue = 1.e+36f ;
		QSNOMELT:missing_value = 1.e+36f ;
	float QSNWCPICE(time, lndgrid) ;
		QSNWCPICE:long_name = "excess snowfall due to snow capping" ;
		QSNWCPICE:units = "mm/s" ;
		QSNWCPICE:cell_methods = "time: mean" ;
		QSNWCPICE:_FillValue = 1.e+36f ;
		QSNWCPICE:missing_value = 1.e+36f ;
	float QSNWCPICE_NODYNLNDUSE(time, lndgrid) ;
		QSNWCPICE_NODYNLNDUSE:long_name = "excess snowfall due to snow capping not including correction for land use change" ;
		QSNWCPICE_NODYNLNDUSE:units = "mm H2O/s" ;
		QSNWCPICE_NODYNLNDUSE:cell_methods = "time: mean" ;
		QSNWCPICE_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QSNWCPICE_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QSOIL(time, lndgrid) ;
		QSOIL:long_name = "Ground evaporation (soil/snow evaporation + soil/snow sublimation - dew)" ;
		QSOIL:units = "mm/s" ;
		QSOIL:cell_methods = "time: mean" ;
		QSOIL:_FillValue = 1.e+36f ;
		QSOIL:missing_value = 1.e+36f ;
	float QVEGE(time, lndgrid) ;
		QVEGE:long_name = "canopy evaporation" ;
		QVEGE:units = "mm/s" ;
		QVEGE:cell_methods = "time: mean" ;
		QVEGE:_FillValue = 1.e+36f ;
		QVEGE:missing_value = 1.e+36f ;
	float QVEGT(time, lndgrid) ;
		QVEGT:long_name = "canopy transpiration" ;
		QVEGT:units = "mm/s" ;
		QVEGT:cell_methods = "time: mean" ;
		QVEGT:_FillValue = 1.e+36f ;
		QVEGT:missing_value = 1.e+36f ;
	float RAIN(time, lndgrid) ;
		RAIN:long_name = "atmospheric rain" ;
		RAIN:units = "mm/s" ;
		RAIN:cell_methods = "time: mean" ;
		RAIN:_FillValue = 1.e+36f ;
		RAIN:missing_value = 1.e+36f ;
	float RETRANSN(time, lndgrid) ;
		RETRANSN:long_name = "plant pool of retranslocated N" ;
		RETRANSN:units = "gN/m^2" ;
		RETRANSN:cell_methods = "time: mean" ;
		RETRANSN:_FillValue = 1.e+36f ;
		RETRANSN:missing_value = 1.e+36f ;
	float RETRANSN_TO_NPOOL(time, lndgrid) ;
		RETRANSN_TO_NPOOL:long_name = "deployment of retranslocated N" ;
		RETRANSN_TO_NPOOL:units = "gN/m^2/s" ;
		RETRANSN_TO_NPOOL:cell_methods = "time: mean" ;
		RETRANSN_TO_NPOOL:_FillValue = 1.e+36f ;
		RETRANSN_TO_NPOOL:missing_value = 1.e+36f ;
	float RH2M(time, lndgrid) ;
		RH2M:long_name = "2m relative humidity" ;
		RH2M:units = "%" ;
		RH2M:cell_methods = "time: mean" ;
		RH2M:_FillValue = 1.e+36f ;
		RH2M:missing_value = 1.e+36f ;
	float RH2M_R(time, lndgrid) ;
		RH2M_R:long_name = "Rural 2m specific humidity" ;
		RH2M_R:units = "%" ;
		RH2M_R:cell_methods = "time: mean" ;
		RH2M_R:_FillValue = 1.e+36f ;
		RH2M_R:missing_value = 1.e+36f ;
	float RH2M_U(time, lndgrid) ;
		RH2M_U:long_name = "Urban 2m relative humidity" ;
		RH2M_U:units = "%" ;
		RH2M_U:cell_methods = "time: mean" ;
		RH2M_U:_FillValue = 1.e+36f ;
		RH2M_U:missing_value = 1.e+36f ;
	float RR(time, lndgrid) ;
		RR:long_name = "root respiration (fine root MR + total root GR)" ;
		RR:units = "gC/m^2/s" ;
		RR:cell_methods = "time: mean" ;
		RR:_FillValue = 1.e+36f ;
		RR:missing_value = 1.e+36f ;
	float SABG(time, lndgrid) ;
		SABG:long_name = "solar rad absorbed by ground" ;
		SABG:units = "W/m^2" ;
		SABG:cell_methods = "time: mean" ;
		SABG:_FillValue = 1.e+36f ;
		SABG:missing_value = 1.e+36f ;
	float SABG_PEN(time, lndgrid) ;
		SABG_PEN:long_name = "Rural solar rad penetrating top soil or snow layer" ;
		SABG_PEN:units = "watt/m^2" ;
		SABG_PEN:cell_methods = "time: mean" ;
		SABG_PEN:_FillValue = 1.e+36f ;
		SABG_PEN:missing_value = 1.e+36f ;
	float SABV(time, lndgrid) ;
		SABV:long_name = "solar rad absorbed by veg" ;
		SABV:units = "W/m^2" ;
		SABV:cell_methods = "time: mean" ;
		SABV:_FillValue = 1.e+36f ;
		SABV:missing_value = 1.e+36f ;
	float SEEDC(time, lndgrid) ;
		SEEDC:long_name = "pool for seeding new PFTs" ;
		SEEDC:units = "gC/m^2" ;
		SEEDC:cell_methods = "time: mean" ;
		SEEDC:_FillValue = 1.e+36f ;
		SEEDC:missing_value = 1.e+36f ;
	float SEEDN(time, lndgrid) ;
		SEEDN:long_name = "pool for seeding new PFTs" ;
		SEEDN:units = "gN/m^2" ;
		SEEDN:cell_methods = "time: mean" ;
		SEEDN:_FillValue = 1.e+36f ;
		SEEDN:missing_value = 1.e+36f ;
	float SMINN(time, lndgrid) ;
		SMINN:long_name = "soil mineral N" ;
		SMINN:units = "gN/m^2" ;
		SMINN:cell_methods = "time: mean" ;
		SMINN:_FillValue = 1.e+36f ;
		SMINN:missing_value = 1.e+36f ;
	float SMINN_TO_NPOOL(time, lndgrid) ;
		SMINN_TO_NPOOL:long_name = "deployment of soil mineral N uptake" ;
		SMINN_TO_NPOOL:units = "gN/m^2/s" ;
		SMINN_TO_NPOOL:cell_methods = "time: mean" ;
		SMINN_TO_NPOOL:_FillValue = 1.e+36f ;
		SMINN_TO_NPOOL:missing_value = 1.e+36f ;
	float SMINN_TO_PLANT(time, lndgrid) ;
		SMINN_TO_PLANT:long_name = "plant uptake of soil mineral N" ;
		SMINN_TO_PLANT:units = "gN/m^2/s" ;
		SMINN_TO_PLANT:cell_methods = "time: mean" ;
		SMINN_TO_PLANT:_FillValue = 1.e+36f ;
		SMINN_TO_PLANT:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L1(time, lndgrid) ;
		SMINN_TO_SOIL1N_L1:long_name = "mineral N flux for decomp. of LITR1to SOIL1" ;
		SMINN_TO_SOIL1N_L1:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L2(time, lndgrid) ;
		SMINN_TO_SOIL1N_L2:long_name = "mineral N flux for decomp. of LITR2to SOIL1" ;
		SMINN_TO_SOIL1N_L2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S2(time, lndgrid) ;
		SMINN_TO_SOIL1N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL1" ;
		SMINN_TO_SOIL1N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S3(time, lndgrid) ;
		SMINN_TO_SOIL1N_S3:long_name = "mineral N flux for decomp. of SOIL3to SOIL1" ;
		SMINN_TO_SOIL1N_S3:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_L3(time, lndgrid) ;
		SMINN_TO_SOIL2N_L3:long_name = "mineral N flux for decomp. of LITR3to SOIL2" ;
		SMINN_TO_SOIL2N_L3:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_L3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_L3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_L3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_S1(time, lndgrid) ;
		SMINN_TO_SOIL2N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL2" ;
		SMINN_TO_SOIL2N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S1(time, lndgrid) ;
		SMINN_TO_SOIL3N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL3" ;
		SMINN_TO_SOIL3N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S2(time, lndgrid) ;
		SMINN_TO_SOIL3N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL3" ;
		SMINN_TO_SOIL3N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S2:missing_value = 1.e+36f ;
	float SMIN_NH4(time, lndgrid) ;
		SMIN_NH4:long_name = "soil mineral NH4" ;
		SMIN_NH4:units = "gN/m^2" ;
		SMIN_NH4:cell_methods = "time: mean" ;
		SMIN_NH4:_FillValue = 1.e+36f ;
		SMIN_NH4:missing_value = 1.e+36f ;
	float SMIN_NH4_vr(time, levdcmp, lndgrid) ;
		SMIN_NH4_vr:long_name = "soil mineral NH4 (vert. res.)" ;
		SMIN_NH4_vr:units = "gN/m^3" ;
		SMIN_NH4_vr:cell_methods = "time: mean" ;
		SMIN_NH4_vr:_FillValue = 1.e+36f ;
		SMIN_NH4_vr:missing_value = 1.e+36f ;
	float SMIN_NO3(time, lndgrid) ;
		SMIN_NO3:long_name = "soil mineral NO3" ;
		SMIN_NO3:units = "gN/m^2" ;
		SMIN_NO3:cell_methods = "time: mean" ;
		SMIN_NO3:_FillValue = 1.e+36f ;
		SMIN_NO3:missing_value = 1.e+36f ;
	float SMIN_NO3_LEACHED(time, lndgrid) ;
		SMIN_NO3_LEACHED:long_name = "soil NO3 pool loss to leaching" ;
		SMIN_NO3_LEACHED:units = "gN/m^2/s" ;
		SMIN_NO3_LEACHED:cell_methods = "time: mean" ;
		SMIN_NO3_LEACHED:_FillValue = 1.e+36f ;
		SMIN_NO3_LEACHED:missing_value = 1.e+36f ;
	float SMIN_NO3_RUNOFF(time, lndgrid) ;
		SMIN_NO3_RUNOFF:long_name = "soil NO3 pool loss to runoff" ;
		SMIN_NO3_RUNOFF:units = "gN/m^2/s" ;
		SMIN_NO3_RUNOFF:cell_methods = "time: mean" ;
		SMIN_NO3_RUNOFF:_FillValue = 1.e+36f ;
		SMIN_NO3_RUNOFF:missing_value = 1.e+36f ;
	float SMIN_NO3_vr(time, levdcmp, lndgrid) ;
		SMIN_NO3_vr:long_name = "soil mineral NO3 (vert. res.)" ;
		SMIN_NO3_vr:units = "gN/m^3" ;
		SMIN_NO3_vr:cell_methods = "time: mean" ;
		SMIN_NO3_vr:_FillValue = 1.e+36f ;
		SMIN_NO3_vr:missing_value = 1.e+36f ;
	float SNOBCMCL(time, lndgrid) ;
		SNOBCMCL:long_name = "mass of BC in snow column" ;
		SNOBCMCL:units = "kg/m2" ;
		SNOBCMCL:cell_methods = "time: mean" ;
		SNOBCMCL:_FillValue = 1.e+36f ;
		SNOBCMCL:missing_value = 1.e+36f ;
	float SNOBCMSL(time, lndgrid) ;
		SNOBCMSL:long_name = "mass of BC in top snow layer" ;
		SNOBCMSL:units = "kg/m2" ;
		SNOBCMSL:cell_methods = "time: mean" ;
		SNOBCMSL:_FillValue = 1.e+36f ;
		SNOBCMSL:missing_value = 1.e+36f ;
	float SNODSTMCL(time, lndgrid) ;
		SNODSTMCL:long_name = "mass of dust in snow column" ;
		SNODSTMCL:units = "kg/m2" ;
		SNODSTMCL:cell_methods = "time: mean" ;
		SNODSTMCL:_FillValue = 1.e+36f ;
		SNODSTMCL:missing_value = 1.e+36f ;
	float SNODSTMSL(time, lndgrid) ;
		SNODSTMSL:long_name = "mass of dust in top snow layer" ;
		SNODSTMSL:units = "kg/m2" ;
		SNODSTMSL:cell_methods = "time: mean" ;
		SNODSTMSL:_FillValue = 1.e+36f ;
		SNODSTMSL:missing_value = 1.e+36f ;
	float SNOOCMCL(time, lndgrid) ;
		SNOOCMCL:long_name = "mass of OC in snow column" ;
		SNOOCMCL:units = "kg/m2" ;
		SNOOCMCL:cell_methods = "time: mean" ;
		SNOOCMCL:_FillValue = 1.e+36f ;
		SNOOCMCL:missing_value = 1.e+36f ;
	float SNOOCMSL(time, lndgrid) ;
		SNOOCMSL:long_name = "mass of OC in top snow layer" ;
		SNOOCMSL:units = "kg/m2" ;
		SNOOCMSL:cell_methods = "time: mean" ;
		SNOOCMSL:_FillValue = 1.e+36f ;
		SNOOCMSL:missing_value = 1.e+36f ;
	float SNOW(time, lndgrid) ;
		SNOW:long_name = "atmospheric snow" ;
		SNOW:units = "mm/s" ;
		SNOW:cell_methods = "time: mean" ;
		SNOW:_FillValue = 1.e+36f ;
		SNOW:missing_value = 1.e+36f ;
	float SNOWDP(time, lndgrid) ;
		SNOWDP:long_name = "gridcell mean snow height" ;
		SNOWDP:units = "m" ;
		SNOWDP:cell_methods = "time: mean" ;
		SNOWDP:_FillValue = 1.e+36f ;
		SNOWDP:missing_value = 1.e+36f ;
	float SNOWICE(time, lndgrid) ;
		SNOWICE:long_name = "snow ice" ;
		SNOWICE:units = "kg/m2" ;
		SNOWICE:cell_methods = "time: mean" ;
		SNOWICE:_FillValue = 1.e+36f ;
		SNOWICE:missing_value = 1.e+36f ;
	float SNOWLIQ(time, lndgrid) ;
		SNOWLIQ:long_name = "snow liquid water" ;
		SNOWLIQ:units = "kg/m2" ;
		SNOWLIQ:cell_methods = "time: mean" ;
		SNOWLIQ:_FillValue = 1.e+36f ;
		SNOWLIQ:missing_value = 1.e+36f ;
	float SNOW_DEPTH(time, lndgrid) ;
		SNOW_DEPTH:long_name = "snow height of snow covered area" ;
		SNOW_DEPTH:units = "m" ;
		SNOW_DEPTH:cell_methods = "time: mean" ;
		SNOW_DEPTH:_FillValue = 1.e+36f ;
		SNOW_DEPTH:missing_value = 1.e+36f ;
	float SNOW_SINKS(time, lndgrid) ;
		SNOW_SINKS:long_name = "snow sinks (liquid water)" ;
		SNOW_SINKS:units = "mm/s" ;
		SNOW_SINKS:cell_methods = "time: mean" ;
		SNOW_SINKS:_FillValue = 1.e+36f ;
		SNOW_SINKS:missing_value = 1.e+36f ;
	float SNOW_SOURCES(time, lndgrid) ;
		SNOW_SOURCES:long_name = "snow sources (liquid water)" ;
		SNOW_SOURCES:units = "mm/s" ;
		SNOW_SOURCES:cell_methods = "time: mean" ;
		SNOW_SOURCES:_FillValue = 1.e+36f ;
		SNOW_SOURCES:missing_value = 1.e+36f ;
	float SOIL1C(time, lndgrid) ;
		SOIL1C:long_name = "SOIL1 C" ;
		SOIL1C:units = "gC/m^2" ;
		SOIL1C:cell_methods = "time: mean" ;
		SOIL1C:_FillValue = 1.e+36f ;
		SOIL1C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL2C(time, lndgrid) ;
		SOIL1C_TO_SOIL2C:long_name = "decomp. of soil 1 C to soil 2 C" ;
		SOIL1C_TO_SOIL2C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL2C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL2C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL2C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL3C(time, lndgrid) ;
		SOIL1C_TO_SOIL3C:long_name = "decomp. of soil 1 C to soil 3 C" ;
		SOIL1C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL1C_vr(time, levdcmp, lndgrid) ;
		SOIL1C_vr:long_name = "SOIL1 C (vertically resolved)" ;
		SOIL1C_vr:units = "gC/m^3" ;
		SOIL1C_vr:cell_methods = "time: mean" ;
		SOIL1C_vr:_FillValue = 1.e+36f ;
		SOIL1C_vr:missing_value = 1.e+36f ;
	float SOIL1N(time, lndgrid) ;
		SOIL1N:long_name = "SOIL1 N" ;
		SOIL1N:units = "gN/m^2" ;
		SOIL1N:cell_methods = "time: mean" ;
		SOIL1N:_FillValue = 1.e+36f ;
		SOIL1N:missing_value = 1.e+36f ;
	float SOIL1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL1N_TNDNCY_VERT_TRANS:long_name = "soil 1 N tendency due to vertical transport" ;
		SOIL1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL2N(time, lndgrid) ;
		SOIL1N_TO_SOIL2N:long_name = "decomp. of soil 1 N to soil 2 N" ;
		SOIL1N_TO_SOIL2N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL2N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL2N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL2N:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL3N(time, lndgrid) ;
		SOIL1N_TO_SOIL3N:long_name = "decomp. of soil 1 N to soil 3 N" ;
		SOIL1N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL1N_vr(time, levdcmp, lndgrid) ;
		SOIL1N_vr:long_name = "SOIL1 N (vertically resolved)" ;
		SOIL1N_vr:units = "gN/m^3" ;
		SOIL1N_vr:cell_methods = "time: mean" ;
		SOIL1N_vr:_FillValue = 1.e+36f ;
		SOIL1N_vr:missing_value = 1.e+36f ;
	float SOIL1_HR_S2(time, lndgrid) ;
		SOIL1_HR_S2:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S2:units = "gC/m^2/s" ;
		SOIL1_HR_S2:cell_methods = "time: mean" ;
		SOIL1_HR_S2:_FillValue = 1.e+36f ;
		SOIL1_HR_S2:missing_value = 1.e+36f ;
	float SOIL1_HR_S3(time, lndgrid) ;
		SOIL1_HR_S3:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S3:units = "gC/m^2/s" ;
		SOIL1_HR_S3:cell_methods = "time: mean" ;
		SOIL1_HR_S3:_FillValue = 1.e+36f ;
		SOIL1_HR_S3:missing_value = 1.e+36f ;
	float SOIL2C(time, lndgrid) ;
		SOIL2C:long_name = "SOIL2 C" ;
		SOIL2C:units = "gC/m^2" ;
		SOIL2C:cell_methods = "time: mean" ;
		SOIL2C:_FillValue = 1.e+36f ;
		SOIL2C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL1C(time, lndgrid) ;
		SOIL2C_TO_SOIL1C:long_name = "decomp. of soil 2 C to soil 1 C" ;
		SOIL2C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL3C(time, lndgrid) ;
		SOIL2C_TO_SOIL3C:long_name = "decomp. of soil 2 C to soil 3 C" ;
		SOIL2C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL2C_vr(time, levdcmp, lndgrid) ;
		SOIL2C_vr:long_name = "SOIL2 C (vertically resolved)" ;
		SOIL2C_vr:units = "gC/m^3" ;
		SOIL2C_vr:cell_methods = "time: mean" ;
		SOIL2C_vr:_FillValue = 1.e+36f ;
		SOIL2C_vr:missing_value = 1.e+36f ;
	float SOIL2N(time, lndgrid) ;
		SOIL2N:long_name = "SOIL2 N" ;
		SOIL2N:units = "gN/m^2" ;
		SOIL2N:cell_methods = "time: mean" ;
		SOIL2N:_FillValue = 1.e+36f ;
		SOIL2N:missing_value = 1.e+36f ;
	float SOIL2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL2N_TNDNCY_VERT_TRANS:long_name = "soil 2 N tendency due to vertical transport" ;
		SOIL2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL1N(time, lndgrid) ;
		SOIL2N_TO_SOIL1N:long_name = "decomp. of soil 2 N to soil 1 N" ;
		SOIL2N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL3N(time, lndgrid) ;
		SOIL2N_TO_SOIL3N:long_name = "decomp. of soil 2 N to soil 3 N" ;
		SOIL2N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL2N_vr(time, levdcmp, lndgrid) ;
		SOIL2N_vr:long_name = "SOIL2 N (vertically resolved)" ;
		SOIL2N_vr:units = "gN/m^3" ;
		SOIL2N_vr:cell_methods = "time: mean" ;
		SOIL2N_vr:_FillValue = 1.e+36f ;
		SOIL2N_vr:missing_value = 1.e+36f ;
	float SOIL2_HR_S1(time, lndgrid) ;
		SOIL2_HR_S1:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S1:units = "gC/m^2/s" ;
		SOIL2_HR_S1:cell_methods = "time: mean" ;
		SOIL2_HR_S1:_FillValue = 1.e+36f ;
		SOIL2_HR_S1:missing_value = 1.e+36f ;
	float SOIL2_HR_S3(time, lndgrid) ;
		SOIL2_HR_S3:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S3:units = "gC/m^2/s" ;
		SOIL2_HR_S3:cell_methods = "time: mean" ;
		SOIL2_HR_S3:_FillValue = 1.e+36f ;
		SOIL2_HR_S3:missing_value = 1.e+36f ;
	float SOIL3C(time, lndgrid) ;
		SOIL3C:long_name = "SOIL3 C" ;
		SOIL3C:units = "gC/m^2" ;
		SOIL3C:cell_methods = "time: mean" ;
		SOIL3C:_FillValue = 1.e+36f ;
		SOIL3C:missing_value = 1.e+36f ;
	float SOIL3C_TO_SOIL1C(time, lndgrid) ;
		SOIL3C_TO_SOIL1C:long_name = "decomp. of soil 3 C to soil 1 C" ;
		SOIL3C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL3C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL3C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL3C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL3C_vr(time, levdcmp, lndgrid) ;
		SOIL3C_vr:long_name = "SOIL3 C (vertically resolved)" ;
		SOIL3C_vr:units = "gC/m^3" ;
		SOIL3C_vr:cell_methods = "time: mean" ;
		SOIL3C_vr:_FillValue = 1.e+36f ;
		SOIL3C_vr:missing_value = 1.e+36f ;
	float SOIL3N(time, lndgrid) ;
		SOIL3N:long_name = "SOIL3 N" ;
		SOIL3N:units = "gN/m^2" ;
		SOIL3N:cell_methods = "time: mean" ;
		SOIL3N:_FillValue = 1.e+36f ;
		SOIL3N:missing_value = 1.e+36f ;
	float SOIL3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL3N_TNDNCY_VERT_TRANS:long_name = "soil 3 N tendency due to vertical transport" ;
		SOIL3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL3N_TO_SOIL1N(time, lndgrid) ;
		SOIL3N_TO_SOIL1N:long_name = "decomp. of soil 3 N to soil 1 N" ;
		SOIL3N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL3N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL3N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL3N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL3N_vr(time, levdcmp, lndgrid) ;
		SOIL3N_vr:long_name = "SOIL3 N (vertically resolved)" ;
		SOIL3N_vr:units = "gN/m^3" ;
		SOIL3N_vr:cell_methods = "time: mean" ;
		SOIL3N_vr:_FillValue = 1.e+36f ;
		SOIL3N_vr:missing_value = 1.e+36f ;
	float SOIL3_HR(time, lndgrid) ;
		SOIL3_HR:long_name = "Het. Resp. from soil 3" ;
		SOIL3_HR:units = "gC/m^2/s" ;
		SOIL3_HR:cell_methods = "time: mean" ;
		SOIL3_HR:_FillValue = 1.e+36f ;
		SOIL3_HR:missing_value = 1.e+36f ;
	float SOILC(time, lndgrid) ;
		SOILC:long_name = "soil C" ;
		SOILC:units = "gC/m^2" ;
		SOILC:cell_methods = "time: mean" ;
		SOILC:_FillValue = 1.e+36f ;
		SOILC:missing_value = 1.e+36f ;
	float SOILC_HR(time, lndgrid) ;
		SOILC_HR:long_name = "soil C heterotrophic respiration" ;
		SOILC_HR:units = "gC/m^2/s" ;
		SOILC_HR:cell_methods = "time: mean" ;
		SOILC_HR:_FillValue = 1.e+36f ;
		SOILC_HR:missing_value = 1.e+36f ;
	float SOILC_LOSS(time, lndgrid) ;
		SOILC_LOSS:long_name = "soil C loss" ;
		SOILC_LOSS:units = "gC/m^2/s" ;
		SOILC_LOSS:cell_methods = "time: mean" ;
		SOILC_LOSS:_FillValue = 1.e+36f ;
		SOILC_LOSS:missing_value = 1.e+36f ;
	float SOILICE(time, levgrnd, lndgrid) ;
		SOILICE:long_name = "soil ice (vegetated landunits only)" ;
		SOILICE:units = "kg/m2" ;
		SOILICE:cell_methods = "time: mean" ;
		SOILICE:_FillValue = 1.e+36f ;
		SOILICE:missing_value = 1.e+36f ;
	float SOILLIQ(time, levgrnd, lndgrid) ;
		SOILLIQ:long_name = "soil liquid water (vegetated landunits only)" ;
		SOILLIQ:units = "kg/m2" ;
		SOILLIQ:cell_methods = "time: mean" ;
		SOILLIQ:_FillValue = 1.e+36f ;
		SOILLIQ:missing_value = 1.e+36f ;
	float SOILPSI(time, levgrnd, lndgrid) ;
		SOILPSI:long_name = "soil water potential in each soil layer" ;
		SOILPSI:units = "MPa" ;
		SOILPSI:cell_methods = "time: mean" ;
		SOILPSI:_FillValue = 1.e+36f ;
		SOILPSI:missing_value = 1.e+36f ;
	float SOILWATER_10CM(time, lndgrid) ;
		SOILWATER_10CM:long_name = "soil liquid water + ice in top 10cm of soil (veg landunits only)" ;
		SOILWATER_10CM:units = "kg/m2" ;
		SOILWATER_10CM:cell_methods = "time: mean" ;
		SOILWATER_10CM:_FillValue = 1.e+36f ;
		SOILWATER_10CM:missing_value = 1.e+36f ;
	float SOMC_FIRE(time, lndgrid) ;
		SOMC_FIRE:long_name = "C loss due to peat burning" ;
		SOMC_FIRE:units = "gC/m^2/s" ;
		SOMC_FIRE:cell_methods = "time: mean" ;
		SOMC_FIRE:_FillValue = 1.e+36f ;
		SOMC_FIRE:missing_value = 1.e+36f ;
	float SOMHR(time, lndgrid) ;
		SOMHR:long_name = "soil organic matter heterotrophic respiration" ;
		SOMHR:units = "gC/m^2/s" ;
		SOMHR:cell_methods = "time: mean" ;
		SOMHR:_FillValue = 1.e+36f ;
		SOMHR:missing_value = 1.e+36f ;
	float SOM_C_LEACHED(time, lndgrid) ;
		SOM_C_LEACHED:long_name = "total flux of C from SOM pools due to leaching" ;
		SOM_C_LEACHED:units = "gC/m^2/s" ;
		SOM_C_LEACHED:cell_methods = "time: mean" ;
		SOM_C_LEACHED:_FillValue = 1.e+36f ;
		SOM_C_LEACHED:missing_value = 1.e+36f ;
	float SR(time, lndgrid) ;
		SR:long_name = "total soil respiration (HR + root resp)" ;
		SR:units = "gC/m^2/s" ;
		SR:cell_methods = "time: mean" ;
		SR:_FillValue = 1.e+36f ;
		SR:missing_value = 1.e+36f ;
	float STORVEGC(time, lndgrid) ;
		STORVEGC:long_name = "stored vegetation carbon, excluding cpool" ;
		STORVEGC:units = "gC/m^2" ;
		STORVEGC:cell_methods = "time: mean" ;
		STORVEGC:_FillValue = 1.e+36f ;
		STORVEGC:missing_value = 1.e+36f ;
	float STORVEGN(time, lndgrid) ;
		STORVEGN:long_name = "stored vegetation nitrogen" ;
		STORVEGN:units = "gN/m^2" ;
		STORVEGN:cell_methods = "time: mean" ;
		STORVEGN:_FillValue = 1.e+36f ;
		STORVEGN:missing_value = 1.e+36f ;
	float SUPPLEMENT_TO_SMINN(time, lndgrid) ;
		SUPPLEMENT_TO_SMINN:long_name = "supplemental N supply" ;
		SUPPLEMENT_TO_SMINN:units = "gN/m^2/s" ;
		SUPPLEMENT_TO_SMINN:cell_methods = "time: mean" ;
		SUPPLEMENT_TO_SMINN:_FillValue = 1.e+36f ;
		SUPPLEMENT_TO_SMINN:missing_value = 1.e+36f ;
	float SoilAlpha(time, lndgrid) ;
		SoilAlpha:long_name = "factor limiting ground evap" ;
		SoilAlpha:units = "unitless" ;
		SoilAlpha:cell_methods = "time: mean" ;
		SoilAlpha:_FillValue = 1.e+36f ;
		SoilAlpha:missing_value = 1.e+36f ;
	float SoilAlpha_U(time, lndgrid) ;
		SoilAlpha_U:long_name = "urban factor limiting ground evap" ;
		SoilAlpha_U:units = "unitless" ;
		SoilAlpha_U:cell_methods = "time: mean" ;
		SoilAlpha_U:_FillValue = 1.e+36f ;
		SoilAlpha_U:missing_value = 1.e+36f ;
	float TAUX(time, lndgrid) ;
		TAUX:long_name = "zonal surface stress" ;
		TAUX:units = "kg/m/s^2" ;
		TAUX:cell_methods = "time: mean" ;
		TAUX:_FillValue = 1.e+36f ;
		TAUX:missing_value = 1.e+36f ;
	float TAUY(time, lndgrid) ;
		TAUY:long_name = "meridional surface stress" ;
		TAUY:units = "kg/m/s^2" ;
		TAUY:cell_methods = "time: mean" ;
		TAUY:_FillValue = 1.e+36f ;
		TAUY:missing_value = 1.e+36f ;
	float TBOT(time, lndgrid) ;
		TBOT:long_name = "atmospheric air temperature" ;
		TBOT:units = "K" ;
		TBOT:cell_methods = "time: mean" ;
		TBOT:_FillValue = 1.e+36f ;
		TBOT:missing_value = 1.e+36f ;
	float TBUILD(time, lndgrid) ;
		TBUILD:long_name = "internal urban building temperature" ;
		TBUILD:units = "K" ;
		TBUILD:cell_methods = "time: mean" ;
		TBUILD:_FillValue = 1.e+36f ;
		TBUILD:missing_value = 1.e+36f ;
	float TG(time, lndgrid) ;
		TG:long_name = "ground temperature" ;
		TG:units = "K" ;
		TG:cell_methods = "time: mean" ;
		TG:_FillValue = 1.e+36f ;
		TG:missing_value = 1.e+36f ;
	float TG_R(time, lndgrid) ;
		TG_R:long_name = "Rural ground temperature" ;
		TG_R:units = "K" ;
		TG_R:cell_methods = "time: mean" ;
		TG_R:_FillValue = 1.e+36f ;
		TG_R:missing_value = 1.e+36f ;
	float TG_U(time, lndgrid) ;
		TG_U:long_name = "Urban ground temperature" ;
		TG_U:units = "K" ;
		TG_U:cell_methods = "time: mean" ;
		TG_U:_FillValue = 1.e+36f ;
		TG_U:missing_value = 1.e+36f ;
	float TH2OSFC(time, lndgrid) ;
		TH2OSFC:long_name = "surface water temperature" ;
		TH2OSFC:units = "K" ;
		TH2OSFC:cell_methods = "time: mean" ;
		TH2OSFC:_FillValue = 1.e+36f ;
		TH2OSFC:missing_value = 1.e+36f ;
	float THBOT(time, lndgrid) ;
		THBOT:long_name = "atmospheric air potential temperature" ;
		THBOT:units = "K" ;
		THBOT:cell_methods = "time: mean" ;
		THBOT:_FillValue = 1.e+36f ;
		THBOT:missing_value = 1.e+36f ;
	float TKE1(time, lndgrid) ;
		TKE1:long_name = "top lake level eddy thermal conductivity" ;
		TKE1:units = "W/(mK)" ;
		TKE1:cell_methods = "time: mean" ;
		TKE1:_FillValue = 1.e+36f ;
		TKE1:missing_value = 1.e+36f ;
	float TLAI(time, lndgrid) ;
		TLAI:long_name = "total projected leaf area index" ;
		TLAI:units = "none" ;
		TLAI:cell_methods = "time: mean" ;
		TLAI:_FillValue = 1.e+36f ;
		TLAI:missing_value = 1.e+36f ;
	float TLAKE(time, levlak, lndgrid) ;
		TLAKE:long_name = "lake temperature" ;
		TLAKE:units = "K" ;
		TLAKE:cell_methods = "time: mean" ;
		TLAKE:_FillValue = 1.e+36f ;
		TLAKE:missing_value = 1.e+36f ;
	float TOTCOLC(time, lndgrid) ;
		TOTCOLC:long_name = "total column carbon, incl veg and cpool" ;
		TOTCOLC:units = "gC/m^2" ;
		TOTCOLC:cell_methods = "time: mean" ;
		TOTCOLC:_FillValue = 1.e+36f ;
		TOTCOLC:missing_value = 1.e+36f ;
	float TOTCOLCH4(time, lndgrid) ;
		TOTCOLCH4:long_name = "total belowground CH4, (0 for non-lake special landunits)" ;
		TOTCOLCH4:units = "gC/m2" ;
		TOTCOLCH4:cell_methods = "time: mean" ;
		TOTCOLCH4:_FillValue = 1.e+36f ;
		TOTCOLCH4:missing_value = 1.e+36f ;
	float TOTCOLN(time, lndgrid) ;
		TOTCOLN:long_name = "total column-level N" ;
		TOTCOLN:units = "gN/m^2" ;
		TOTCOLN:cell_methods = "time: mean" ;
		TOTCOLN:_FillValue = 1.e+36f ;
		TOTCOLN:missing_value = 1.e+36f ;
	float TOTECOSYSC(time, lndgrid) ;
		TOTECOSYSC:long_name = "total ecosystem carbon, incl veg but excl cpool" ;
		TOTECOSYSC:units = "gC/m^2" ;
		TOTECOSYSC:cell_methods = "time: mean" ;
		TOTECOSYSC:_FillValue = 1.e+36f ;
		TOTECOSYSC:missing_value = 1.e+36f ;
	float TOTECOSYSN(time, lndgrid) ;
		TOTECOSYSN:long_name = "total ecosystem N" ;
		TOTECOSYSN:units = "gN/m^2" ;
		TOTECOSYSN:cell_methods = "time: mean" ;
		TOTECOSYSN:_FillValue = 1.e+36f ;
		TOTECOSYSN:missing_value = 1.e+36f ;
	float TOTLITC(time, lndgrid) ;
		TOTLITC:long_name = "total litter carbon" ;
		TOTLITC:units = "gC/m^2" ;
		TOTLITC:cell_methods = "time: mean" ;
		TOTLITC:_FillValue = 1.e+36f ;
		TOTLITC:missing_value = 1.e+36f ;
	float TOTLITC_1m(time, lndgrid) ;
		TOTLITC_1m:long_name = "total litter carbon to 1 meter depth" ;
		TOTLITC_1m:units = "gC/m^2" ;
		TOTLITC_1m:cell_methods = "time: mean" ;
		TOTLITC_1m:_FillValue = 1.e+36f ;
		TOTLITC_1m:missing_value = 1.e+36f ;
	float TOTLITN(time, lndgrid) ;
		TOTLITN:long_name = "total litter N" ;
		TOTLITN:units = "gN/m^2" ;
		TOTLITN:cell_methods = "time: mean" ;
		TOTLITN:_FillValue = 1.e+36f ;
		TOTLITN:missing_value = 1.e+36f ;
	float TOTLITN_1m(time, lndgrid) ;
		TOTLITN_1m:long_name = "total litter N to 1 meter" ;
		TOTLITN_1m:units = "gN/m^2" ;
		TOTLITN_1m:cell_methods = "time: mean" ;
		TOTLITN_1m:_FillValue = 1.e+36f ;
		TOTLITN_1m:missing_value = 1.e+36f ;
	float TOTPFTC(time, lndgrid) ;
		TOTPFTC:long_name = "total pft-level carbon, including cpool" ;
		TOTPFTC:units = "gC/m^2" ;
		TOTPFTC:cell_methods = "time: mean" ;
		TOTPFTC:_FillValue = 1.e+36f ;
		TOTPFTC:missing_value = 1.e+36f ;
	float TOTPFTN(time, lndgrid) ;
		TOTPFTN:long_name = "total PFT-level nitrogen" ;
		TOTPFTN:units = "gN/m^2" ;
		TOTPFTN:cell_methods = "time: mean" ;
		TOTPFTN:_FillValue = 1.e+36f ;
		TOTPFTN:missing_value = 1.e+36f ;
	float TOTPRODC(time, lndgrid) ;
		TOTPRODC:long_name = "total wood product C" ;
		TOTPRODC:units = "gC/m^2" ;
		TOTPRODC:cell_methods = "time: mean" ;
		TOTPRODC:_FillValue = 1.e+36f ;
		TOTPRODC:missing_value = 1.e+36f ;
	float TOTPRODN(time, lndgrid) ;
		TOTPRODN:long_name = "total wood product N" ;
		TOTPRODN:units = "gN/m^2" ;
		TOTPRODN:cell_methods = "time: mean" ;
		TOTPRODN:_FillValue = 1.e+36f ;
		TOTPRODN:missing_value = 1.e+36f ;
	float TOTSOMC(time, lndgrid) ;
		TOTSOMC:long_name = "total soil organic matter carbon" ;
		TOTSOMC:units = "gC/m^2" ;
		TOTSOMC:cell_methods = "time: mean" ;
		TOTSOMC:_FillValue = 1.e+36f ;
		TOTSOMC:missing_value = 1.e+36f ;
	float TOTSOMC_1m(time, lndgrid) ;
		TOTSOMC_1m:long_name = "total soil organic matter carbon to 1 meter depth" ;
		TOTSOMC_1m:units = "gC/m^2" ;
		TOTSOMC_1m:cell_methods = "time: mean" ;
		TOTSOMC_1m:_FillValue = 1.e+36f ;
		TOTSOMC_1m:missing_value = 1.e+36f ;
	float TOTSOMN(time, lndgrid) ;
		TOTSOMN:long_name = "total soil organic matter N" ;
		TOTSOMN:units = "gN/m^2" ;
		TOTSOMN:cell_methods = "time: mean" ;
		TOTSOMN:_FillValue = 1.e+36f ;
		TOTSOMN:missing_value = 1.e+36f ;
	float TOTSOMN_1m(time, lndgrid) ;
		TOTSOMN_1m:long_name = "total soil organic matter N to 1 meter" ;
		TOTSOMN_1m:units = "gN/m^2" ;
		TOTSOMN_1m:cell_methods = "time: mean" ;
		TOTSOMN_1m:_FillValue = 1.e+36f ;
		TOTSOMN_1m:missing_value = 1.e+36f ;
	float TOTVEGC(time, lndgrid) ;
		TOTVEGC:long_name = "total vegetation carbon, excluding cpool" ;
		TOTVEGC:units = "gC/m^2" ;
		TOTVEGC:cell_methods = "time: mean" ;
		TOTVEGC:_FillValue = 1.e+36f ;
		TOTVEGC:missing_value = 1.e+36f ;
	float TOTVEGN(time, lndgrid) ;
		TOTVEGN:long_name = "total vegetation nitrogen" ;
		TOTVEGN:units = "gN/m^2" ;
		TOTVEGN:cell_methods = "time: mean" ;
		TOTVEGN:_FillValue = 1.e+36f ;
		TOTVEGN:missing_value = 1.e+36f ;
	float TREFMNAV(time, lndgrid) ;
		TREFMNAV:long_name = "daily minimum of average 2-m temperature" ;
		TREFMNAV:units = "K" ;
		TREFMNAV:cell_methods = "time: mean" ;
		TREFMNAV:_FillValue = 1.e+36f ;
		TREFMNAV:missing_value = 1.e+36f ;
	float TREFMNAV_R(time, lndgrid) ;
		TREFMNAV_R:long_name = "Rural daily minimum of average 2-m temperature" ;
		TREFMNAV_R:units = "K" ;
		TREFMNAV_R:cell_methods = "time: mean" ;
		TREFMNAV_R:_FillValue = 1.e+36f ;
		TREFMNAV_R:missing_value = 1.e+36f ;
	float TREFMNAV_U(time, lndgrid) ;
		TREFMNAV_U:long_name = "Urban daily minimum of average 2-m temperature" ;
		TREFMNAV_U:units = "K" ;
		TREFMNAV_U:cell_methods = "time: mean" ;
		TREFMNAV_U:_FillValue = 1.e+36f ;
		TREFMNAV_U:missing_value = 1.e+36f ;
	float TREFMXAV(time, lndgrid) ;
		TREFMXAV:long_name = "daily maximum of average 2-m temperature" ;
		TREFMXAV:units = "K" ;
		TREFMXAV:cell_methods = "time: mean" ;
		TREFMXAV:_FillValue = 1.e+36f ;
		TREFMXAV:missing_value = 1.e+36f ;
	float TREFMXAV_R(time, lndgrid) ;
		TREFMXAV_R:long_name = "Rural daily maximum of average 2-m temperature" ;
		TREFMXAV_R:units = "K" ;
		TREFMXAV_R:cell_methods = "time: mean" ;
		TREFMXAV_R:_FillValue = 1.e+36f ;
		TREFMXAV_R:missing_value = 1.e+36f ;
	float TREFMXAV_U(time, lndgrid) ;
		TREFMXAV_U:long_name = "Urban daily maximum of average 2-m temperature" ;
		TREFMXAV_U:units = "K" ;
		TREFMXAV_U:cell_methods = "time: mean" ;
		TREFMXAV_U:_FillValue = 1.e+36f ;
		TREFMXAV_U:missing_value = 1.e+36f ;
	float TSA(time, lndgrid) ;
		TSA:long_name = "2m air temperature" ;
		TSA:units = "K" ;
		TSA:cell_methods = "time: mean" ;
		TSA:_FillValue = 1.e+36f ;
		TSA:missing_value = 1.e+36f ;
	float TSAI(time, lndgrid) ;
		TSAI:long_name = "total projected stem area index" ;
		TSAI:units = "none" ;
		TSAI:cell_methods = "time: mean" ;
		TSAI:_FillValue = 1.e+36f ;
		TSAI:missing_value = 1.e+36f ;
	float TSA_R(time, lndgrid) ;
		TSA_R:long_name = "Rural 2m air temperature" ;
		TSA_R:units = "K" ;
		TSA_R:cell_methods = "time: mean" ;
		TSA_R:_FillValue = 1.e+36f ;
		TSA_R:missing_value = 1.e+36f ;
	float TSA_U(time, lndgrid) ;
		TSA_U:long_name = "Urban 2m air temperature" ;
		TSA_U:units = "K" ;
		TSA_U:cell_methods = "time: mean" ;
		TSA_U:_FillValue = 1.e+36f ;
		TSA_U:missing_value = 1.e+36f ;
	float TSOI(time, levgrnd, lndgrid) ;
		TSOI:long_name = "soil temperature (vegetated landunits only)" ;
		TSOI:units = "K" ;
		TSOI:cell_methods = "time: mean" ;
		TSOI:_FillValue = 1.e+36f ;
		TSOI:missing_value = 1.e+36f ;
	float TSOI_10CM(time, lndgrid) ;
		TSOI_10CM:long_name = "soil temperature in top 10cm of soil" ;
		TSOI_10CM:units = "K" ;
		TSOI_10CM:cell_methods = "time: mean" ;
		TSOI_10CM:_FillValue = 1.e+36f ;
		TSOI_10CM:missing_value = 1.e+36f ;
	float TSOI_ICE(time, levgrnd, lndgrid) ;
		TSOI_ICE:long_name = "soil temperature (ice landunits only)" ;
		TSOI_ICE:units = "K" ;
		TSOI_ICE:cell_methods = "time: mean" ;
		TSOI_ICE:_FillValue = 1.e+36f ;
		TSOI_ICE:missing_value = 1.e+36f ;
	float TV(time, lndgrid) ;
		TV:long_name = "vegetation temperature" ;
		TV:units = "K" ;
		TV:cell_methods = "time: mean" ;
		TV:_FillValue = 1.e+36f ;
		TV:missing_value = 1.e+36f ;
	float TWS(time, lndgrid) ;
		TWS:long_name = "total water storage" ;
		TWS:units = "mm" ;
		TWS:cell_methods = "time: mean" ;
		TWS:_FillValue = 1.e+36f ;
		TWS:missing_value = 1.e+36f ;
	float T_SCALAR(time, levdcmp, lndgrid) ;
		T_SCALAR:long_name = "temperature inhibition of decomposition" ;
		T_SCALAR:units = "unitless" ;
		T_SCALAR:cell_methods = "time: mean" ;
		T_SCALAR:_FillValue = 1.e+36f ;
		T_SCALAR:missing_value = 1.e+36f ;
	float U10(time, lndgrid) ;
		U10:long_name = "10-m wind" ;
		U10:units = "m/s" ;
		U10:cell_methods = "time: mean" ;
		U10:_FillValue = 1.e+36f ;
		U10:missing_value = 1.e+36f ;
	float URBAN_AC(time, lndgrid) ;
		URBAN_AC:long_name = "urban air conditioning flux" ;
		URBAN_AC:units = "W/m^2" ;
		URBAN_AC:cell_methods = "time: mean" ;
		URBAN_AC:_FillValue = 1.e+36f ;
		URBAN_AC:missing_value = 1.e+36f ;
	float URBAN_HEAT(time, lndgrid) ;
		URBAN_HEAT:long_name = "urban heating flux" ;
		URBAN_HEAT:units = "W/m^2" ;
		URBAN_HEAT:cell_methods = "time: mean" ;
		URBAN_HEAT:_FillValue = 1.e+36f ;
		URBAN_HEAT:missing_value = 1.e+36f ;
	float VOCFLXT(time, lndgrid) ;
		VOCFLXT:long_name = "total VOC flux into atmosphere" ;
		VOCFLXT:units = "moles/m2/sec" ;
		VOCFLXT:cell_methods = "time: mean" ;
		VOCFLXT:_FillValue = 1.e+36f ;
		VOCFLXT:missing_value = 1.e+36f ;
	float VOLR(time, lndgrid) ;
		VOLR:long_name = "river channel water storage" ;
		VOLR:units = "m3" ;
		VOLR:cell_methods = "time: mean" ;
		VOLR:_FillValue = 1.e+36f ;
		VOLR:missing_value = 1.e+36f ;
	float WA(time, lndgrid) ;
		WA:long_name = "water in the unconfined aquifer (vegetated landunits only)" ;
		WA:units = "mm" ;
		WA:cell_methods = "time: mean" ;
		WA:_FillValue = 1.e+36f ;
		WA:missing_value = 1.e+36f ;
	float WASTEHEAT(time, lndgrid) ;
		WASTEHEAT:long_name = "sensible heat flux from heating/cooling sources of urban waste heat" ;
		WASTEHEAT:units = "W/m^2" ;
		WASTEHEAT:cell_methods = "time: mean" ;
		WASTEHEAT:_FillValue = 1.e+36f ;
		WASTEHEAT:missing_value = 1.e+36f ;
	float WF(time, lndgrid) ;
		WF:long_name = "soil water as frac. of whc for top 0.05 m" ;
		WF:units = "proportion" ;
		WF:cell_methods = "time: mean" ;
		WF:_FillValue = 1.e+36f ;
		WF:missing_value = 1.e+36f ;
	float WIND(time, lndgrid) ;
		WIND:long_name = "atmospheric wind velocity magnitude" ;
		WIND:units = "m/s" ;
		WIND:cell_methods = "time: mean" ;
		WIND:_FillValue = 1.e+36f ;
		WIND:missing_value = 1.e+36f ;
	float WOODC(time, lndgrid) ;
		WOODC:long_name = "wood C" ;
		WOODC:units = "gC/m^2" ;
		WOODC:cell_methods = "time: mean" ;
		WOODC:_FillValue = 1.e+36f ;
		WOODC:missing_value = 1.e+36f ;
	float WOODC_ALLOC(time, lndgrid) ;
		WOODC_ALLOC:long_name = "wood C allocation" ;
		WOODC_ALLOC:units = "gC/m^2/s" ;
		WOODC_ALLOC:cell_methods = "time: mean" ;
		WOODC_ALLOC:_FillValue = 1.e+36f ;
		WOODC_ALLOC:missing_value = 1.e+36f ;
	float WOODC_LOSS(time, lndgrid) ;
		WOODC_LOSS:long_name = "wood C loss" ;
		WOODC_LOSS:units = "gC/m^2/s" ;
		WOODC_LOSS:cell_methods = "time: mean" ;
		WOODC_LOSS:_FillValue = 1.e+36f ;
		WOODC_LOSS:missing_value = 1.e+36f ;
	float WOOD_HARVESTC(time, lndgrid) ;
		WOOD_HARVESTC:long_name = "wood harvest carbon (to product pools)" ;
		WOOD_HARVESTC:units = "gC/m^2/s" ;
		WOOD_HARVESTC:cell_methods = "time: mean" ;
		WOOD_HARVESTC:_FillValue = 1.e+36f ;
		WOOD_HARVESTC:missing_value = 1.e+36f ;
	float WOOD_HARVESTN(time, lndgrid) ;
		WOOD_HARVESTN:long_name = "wood harvest N (to product pools)" ;
		WOOD_HARVESTN:units = "gN/m^2/s" ;
		WOOD_HARVESTN:cell_methods = "time: mean" ;
		WOOD_HARVESTN:_FillValue = 1.e+36f ;
		WOOD_HARVESTN:missing_value = 1.e+36f ;
	float WTGQ(time, lndgrid) ;
		WTGQ:long_name = "surface tracer conductance" ;
		WTGQ:units = "m/s" ;
		WTGQ:cell_methods = "time: mean" ;
		WTGQ:_FillValue = 1.e+36f ;
		WTGQ:missing_value = 1.e+36f ;
	float W_SCALAR(time, levdcmp, lndgrid) ;
		W_SCALAR:long_name = "Moisture (dryness) inhibition of decomposition" ;
		W_SCALAR:units = "unitless" ;
		W_SCALAR:cell_methods = "time: mean" ;
		W_SCALAR:_FillValue = 1.e+36f ;
		W_SCALAR:missing_value = 1.e+36f ;
	float XSMRPOOL(time, lndgrid) ;
		XSMRPOOL:long_name = "temporary photosynthate C pool" ;
		XSMRPOOL:units = "gC/m^2" ;
		XSMRPOOL:cell_methods = "time: mean" ;
		XSMRPOOL:_FillValue = 1.e+36f ;
		XSMRPOOL:missing_value = 1.e+36f ;
	float XSMRPOOL_RECOVER(time, lndgrid) ;
		XSMRPOOL_RECOVER:long_name = "C flux assigned to recovery of negative xsmrpool" ;
		XSMRPOOL_RECOVER:units = "gC/m^2/s" ;
		XSMRPOOL_RECOVER:cell_methods = "time: mean" ;
		XSMRPOOL_RECOVER:_FillValue = 1.e+36f ;
		XSMRPOOL_RECOVER:missing_value = 1.e+36f ;
	float ZBOT(time, lndgrid) ;
		ZBOT:long_name = "atmospheric reference height" ;
		ZBOT:units = "m" ;
		ZBOT:cell_methods = "time: mean" ;
		ZBOT:_FillValue = 1.e+36f ;
		ZBOT:missing_value = 1.e+36f ;
	float ZWT(time, lndgrid) ;
		ZWT:long_name = "water table depth (vegetated landunits only)" ;
		ZWT:units = "m" ;
		ZWT:cell_methods = "time: mean" ;
		ZWT:_FillValue = 1.e+36f ;
		ZWT:missing_value = 1.e+36f ;
	float ZWT_CH4_UNSAT(time, lndgrid) ;
		ZWT_CH4_UNSAT:long_name = "depth of water table for methane production used in non-inundated area" ;
		ZWT_CH4_UNSAT:units = "m" ;
		ZWT_CH4_UNSAT:cell_methods = "time: mean" ;
		ZWT_CH4_UNSAT:_FillValue = 1.e+36f ;
		ZWT_CH4_UNSAT:missing_value = 1.e+36f ;
	float ZWT_PERCH(time, lndgrid) ;
		ZWT_PERCH:long_name = "perched water table depth (vegetated landunits only)" ;
		ZWT_PERCH:units = "m" ;
		ZWT_PERCH:cell_methods = "time: mean" ;
		ZWT_PERCH:_FillValue = 1.e+36f ;
		ZWT_PERCH:missing_value = 1.e+36f ;
	float o2_decomp_depth_unsat(time, levgrnd, lndgrid) ;
		o2_decomp_depth_unsat:long_name = "o2_decomp_depth_unsat" ;
		o2_decomp_depth_unsat:units = "mol/m3/2" ;
		o2_decomp_depth_unsat:cell_methods = "time: mean" ;
		o2_decomp_depth_unsat:_FillValue = 1.e+36f ;
		o2_decomp_depth_unsat:missing_value = 1.e+36f ;

// global attributes:
		:title = "CLM History file information" ;
		:comment = "NOTE: None of the variables are weighted by land fraction!" ;
		:Conventions = "CF-1.0" ;
		:history = "created on 02/14/14 17:22:10" ;
		:source = "Community Land Model CLM4.0" ;
		:hostname = "userdefined" ;
		:username = "bandre" ;
		:version = "" ;
		:revision_id = "$Id: histFileMod.F90 42903 2012-12-21 15:32:10Z muszala $" ;
		:case_title = "UNSET" ;
		:case_id = "ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-1" ;
		:Surface_dataset = "surfdata_13x26pt_US-Brw_simyr1850.nc" ;
		:Initial_conditions_dataset = "arbitrary initialization" ;
		:PFT_physiological_constants_dataset = "clm_params.c130821.nc" ;
		:Time_constant_3Dvars_filename = "./ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-1.clm2.h0.0001-01-01-00000.nc" ;
		:Time_constant_3Dvars = "ZSOI:DZSOI:WATSAT:SUCSAT:BSW:HKSAT:ZLAKE:DZLAKE" ;
data:

 levgrnd = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 levlak = 0.05, 0.6, 2.1, 4.6, 8.1, 12.6, 18.6, 25.6, 34.325, 44.775 ;

 levdcmp = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 time = 1 ;

 mcdate = 10102 ;

 mcsec = 0 ;

 mdcur = 1 ;

 mscur = 0 ;

 nstep = 48 ;

 time_bounds =
  0, 1 ;

 date_written =
  "02/14/14" ;

 time_written =
  "17:22:10" ;

 lon = -156.6089, -156.6089, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6083, -156.6082, -156.608, -156.608, -156.6078, -156.6078, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, 
    -156.6069, -156.6069, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6063, -156.6062, -156.6089, -156.6089, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6083, -156.6082, -156.608, -156.608, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6074, -156.6073, 
    -156.6071, -156.6071, -156.6069, -156.6069, -156.6067, -156.6066, 
    -156.6065, -156.6064, -156.6063, -156.6062, -156.6089, -156.6089, 
    -156.6087, -156.6086, -156.6085, -156.6084, -156.6083, -156.6082, 
    -156.608, -156.608, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6074, -156.6073, -156.6071, -156.6071, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6065, -156.6064, -156.6062, -156.6062, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6082, -156.6082, -156.608, -156.608, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6071, -156.6071, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6062, -156.6062, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6082, -156.6082, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6073, -156.6073, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6067, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6062, -156.6089, -156.6088, 
    -156.6087, -156.6086, -156.6084, -156.6084, -156.6082, -156.6082, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6073, -156.6073, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6064, -156.6064, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6084, -156.6084, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6073, -156.6073, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6064, -156.6064, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6084, -156.6084, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6075, -156.6075, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6061, -156.6089, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6084, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6075, -156.6075, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6066, -156.6066, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6086, -156.6086, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6075, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6066, -156.6066, -156.6064, -156.6063, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6086, -156.6086, 
    -156.6084, -156.6083, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6077, -156.6077, -156.6075, -156.6074, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6068, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6063, -156.6062, -156.6061, -156.6088, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6083, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6077, -156.6077, -156.6075, -156.6074, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6068, -156.6068, 
    -156.6066, -156.6065, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6088, -156.6088, -156.6086, -156.6085, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.6079, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6068, -156.6068, -156.6066, -156.6065, -156.6064, -156.6063, 
    -156.6062, -156.6061 ;

 lat = 71.27904, 71.27901, 71.27903, 71.27901, 71.27901, 71.27903, 71.27901, 
    71.27903, 71.279, 71.27902, 71.27902, 71.279, 71.27899, 71.27901, 
    71.27901, 71.27899, 71.27899, 71.27901, 71.27898, 71.27901, 71.27901, 
    71.27898, 71.27901, 71.27898, 71.27898, 71.279, 71.27911, 71.27908, 
    71.27911, 71.27908, 71.27908, 71.2791, 71.27908, 71.2791, 71.2791, 
    71.27907, 71.27907, 71.27909, 71.27909, 71.27907, 71.27909, 71.27906, 
    71.27906, 71.27908, 71.27906, 71.27908, 71.27905, 71.27908, 71.27908, 
    71.27905, 71.27908, 71.27905, 71.27915, 71.27918, 71.27915, 71.27917, 
    71.27917, 71.27915, 71.27917, 71.27914, 71.27914, 71.27917, 71.27914, 
    71.27917, 71.27916, 71.27914, 71.27914, 71.27916, 71.27914, 71.27916, 
    71.27913, 71.27915, 71.27913, 71.27915, 71.27915, 71.27912, 71.27914, 
    71.27912, 71.27923, 71.27925, 71.27923, 71.27925, 71.27924, 71.27922, 
    71.27922, 71.27924, 71.27921, 71.27924, 71.27921, 71.27924, 71.27924, 
    71.27921, 71.27921, 71.27923, 71.27923, 71.27921, 71.27923, 71.2792, 
    71.27922, 71.2792, 71.27922, 71.2792, 71.27922, 71.27919, 71.27932, 
    71.2793, 71.2793, 71.27932, 71.2793, 71.27932, 71.27931, 71.27929, 
    71.27929, 71.27931, 71.27931, 71.27928, 71.27928, 71.2793, 71.27928, 
    71.2793, 71.27927, 71.2793, 71.27927, 71.2793, 71.2793, 71.27927, 
    71.27929, 71.27927, 71.27927, 71.27929, 71.27937, 71.2794, 71.27937, 
    71.27939, 71.27939, 71.27937, 71.27937, 71.27939, 71.27938, 71.27936, 
    71.27936, 71.27938, 71.27935, 71.27937, 71.27935, 71.27937, 71.27935, 
    71.27937, 71.27934, 71.27937, 71.27937, 71.27934, 71.27937, 71.27934, 
    71.27934, 71.27936, 71.27944, 71.27946, 71.27946, 71.27944, 71.27946, 
    71.27943, 71.27943, 71.27946, 71.27946, 71.27943, 71.27945, 71.27943, 
    71.27943, 71.27945, 71.27942, 71.27944, 71.27942, 71.27944, 71.27942, 
    71.27944, 71.27943, 71.27941, 71.27943, 71.27941, 71.27943, 71.2794, 
    71.27951, 71.27953, 71.27951, 71.27953, 71.27953, 71.27951, 71.2795, 
    71.27953, 71.27953, 71.2795, 71.27953, 71.2795, 71.2795, 71.27952, 
    71.2795, 71.27952, 71.27949, 71.27951, 71.27949, 71.27951, 71.27951, 
    71.27949, 71.27951, 71.27948, 71.27948, 71.2795, 71.27959, 71.27961, 
    71.27961, 71.27958, 71.2796, 71.27958, 71.27958, 71.2796, 71.2796, 
    71.27957, 71.27957, 71.27959, 71.27957, 71.27959, 71.27959, 71.27956, 
    71.27959, 71.27956, 71.27956, 71.27959, 71.27958, 71.27956, 71.27958, 
    71.27956, 71.27958, 71.27955, 71.27966, 71.27968, 71.27968, 71.27966, 
    71.27968, 71.27965, 71.27967, 71.27965, 71.27967, 71.27965, 71.27967, 
    71.27964, 71.27966, 71.27964, 71.27964, 71.27966, 71.27963, 71.27966, 
    71.27966, 71.27963, 71.27963, 71.27966, 71.27962, 71.27965, 71.27962, 
    71.27965, 71.27973, 71.27975, 71.27975, 71.27972, 71.27975, 71.27972, 
    71.27972, 71.27975, 71.27974, 71.27972, 71.27974, 71.27972, 71.27974, 
    71.27971, 71.27973, 71.27971, 71.27973, 71.27971, 71.27972, 71.2797, 
    71.2797, 71.27972, 71.27972, 71.27969, 71.27972, 71.27969, 71.27982, 
    71.2798, 71.2798, 71.27982, 71.27982, 71.27979, 71.27982, 71.27979, 
    71.27982, 71.27979, 71.27979, 71.27981, 71.27981, 71.27979, 71.27981, 
    71.27978, 71.2798, 71.27978, 71.27978, 71.2798, 71.27977, 71.27979, 
    71.27977, 71.27979, 71.27977, 71.27979, 71.2799, 71.27987, 71.27987, 
    71.27989, 71.27987, 71.27989, 71.27988, 71.27986, 71.27986, 71.27988, 
    71.27988, 71.27985, 71.27988, 71.27985, 71.27985, 71.27988, 71.27988, 
    71.27985, 71.27987, 71.27985, 71.27985, 71.27987, 71.27984, 71.27986, 
    71.27984, 71.27985 ;

 area = 9.902211e-05, 9.902174e-05, 9.902174e-05, 9.902209e-05, 9.902172e-05, 
    9.902208e-05, 9.902207e-05, 9.902169e-05, 9.902168e-05, 9.902204e-05, 
    9.902203e-05, 9.902166e-05, 9.902201e-05, 9.902164e-05, 9.902163e-05, 
    9.902199e-05, 9.902198e-05, 9.902161e-05, 9.902196e-05, 9.902159e-05, 
    9.902158e-05, 9.902194e-05, 9.902156e-05, 9.902192e-05, 9.902155e-05, 
    4.951087e-05, 9.902174e-05, 9.902138e-05, 9.902137e-05, 9.902173e-05, 
    9.902172e-05, 9.902135e-05, 9.90217e-05, 9.902133e-05, 9.902168e-05, 
    9.902132e-05, 9.90213e-05, 9.902166e-05, 9.902164e-05, 9.902128e-05, 
    9.902163e-05, 9.902126e-05, 9.902161e-05, 9.902124e-05, 9.902123e-05, 
    9.902159e-05, 9.902121e-05, 9.902157e-05, 9.902119e-05, 9.902156e-05, 
    9.902118e-05, 9.902155e-05, 9.902102e-05, 9.902138e-05, 9.902137e-05, 
    9.9021e-05, 9.902135e-05, 9.902099e-05, 9.902097e-05, 9.902133e-05, 
    9.902132e-05, 9.902095e-05, 9.90213e-05, 9.902093e-05, 9.902128e-05, 
    9.902092e-05, 9.902126e-05, 9.90209e-05, 9.902124e-05, 9.902088e-05, 
    9.902123e-05, 9.902086e-05, 9.902084e-05, 9.902121e-05, 9.902119e-05, 
    9.902083e-05, 9.902118e-05, 9.902081e-05, 9.902065e-05, 9.902102e-05, 
    9.9021e-05, 9.902064e-05, 9.902099e-05, 9.902062e-05, 9.902097e-05, 
    9.90206e-05, 9.902095e-05, 9.902059e-05, 9.902094e-05, 9.902057e-05, 
    9.902092e-05, 9.902055e-05, 9.902054e-05, 9.90209e-05, 9.902052e-05, 
    9.902088e-05, 9.902086e-05, 9.90205e-05, 9.902048e-05, 9.902084e-05, 
    9.902046e-05, 9.902083e-05, 9.902046e-05, 9.902081e-05, 9.902029e-05, 
    9.902065e-05, 9.902064e-05, 9.902028e-05, 9.902062e-05, 9.902026e-05, 
    9.902024e-05, 9.90206e-05, 9.902059e-05, 9.902022e-05, 9.90202e-05, 
    9.902057e-05, 9.902019e-05, 9.902055e-05, 9.902054e-05, 9.902017e-05, 
    9.902052e-05, 9.902015e-05, 9.902014e-05, 9.90205e-05, 9.902048e-05, 
    9.902012e-05, 9.902046e-05, 9.90201e-05, 9.902046e-05, 9.902009e-05, 
    9.901992e-05, 9.902028e-05, 9.901991e-05, 9.902028e-05, 9.902026e-05, 
    9.901989e-05, 9.901988e-05, 9.902024e-05, 9.902022e-05, 9.901986e-05, 
    9.90202e-05, 9.901984e-05, 9.901982e-05, 9.902019e-05, 9.90198e-05, 
    9.902017e-05, 9.901979e-05, 9.902015e-05, 9.901977e-05, 9.902013e-05, 
    9.902012e-05, 9.901975e-05, 9.90201e-05, 9.901973e-05, 9.901972e-05, 
    9.902009e-05, 9.901955e-05, 9.901992e-05, 9.901991e-05, 9.901955e-05, 
    9.90199e-05, 9.901953e-05, 9.901951e-05, 9.901988e-05, 9.901986e-05, 
    9.901949e-05, 9.901984e-05, 9.901947e-05, 9.901946e-05, 9.901982e-05, 
    9.901944e-05, 9.90198e-05, 9.901942e-05, 9.901979e-05, 9.90194e-05, 
    9.901977e-05, 9.901975e-05, 9.901939e-05, 9.901974e-05, 9.901937e-05, 
    9.901972e-05, 9.901936e-05, 9.901919e-05, 9.901955e-05, 9.901918e-05, 
    9.901955e-05, 9.901953e-05, 9.901916e-05, 9.901915e-05, 9.901951e-05, 
    9.90195e-05, 9.901913e-05, 9.901911e-05, 9.901947e-05, 9.90191e-05, 
    9.901946e-05, 9.901907e-05, 9.901944e-05, 9.901906e-05, 9.901942e-05, 
    9.901904e-05, 9.90194e-05, 9.901939e-05, 9.901902e-05, 9.901937e-05, 
    9.9019e-05, 9.901899e-05, 9.901936e-05, 9.901919e-05, 9.901883e-05, 
    9.901882e-05, 9.901918e-05, 9.90188e-05, 9.901916e-05, 9.901915e-05, 
    9.901878e-05, 9.901877e-05, 9.901913e-05, 9.901911e-05, 9.901875e-05, 
    9.901873e-05, 9.90191e-05, 9.901871e-05, 9.901907e-05, 9.90187e-05, 
    9.901906e-05, 9.901867e-05, 9.901904e-05, 9.901902e-05, 9.901866e-05, 
    9.901901e-05, 9.901864e-05, 9.901863e-05, 9.901899e-05, 9.901846e-05, 
    9.901883e-05, 9.901846e-05, 9.901882e-05, 9.90188e-05, 9.901843e-05, 
    9.901842e-05, 9.901878e-05, 9.90184e-05, 9.901876e-05, 9.901838e-05, 
    9.901875e-05, 9.901873e-05, 9.901836e-05, 9.901835e-05, 9.901871e-05, 
    9.90187e-05, 9.901833e-05, 9.901867e-05, 9.901831e-05, 9.901866e-05, 
    9.90183e-05, 9.901864e-05, 9.901827e-05, 9.901863e-05, 9.901827e-05, 
    9.90181e-05, 9.901846e-05, 9.901809e-05, 9.901846e-05, 9.901843e-05, 
    9.901807e-05, 9.901842e-05, 9.901806e-05, 9.901803e-05, 9.90184e-05, 
    9.901802e-05, 9.901838e-05, 9.901837e-05, 9.9018e-05, 9.901798e-05, 
    9.901835e-05, 9.901797e-05, 9.901833e-05, 9.901795e-05, 9.901831e-05, 
    9.901793e-05, 9.90183e-05, 9.901827e-05, 9.901791e-05, 9.901827e-05, 
    9.90179e-05, 9.90181e-05, 9.901774e-05, 9.901809e-05, 9.901772e-05, 
    9.901771e-05, 9.901807e-05, 9.901769e-05, 9.901806e-05, 9.901803e-05, 
    9.901767e-05, 9.901766e-05, 9.901802e-05, 9.9018e-05, 9.901763e-05, 
    9.901798e-05, 9.901762e-05, 9.90176e-05, 9.901796e-05, 9.901758e-05, 
    9.901795e-05, 9.901757e-05, 9.901793e-05, 9.901791e-05, 9.901755e-05, 
    9.90179e-05, 9.901754e-05, 9.901774e-05, 9.901737e-05, 9.901773e-05, 
    9.901736e-05, 9.901734e-05, 9.901771e-05, 9.901733e-05, 9.901768e-05, 
    9.901731e-05, 9.901767e-05, 9.901766e-05, 9.901728e-05, 9.901727e-05, 
    9.901763e-05, 9.901762e-05, 9.901726e-05, 9.901723e-05, 9.90176e-05, 
    9.901722e-05, 9.901758e-05, 9.901757e-05, 9.90172e-05, 9.901755e-05, 
    9.901718e-05, 9.901718e-05, 9.901754e-05 ;

 topo = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0 ;

 landfrac = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 landmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 pftmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 ACTUAL_IMMOB =
  4.718843e-14, 4.731617e-14, 4.729135e-14, 4.739429e-14, 4.733722e-14, 
    4.740459e-14, 4.721436e-14, 4.732122e-14, 4.725302e-14, 4.719996e-14, 
    4.759375e-14, 4.739888e-14, 4.779601e-14, 4.767194e-14, 4.798338e-14, 
    4.777668e-14, 4.802502e-14, 4.797746e-14, 4.812065e-14, 4.807965e-14, 
    4.826253e-14, 4.813958e-14, 4.835728e-14, 4.82332e-14, 4.82526e-14, 
    4.813551e-14, 4.743816e-14, 4.75695e-14, 4.743037e-14, 4.744911e-14, 
    4.744071e-14, 4.733838e-14, 4.728676e-14, 4.717869e-14, 4.719832e-14, 
    4.727771e-14, 4.745753e-14, 4.739655e-14, 4.755027e-14, 4.754681e-14, 
    4.77177e-14, 4.764068e-14, 4.792754e-14, 4.784611e-14, 4.808136e-14, 
    4.802223e-14, 4.807858e-14, 4.80615e-14, 4.80788e-14, 4.799207e-14, 
    4.802923e-14, 4.79529e-14, 4.76551e-14, 4.774269e-14, 4.748123e-14, 
    4.732369e-14, 4.721904e-14, 4.714469e-14, 4.715521e-14, 4.717524e-14, 
    4.727817e-14, 4.737491e-14, 4.744856e-14, 4.74978e-14, 4.754631e-14, 
    4.76929e-14, 4.77705e-14, 4.794399e-14, 4.791273e-14, 4.796571e-14, 
    4.801635e-14, 4.810127e-14, 4.80873e-14, 4.81247e-14, 4.796434e-14, 
    4.807092e-14, 4.789491e-14, 4.794307e-14, 4.755935e-14, 4.741301e-14, 
    4.735064e-14, 4.729612e-14, 4.716329e-14, 4.725503e-14, 4.721886e-14, 
    4.730491e-14, 4.735953e-14, 4.733252e-14, 4.749915e-14, 4.743439e-14, 
    4.77751e-14, 4.762847e-14, 4.801044e-14, 4.791915e-14, 4.803232e-14, 
    4.797459e-14, 4.807348e-14, 4.798448e-14, 4.813862e-14, 4.817214e-14, 
    4.814923e-14, 4.823726e-14, 4.797954e-14, 4.807857e-14, 4.733176e-14, 
    4.733616e-14, 4.735669e-14, 4.726641e-14, 4.726089e-14, 4.717814e-14, 
    4.725179e-14, 4.728313e-14, 4.73627e-14, 4.740972e-14, 4.745441e-14, 
    4.755261e-14, 4.766216e-14, 4.781523e-14, 4.792507e-14, 4.799865e-14, 
    4.795354e-14, 4.799337e-14, 4.794884e-14, 4.792798e-14, 4.815957e-14, 
    4.802957e-14, 4.82246e-14, 4.821382e-14, 4.812558e-14, 4.821504e-14, 
    4.733926e-14, 4.731391e-14, 4.722581e-14, 4.729476e-14, 4.716913e-14, 
    4.723945e-14, 4.727985e-14, 4.743571e-14, 4.746996e-14, 4.750167e-14, 
    4.756431e-14, 4.764462e-14, 4.778537e-14, 4.79077e-14, 4.80193e-14, 
    4.801113e-14, 4.801401e-14, 4.803891e-14, 4.797719e-14, 4.804904e-14, 
    4.806108e-14, 4.802957e-14, 4.821238e-14, 4.816018e-14, 4.821359e-14, 
    4.817961e-14, 4.732215e-14, 4.736481e-14, 4.734176e-14, 4.738509e-14, 
    4.735455e-14, 4.749024e-14, 4.753089e-14, 4.772097e-14, 4.764303e-14, 
    4.776708e-14, 4.765565e-14, 4.76754e-14, 4.777107e-14, 4.766168e-14, 
    4.790093e-14, 4.773873e-14, 4.803988e-14, 4.787804e-14, 4.805001e-14, 
    4.801882e-14, 4.807047e-14, 4.81167e-14, 4.817485e-14, 4.828204e-14, 
    4.825723e-14, 4.834684e-14, 4.742838e-14, 4.748364e-14, 4.74788e-14, 
    4.753663e-14, 4.757937e-14, 4.767199e-14, 4.782037e-14, 4.77646e-14, 
    4.786698e-14, 4.788749e-14, 4.773198e-14, 4.782748e-14, 4.752063e-14, 
    4.757023e-14, 4.754072e-14, 4.743272e-14, 4.777742e-14, 4.760063e-14, 
    4.792688e-14, 4.783129e-14, 4.81101e-14, 4.797148e-14, 4.824357e-14, 
    4.835962e-14, 4.846886e-14, 4.859624e-14, 4.751382e-14, 4.747628e-14, 
    4.754351e-14, 4.763642e-14, 4.772264e-14, 4.783712e-14, 4.784884e-14, 
    4.787026e-14, 4.792575e-14, 4.797239e-14, 4.787701e-14, 4.798408e-14, 
    4.758168e-14, 4.779276e-14, 4.746206e-14, 4.75617e-14, 4.763096e-14, 
    4.760061e-14, 4.775823e-14, 4.779534e-14, 4.794599e-14, 4.786817e-14, 
    4.833096e-14, 4.812642e-14, 4.869322e-14, 4.853509e-14, 4.746315e-14, 
    4.75137e-14, 4.768943e-14, 4.760585e-14, 4.784477e-14, 4.790347e-14, 
    4.795121e-14, 4.801216e-14, 4.801876e-14, 4.805486e-14, 4.79957e-14, 
    4.805254e-14, 4.783736e-14, 4.793356e-14, 4.766938e-14, 4.773373e-14, 
    4.770414e-14, 4.767166e-14, 4.777188e-14, 4.787851e-14, 4.788083e-14, 
    4.791497e-14, 4.801111e-14, 4.784574e-14, 4.835726e-14, 4.804153e-14, 
    4.75688e-14, 4.7666e-14, 4.767993e-14, 4.764228e-14, 4.789758e-14, 
    4.780515e-14, 4.805399e-14, 4.798679e-14, 4.809689e-14, 4.804219e-14, 
    4.803414e-14, 4.796385e-14, 4.792006e-14, 4.780938e-14, 4.771925e-14, 
    4.764775e-14, 4.766438e-14, 4.774291e-14, 4.788504e-14, 4.801934e-14, 
    4.798992e-14, 4.808852e-14, 4.782746e-14, 4.793696e-14, 4.789463e-14, 
    4.800499e-14, 4.776311e-14, 4.796898e-14, 4.771041e-14, 4.773311e-14, 
    4.780331e-14, 4.794436e-14, 4.797561e-14, 4.800889e-14, 4.798837e-14, 
    4.788862e-14, 4.787232e-14, 4.780162e-14, 4.778207e-14, 4.772817e-14, 
    4.768351e-14, 4.772431e-14, 4.776713e-14, 4.788868e-14, 4.799812e-14, 
    4.811735e-14, 4.814652e-14, 4.828552e-14, 4.817232e-14, 4.8359e-14, 
    4.820022e-14, 4.847499e-14, 4.798096e-14, 4.819564e-14, 4.780652e-14, 
    4.784852e-14, 4.792437e-14, 4.809829e-14, 4.800447e-14, 4.811421e-14, 
    4.787169e-14, 4.77456e-14, 4.771301e-14, 4.765209e-14, 4.77144e-14, 
    4.770933e-14, 4.776893e-14, 4.774978e-14, 4.789272e-14, 4.781598e-14, 
    4.803392e-14, 4.811335e-14, 4.833744e-14, 4.847456e-14, 4.861405e-14, 
    4.867555e-14, 4.869427e-14, 4.870209e-14 ;

 AGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX_LASTYEAR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 AR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_CROP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_PEATF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BCDEP =
  8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 8.212629e-15, 
    8.212629e-15, 8.212629e-15, 8.212629e-15 ;

 BGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BTRAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BUILDHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4PROD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_DIFF_SAT =
  -1.764688e-14, -1.766985e-14, -1.766537e-14, -1.76839e-14, -1.76736e-14, 
    -1.768575e-14, -1.765151e-14, -1.767078e-14, -1.765847e-14, 
    -1.764891e-14, -1.771985e-14, -1.768472e-14, -1.775594e-14, 
    -1.773367e-14, -1.778942e-14, -1.775251e-14, -1.779683e-14, 
    -1.778829e-14, -1.781381e-14, -1.78065e-14, -1.783921e-14, -1.781718e-14, 
    -1.785601e-14, -1.783392e-14, -1.78374e-14, -1.781646e-14, -1.769174e-14, 
    -1.771551e-14, -1.769034e-14, -1.769373e-14, -1.76922e-14, -1.767384e-14, 
    -1.766462e-14, -1.764508e-14, -1.764862e-14, -1.766294e-14, 
    -1.769526e-14, -1.768426e-14, -1.771183e-14, -1.771121e-14, 
    -1.774186e-14, -1.772805e-14, -1.777938e-14, -1.77648e-14, -1.780681e-14, 
    -1.779627e-14, -1.780632e-14, -1.780327e-14, -1.780636e-14, -1.77909e-14, 
    -1.779753e-14, -1.77839e-14, -1.773065e-14, -1.774635e-14, -1.769949e-14, 
    -1.76713e-14, -1.765237e-14, -1.763897e-14, -1.764086e-14, -1.764449e-14, 
    -1.766303e-14, -1.768037e-14, -1.769358e-14, -1.770242e-14, 
    -1.771112e-14, -1.773756e-14, -1.775137e-14, -1.778235e-14, 
    -1.777672e-14, -1.778622e-14, -1.779522e-14, -1.781038e-14, 
    -1.780787e-14, -1.781456e-14, -1.778593e-14, -1.780499e-14, 
    -1.777351e-14, -1.778214e-14, -1.77137e-14, -1.768721e-14, -1.767613e-14, 
    -1.766624e-14, -1.764233e-14, -1.765886e-14, -1.765235e-14, 
    -1.766778e-14, -1.767761e-14, -1.767274e-14, -1.770267e-14, 
    -1.769105e-14, -1.775219e-14, -1.77259e-14, -1.779417e-14, -1.777787e-14, 
    -1.779806e-14, -1.778775e-14, -1.780543e-14, -1.778952e-14, 
    -1.781703e-14, -1.782303e-14, -1.781894e-14, -1.783459e-14, 
    -1.778864e-14, -1.780634e-14, -1.767261e-14, -1.767341e-14, 
    -1.767709e-14, -1.766091e-14, -1.765991e-14, -1.764499e-14, 
    -1.765824e-14, -1.76639e-14, -1.767816e-14, -1.768663e-14, -1.769465e-14, 
    -1.771227e-14, -1.773195e-14, -1.775933e-14, -1.777893e-14, 
    -1.779205e-14, -1.778399e-14, -1.779111e-14, -1.778316e-14, 
    -1.777942e-14, -1.78208e-14, -1.779761e-14, -1.783234e-14, -1.783042e-14, 
    -1.781473e-14, -1.783063e-14, -1.767396e-14, -1.766939e-14, 
    -1.765358e-14, -1.766596e-14, -1.764336e-14, -1.765604e-14, 
    -1.766335e-14, -1.769134e-14, -1.769743e-14, -1.770314e-14, 
    -1.771436e-14, -1.772876e-14, -1.775399e-14, -1.777585e-14, 
    -1.779573e-14, -1.779427e-14, -1.779479e-14, -1.779925e-14, 
    -1.778823e-14, -1.780105e-14, -1.780322e-14, -1.779758e-14, 
    -1.783016e-14, -1.782086e-14, -1.783038e-14, -1.782432e-14, 
    -1.767087e-14, -1.767855e-14, -1.767441e-14, -1.768221e-14, 
    -1.767673e-14, -1.770114e-14, -1.770845e-14, -1.774251e-14, 
    -1.772849e-14, -1.775073e-14, -1.773073e-14, -1.773429e-14, 
    -1.775155e-14, -1.77318e-14, -1.777469e-14, -1.774571e-14, -1.779942e-14, 
    -1.777065e-14, -1.780122e-14, -1.779565e-14, -1.780486e-14, 
    -1.781313e-14, -1.782348e-14, -1.784261e-14, -1.783818e-14, 
    -1.785412e-14, -1.768997e-14, -1.769993e-14, -1.769901e-14, 
    -1.770939e-14, -1.771708e-14, -1.773365e-14, -1.776022e-14, 
    -1.775023e-14, -1.776853e-14, -1.777221e-14, -1.774438e-14, 
    -1.776152e-14, -1.770656e-14, -1.77155e-14, -1.771015e-14, -1.769078e-14, 
    -1.775259e-14, -1.772095e-14, -1.777926e-14, -1.776217e-14, 
    -1.781195e-14, -1.778727e-14, -1.783574e-14, -1.78565e-14, -1.78758e-14, 
    -1.789852e-14, -1.770531e-14, -1.769856e-14, -1.771062e-14, 
    -1.772735e-14, -1.774274e-14, -1.776322e-14, -1.776529e-14, 
    -1.776913e-14, -1.777903e-14, -1.778736e-14, -1.777039e-14, 
    -1.778945e-14, -1.771766e-14, -1.775531e-14, -1.769604e-14, 
    -1.771398e-14, -1.772635e-14, -1.772088e-14, -1.774907e-14, 
    -1.775572e-14, -1.77827e-14, -1.776874e-14, -1.785142e-14, -1.781493e-14, 
    -1.791565e-14, -1.788764e-14, -1.76962e-14, -1.770527e-14, -1.773682e-14, 
    -1.772182e-14, -1.776456e-14, -1.777507e-14, -1.778357e-14, -1.77945e-14, 
    -1.779564e-14, -1.78021e-14, -1.779152e-14, -1.780167e-14, -1.776326e-14, 
    -1.778044e-14, -1.773317e-14, -1.774472e-14, -1.77394e-14, -1.773358e-14, 
    -1.775152e-14, -1.777066e-14, -1.777101e-14, -1.777715e-14, 
    -1.779456e-14, -1.776473e-14, -1.785624e-14, -1.779995e-14, 
    -1.771515e-14, -1.773267e-14, -1.773509e-14, -1.772832e-14, 
    -1.777402e-14, -1.77575e-14, -1.780194e-14, -1.778993e-14, -1.780958e-14, 
    -1.779982e-14, -1.779839e-14, -1.778584e-14, -1.777803e-14, 
    -1.775827e-14, -1.774214e-14, -1.772929e-14, -1.773228e-14, 
    -1.774638e-14, -1.777182e-14, -1.779578e-14, -1.779054e-14, 
    -1.780808e-14, -1.776147e-14, -1.778108e-14, -1.777353e-14, 
    -1.779319e-14, -1.774998e-14, -1.778699e-14, -1.774052e-14, 
    -1.774459e-14, -1.775717e-14, -1.778245e-14, -1.778794e-14, 
    -1.779391e-14, -1.779021e-14, -1.777245e-14, -1.776951e-14, 
    -1.775684e-14, -1.775338e-14, -1.77437e-14, -1.77357e-14, -1.774302e-14, 
    -1.775072e-14, -1.777243e-14, -1.779199e-14, -1.781326e-14, 
    -1.781842e-14, -1.784336e-14, -1.782316e-14, -1.785656e-14, 
    -1.782831e-14, -1.787709e-14, -1.778904e-14, -1.782734e-14, 
    -1.775772e-14, -1.776522e-14, -1.777887e-14, -1.780993e-14, -1.77931e-14, 
    -1.781275e-14, -1.776939e-14, -1.77469e-14, -1.774099e-14, -1.773009e-14, 
    -1.774124e-14, -1.774033e-14, -1.775099e-14, -1.774756e-14, 
    -1.777315e-14, -1.775941e-14, -1.779837e-14, -1.781257e-14, 
    -1.785247e-14, -1.787689e-14, -1.790157e-14, -1.791248e-14, -1.79158e-14, 
    -1.791718e-14 ;

 CH4_SURF_DIFF_UNSAT =
  1.391905e-11, 1.379071e-11, 1.381577e-11, 1.371146e-11, 1.376944e-11, 
    1.370097e-11, 1.389314e-11, 1.378559e-11, 1.385436e-11, 1.390755e-11, 
    1.350647e-11, 1.370679e-11, 1.321951e-11, 1.333741e-11, 1.303696e-11, 
    1.323801e-11, 1.299567e-11, 1.304284e-11, 1.289988e-11, 1.294113e-11, 
    1.275513e-11, 1.288076e-11, 1.26569e-11, 1.278532e-11, 1.276537e-11, 
    1.288487e-11, 1.366673e-11, 1.353159e-11, 1.367469e-11, 1.365552e-11, 
    1.366413e-11, 1.376824e-11, 1.382037e-11, 1.392879e-11, 1.390919e-11, 
    1.382951e-11, 1.364689e-11, 1.370919e-11, 1.355157e-11, 1.355516e-11, 
    1.329422e-11, 1.336675e-11, 1.309195e-11, 1.317128e-11, 1.293942e-11, 
    1.299848e-11, 1.29422e-11, 1.295931e-11, 1.294198e-11, 1.30284e-11, 
    1.29915e-11, 1.306706e-11, 1.335323e-11, 1.327048e-11, 1.362262e-11, 
    1.378306e-11, 1.388844e-11, 1.396265e-11, 1.395219e-11, 1.393222e-11, 
    1.382905e-11, 1.373121e-11, 1.365611e-11, 1.360562e-11, 1.355567e-11, 
    1.331761e-11, 1.324394e-11, 1.307579e-11, 1.310646e-11, 1.305442e-11, 
    1.300433e-11, 1.29194e-11, 1.293345e-11, 1.289578e-11, 1.30558e-11, 
    1.294986e-11, 1.312386e-11, 1.307672e-11, 1.354207e-11, 1.369242e-11, 
    1.375578e-11, 1.381096e-11, 1.394414e-11, 1.385233e-11, 1.388861e-11, 
    1.380211e-11, 1.374682e-11, 1.37742e-11, 1.360424e-11, 1.367059e-11, 
    1.323954e-11, 1.337814e-11, 1.301019e-11, 1.310018e-11, 1.298844e-11, 
    1.304569e-11, 1.294731e-11, 1.303591e-11, 1.288171e-11, 1.284769e-11, 
    1.287096e-11, 1.278118e-11, 1.304079e-11, 1.29422e-11, 1.377497e-11, 
    1.377051e-11, 1.37497e-11, 1.384088e-11, 1.384643e-11, 1.392933e-11, 
    1.38556e-11, 1.382406e-11, 1.374361e-11, 1.369577e-11, 1.365012e-11, 
    1.354915e-11, 1.334659e-11, 1.320106e-11, 1.309438e-11, 1.302189e-11, 
    1.306643e-11, 1.302712e-11, 1.307105e-11, 1.309154e-11, 1.286046e-11, 
    1.299116e-11, 1.279416e-11, 1.28052e-11, 1.289488e-11, 1.280396e-11, 
    1.376737e-11, 1.379303e-11, 1.388166e-11, 1.381235e-11, 1.393832e-11, 
    1.386798e-11, 1.382734e-11, 1.366921e-11, 1.363419e-11, 1.360163e-11, 
    1.353707e-11, 1.336306e-11, 1.322973e-11, 1.311136e-11, 1.30014e-11, 
    1.300952e-11, 1.300666e-11, 1.298187e-11, 1.304311e-11, 1.297177e-11, 
    1.295972e-11, 1.299117e-11, 1.280668e-11, 1.285987e-11, 1.280544e-11, 
    1.284011e-11, 1.378469e-11, 1.374147e-11, 1.376484e-11, 1.372085e-11, 
    1.375186e-11, 1.361335e-11, 1.357152e-11, 1.329109e-11, 1.336454e-11, 
    1.324722e-11, 1.335272e-11, 1.333416e-11, 1.324336e-11, 1.334707e-11, 
    1.311795e-11, 1.327421e-11, 1.298091e-11, 1.314024e-11, 1.29708e-11, 
    1.300188e-11, 1.295034e-11, 1.290386e-11, 1.284496e-11, 1.273504e-11, 
    1.276064e-11, 1.266782e-11, 1.367674e-11, 1.362014e-11, 1.362513e-11, 
    1.356565e-11, 1.352148e-11, 1.333738e-11, 1.319612e-11, 1.324962e-11, 
    1.315105e-11, 1.313108e-11, 1.328069e-11, 1.318925e-11, 1.358212e-11, 
    1.35309e-11, 1.356142e-11, 1.367228e-11, 1.323733e-11, 1.349942e-11, 
    1.30926e-11, 1.318559e-11, 1.291051e-11, 1.304872e-11, 1.277469e-11, 
    1.265443e-11, 1.25396e-11, 1.240352e-11, 1.358914e-11, 1.362772e-11, 
    1.355856e-11, 1.337069e-11, 1.328954e-11, 1.317996e-11, 1.316864e-11, 
    1.314786e-11, 1.309372e-11, 1.304786e-11, 1.314128e-11, 1.303631e-11, 
    1.351899e-11, 1.322265e-11, 1.364228e-11, 1.353971e-11, 1.337581e-11, 
    1.349947e-11, 1.32557e-11, 1.32202e-11, 1.307383e-11, 1.314991e-11, 
    1.268428e-11, 1.289401e-11, 1.229859e-11, 1.24691e-11, 1.364117e-11, 
    1.358927e-11, 1.332093e-11, 1.349403e-11, 1.317258e-11, 1.31155e-11, 
    1.306873e-11, 1.300847e-11, 1.300193e-11, 1.296594e-11, 1.302482e-11, 
    1.296827e-11, 1.317973e-11, 1.308606e-11, 1.333983e-11, 1.327902e-11, 
    1.330707e-11, 1.333769e-11, 1.324267e-11, 1.313982e-11, 1.31376e-11, 
    1.310425e-11, 1.300939e-11, 1.317164e-11, 1.26568e-11, 1.297914e-11, 
    1.353243e-11, 1.334296e-11, 1.33299e-11, 1.336525e-11, 1.312125e-11, 
    1.321077e-11, 1.296682e-11, 1.303363e-11, 1.292382e-11, 1.297861e-11, 
    1.298663e-11, 1.305628e-11, 1.309929e-11, 1.320669e-11, 1.329275e-11, 
    1.336014e-11, 1.334454e-11, 1.327028e-11, 1.313347e-11, 1.300134e-11, 
    1.303051e-11, 1.293223e-11, 1.318929e-11, 1.30827e-11, 1.312411e-11, 
    1.30156e-11, 1.325104e-11, 1.30511e-11, 1.330114e-11, 1.327961e-11, 
    1.321253e-11, 1.307541e-11, 1.304468e-11, 1.301172e-11, 1.303207e-11, 
    1.312996e-11, 1.314586e-11, 1.321417e-11, 1.32329e-11, 1.328431e-11, 
    1.332654e-11, 1.328796e-11, 1.324719e-11, 1.312992e-11, 1.302239e-11, 
    1.29032e-11, 1.287372e-11, 1.273137e-11, 1.284746e-11, 1.265497e-11, 
    1.281893e-11, 1.253299e-11, 1.303932e-11, 1.282369e-11, 1.320946e-11, 
    1.316895e-11, 1.309504e-11, 1.292235e-11, 1.301612e-11, 1.290633e-11, 
    1.314648e-11, 1.32677e-11, 1.329868e-11, 1.335606e-11, 1.329736e-11, 
    1.330216e-11, 1.324549e-11, 1.326376e-11, 1.312599e-11, 1.320037e-11, 
    1.298683e-11, 1.290721e-11, 1.26776e-11, 1.253351e-11, 1.23844e-11, 
    1.231782e-11, 1.229747e-11, 1.228895e-11 ;

 CH4_SURF_EBUL_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_EBUL_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_CTRUNC =
  2.007731e-23, 2.007729e-23, 2.00773e-23, 2.007729e-23, 2.007729e-23, 
    2.007729e-23, 2.00773e-23, 2.007729e-23, 2.00773e-23, 2.00773e-23, 
    2.007727e-23, 2.007729e-23, 2.007726e-23, 2.007727e-23, 2.007724e-23, 
    2.007726e-23, 2.007724e-23, 2.007724e-23, 2.007723e-23, 2.007723e-23, 
    2.007722e-23, 2.007723e-23, 2.007721e-23, 2.007722e-23, 2.007722e-23, 
    2.007723e-23, 2.007728e-23, 2.007728e-23, 2.007729e-23, 2.007728e-23, 
    2.007728e-23, 2.007729e-23, 2.00773e-23, 2.007731e-23, 2.00773e-23, 
    2.00773e-23, 2.007728e-23, 2.007729e-23, 2.007728e-23, 2.007728e-23, 
    2.007726e-23, 2.007727e-23, 2.007725e-23, 2.007725e-23, 2.007723e-23, 
    2.007724e-23, 2.007723e-23, 2.007724e-23, 2.007723e-23, 2.007724e-23, 
    2.007724e-23, 2.007725e-23, 2.007727e-23, 2.007726e-23, 2.007728e-23, 
    2.007729e-23, 2.00773e-23, 2.007731e-23, 2.007731e-23, 2.007731e-23, 
    2.00773e-23, 2.007729e-23, 2.007728e-23, 2.007728e-23, 2.007728e-23, 
    2.007727e-23, 2.007726e-23, 2.007725e-23, 2.007725e-23, 2.007724e-23, 
    2.007724e-23, 2.007723e-23, 2.007723e-23, 2.007723e-23, 2.007724e-23, 
    2.007724e-23, 2.007725e-23, 2.007725e-23, 2.007728e-23, 2.007729e-23, 
    2.007729e-23, 2.00773e-23, 2.007731e-23, 2.00773e-23, 2.00773e-23, 
    2.00773e-23, 2.007729e-23, 2.007729e-23, 2.007728e-23, 2.007728e-23, 
    2.007726e-23, 2.007727e-23, 2.007724e-23, 2.007725e-23, 2.007724e-23, 
    2.007724e-23, 2.007724e-23, 2.007724e-23, 2.007723e-23, 2.007723e-23, 
    2.007723e-23, 2.007722e-23, 2.007724e-23, 2.007723e-23, 2.007729e-23, 
    2.007729e-23, 2.007729e-23, 2.00773e-23, 2.00773e-23, 2.007731e-23, 
    2.00773e-23, 2.00773e-23, 2.007729e-23, 2.007729e-23, 2.007728e-23, 
    2.007728e-23, 2.007727e-23, 2.007725e-23, 2.007725e-23, 2.007724e-23, 
    2.007725e-23, 2.007724e-23, 2.007725e-23, 2.007725e-23, 2.007723e-23, 
    2.007724e-23, 2.007722e-23, 2.007722e-23, 2.007723e-23, 2.007722e-23, 
    2.007729e-23, 2.007729e-23, 2.00773e-23, 2.00773e-23, 2.007731e-23, 
    2.00773e-23, 2.00773e-23, 2.007728e-23, 2.007728e-23, 2.007728e-23, 
    2.007728e-23, 2.007727e-23, 2.007726e-23, 2.007725e-23, 2.007724e-23, 
    2.007724e-23, 2.007724e-23, 2.007724e-23, 2.007724e-23, 2.007724e-23, 
    2.007724e-23, 2.007724e-23, 2.007722e-23, 2.007723e-23, 2.007722e-23, 
    2.007723e-23, 2.007729e-23, 2.007729e-23, 2.007729e-23, 2.007729e-23, 
    2.007729e-23, 2.007728e-23, 2.007728e-23, 2.007726e-23, 2.007727e-23, 
    2.007726e-23, 2.007727e-23, 2.007727e-23, 2.007726e-23, 2.007727e-23, 
    2.007725e-23, 2.007726e-23, 2.007724e-23, 2.007725e-23, 2.007724e-23, 
    2.007724e-23, 2.007724e-23, 2.007723e-23, 2.007723e-23, 2.007722e-23, 
    2.007722e-23, 2.007721e-23, 2.007729e-23, 2.007728e-23, 2.007728e-23, 
    2.007728e-23, 2.007727e-23, 2.007727e-23, 2.007725e-23, 2.007726e-23, 
    2.007725e-23, 2.007725e-23, 2.007726e-23, 2.007725e-23, 2.007728e-23, 
    2.007728e-23, 2.007728e-23, 2.007728e-23, 2.007726e-23, 2.007727e-23, 
    2.007725e-23, 2.007725e-23, 2.007723e-23, 2.007724e-23, 2.007722e-23, 
    2.007721e-23, 2.00772e-23, 2.007719e-23, 2.007728e-23, 2.007728e-23, 
    2.007728e-23, 2.007727e-23, 2.007726e-23, 2.007725e-23, 2.007725e-23, 
    2.007725e-23, 2.007725e-23, 2.007724e-23, 2.007725e-23, 2.007724e-23, 
    2.007727e-23, 2.007726e-23, 2.007728e-23, 2.007728e-23, 2.007727e-23, 
    2.007727e-23, 2.007726e-23, 2.007726e-23, 2.007725e-23, 2.007725e-23, 
    2.007722e-23, 2.007723e-23, 2.007719e-23, 2.00772e-23, 2.007728e-23, 
    2.007728e-23, 2.007727e-23, 2.007727e-23, 2.007725e-23, 2.007725e-23, 
    2.007725e-23, 2.007724e-23, 2.007724e-23, 2.007724e-23, 2.007724e-23, 
    2.007724e-23, 2.007725e-23, 2.007725e-23, 2.007727e-23, 2.007726e-23, 
    2.007726e-23, 2.007727e-23, 2.007726e-23, 2.007725e-23, 2.007725e-23, 
    2.007725e-23, 2.007724e-23, 2.007725e-23, 2.007721e-23, 2.007724e-23, 
    2.007728e-23, 2.007727e-23, 2.007727e-23, 2.007727e-23, 2.007725e-23, 
    2.007726e-23, 2.007724e-23, 2.007724e-23, 2.007723e-23, 2.007724e-23, 
    2.007724e-23, 2.007724e-23, 2.007725e-23, 2.007726e-23, 2.007726e-23, 
    2.007727e-23, 2.007727e-23, 2.007726e-23, 2.007725e-23, 2.007724e-23, 
    2.007724e-23, 2.007723e-23, 2.007725e-23, 2.007725e-23, 2.007725e-23, 
    2.007724e-23, 2.007726e-23, 2.007724e-23, 2.007726e-23, 2.007726e-23, 
    2.007726e-23, 2.007725e-23, 2.007724e-23, 2.007724e-23, 2.007724e-23, 
    2.007725e-23, 2.007725e-23, 2.007726e-23, 2.007726e-23, 2.007726e-23, 
    2.007727e-23, 2.007726e-23, 2.007726e-23, 2.007725e-23, 2.007724e-23, 
    2.007723e-23, 2.007723e-23, 2.007722e-23, 2.007723e-23, 2.007721e-23, 
    2.007722e-23, 2.00772e-23, 2.007724e-23, 2.007723e-23, 2.007726e-23, 
    2.007725e-23, 2.007725e-23, 2.007723e-23, 2.007724e-23, 2.007723e-23, 
    2.007725e-23, 2.007726e-23, 2.007726e-23, 2.007727e-23, 2.007726e-23, 
    2.007726e-23, 2.007726e-23, 2.007726e-23, 2.007725e-23, 2.007725e-23, 
    2.007724e-23, 2.007723e-23, 2.007721e-23, 2.00772e-23, 2.007719e-23, 
    2.007719e-23, 2.007719e-23, 2.007719e-23 ;

 COL_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_NTRUNC =
  2.052861e-24, 2.05286e-24, 2.05286e-24, 2.052859e-24, 2.05286e-24, 
    2.052859e-24, 2.052861e-24, 2.05286e-24, 2.052861e-24, 2.052861e-24, 
    2.052857e-24, 2.052859e-24, 2.052855e-24, 2.052856e-24, 2.052853e-24, 
    2.052855e-24, 2.052852e-24, 2.052853e-24, 2.052851e-24, 2.052852e-24, 
    2.05285e-24, 2.052851e-24, 2.052848e-24, 2.05285e-24, 2.05285e-24, 
    2.052851e-24, 2.052859e-24, 2.052857e-24, 2.052859e-24, 2.052858e-24, 
    2.052858e-24, 2.05286e-24, 2.05286e-24, 2.052861e-24, 2.052861e-24, 
    2.05286e-24, 2.052858e-24, 2.052859e-24, 2.052857e-24, 2.052857e-24, 
    2.052855e-24, 2.052856e-24, 2.052853e-24, 2.052854e-24, 2.052852e-24, 
    2.052852e-24, 2.052852e-24, 2.052852e-24, 2.052852e-24, 2.052853e-24, 
    2.052852e-24, 2.052853e-24, 2.052856e-24, 2.052855e-24, 2.052858e-24, 
    2.05286e-24, 2.052861e-24, 2.052862e-24, 2.052862e-24, 2.052861e-24, 
    2.05286e-24, 2.052859e-24, 2.052858e-24, 2.052858e-24, 2.052857e-24, 
    2.052856e-24, 2.052855e-24, 2.052853e-24, 2.052853e-24, 2.052853e-24, 
    2.052852e-24, 2.052851e-24, 2.052851e-24, 2.052851e-24, 2.052853e-24, 
    2.052852e-24, 2.052854e-24, 2.052853e-24, 2.052857e-24, 2.052859e-24, 
    2.052859e-24, 2.05286e-24, 2.052862e-24, 2.052861e-24, 2.052861e-24, 
    2.05286e-24, 2.052859e-24, 2.05286e-24, 2.052858e-24, 2.052859e-24, 
    2.052855e-24, 2.052856e-24, 2.052852e-24, 2.052853e-24, 2.052852e-24, 
    2.052853e-24, 2.052852e-24, 2.052853e-24, 2.052851e-24, 2.052851e-24, 
    2.052851e-24, 2.05285e-24, 2.052853e-24, 2.052852e-24, 2.05286e-24, 
    2.05286e-24, 2.052859e-24, 2.05286e-24, 2.05286e-24, 2.052861e-24, 
    2.052861e-24, 2.05286e-24, 2.052859e-24, 2.052859e-24, 2.052858e-24, 
    2.052857e-24, 2.052856e-24, 2.052855e-24, 2.052853e-24, 2.052852e-24, 
    2.052853e-24, 2.052853e-24, 2.052853e-24, 2.052853e-24, 2.052851e-24, 
    2.052852e-24, 2.05285e-24, 2.05285e-24, 2.052851e-24, 2.05285e-24, 
    2.05286e-24, 2.05286e-24, 2.052861e-24, 2.05286e-24, 2.052861e-24, 
    2.052861e-24, 2.05286e-24, 2.052859e-24, 2.052858e-24, 2.052858e-24, 
    2.052857e-24, 2.052856e-24, 2.052855e-24, 2.052853e-24, 2.052852e-24, 
    2.052852e-24, 2.052852e-24, 2.052852e-24, 2.052853e-24, 2.052852e-24, 
    2.052852e-24, 2.052852e-24, 2.05285e-24, 2.052851e-24, 2.05285e-24, 
    2.05285e-24, 2.05286e-24, 2.052859e-24, 2.05286e-24, 2.052859e-24, 
    2.052859e-24, 2.052858e-24, 2.052857e-24, 2.052855e-24, 2.052856e-24, 
    2.052855e-24, 2.052856e-24, 2.052856e-24, 2.052855e-24, 2.052856e-24, 
    2.052854e-24, 2.052855e-24, 2.052852e-24, 2.052854e-24, 2.052852e-24, 
    2.052852e-24, 2.052852e-24, 2.052851e-24, 2.05285e-24, 2.052849e-24, 
    2.05285e-24, 2.052849e-24, 2.052859e-24, 2.052858e-24, 2.052858e-24, 
    2.052857e-24, 2.052857e-24, 2.052856e-24, 2.052854e-24, 2.052855e-24, 
    2.052854e-24, 2.052854e-24, 2.052855e-24, 2.052854e-24, 2.052858e-24, 
    2.052857e-24, 2.052857e-24, 2.052859e-24, 2.052855e-24, 2.052857e-24, 
    2.052853e-24, 2.052854e-24, 2.052851e-24, 2.052853e-24, 2.05285e-24, 
    2.052848e-24, 2.052847e-24, 2.052846e-24, 2.052858e-24, 2.052858e-24, 
    2.052857e-24, 2.052856e-24, 2.052855e-24, 2.052854e-24, 2.052854e-24, 
    2.052854e-24, 2.052853e-24, 2.052853e-24, 2.052854e-24, 2.052853e-24, 
    2.052857e-24, 2.052855e-24, 2.052858e-24, 2.052857e-24, 2.052856e-24, 
    2.052857e-24, 2.052855e-24, 2.052855e-24, 2.052853e-24, 2.052854e-24, 
    2.052849e-24, 2.052851e-24, 2.052845e-24, 2.052846e-24, 2.052858e-24, 
    2.052858e-24, 2.052856e-24, 2.052857e-24, 2.052854e-24, 2.052854e-24, 
    2.052853e-24, 2.052852e-24, 2.052852e-24, 2.052852e-24, 2.052852e-24, 
    2.052852e-24, 2.052854e-24, 2.052853e-24, 2.052856e-24, 2.052855e-24, 
    2.052856e-24, 2.052856e-24, 2.052855e-24, 2.052854e-24, 2.052854e-24, 
    2.052853e-24, 2.052852e-24, 2.052854e-24, 2.052848e-24, 2.052852e-24, 
    2.052857e-24, 2.052856e-24, 2.052856e-24, 2.052856e-24, 2.052854e-24, 
    2.052855e-24, 2.052852e-24, 2.052853e-24, 2.052851e-24, 2.052852e-24, 
    2.052852e-24, 2.052853e-24, 2.052853e-24, 2.052855e-24, 2.052855e-24, 
    2.052856e-24, 2.052856e-24, 2.052855e-24, 2.052854e-24, 2.052852e-24, 
    2.052853e-24, 2.052851e-24, 2.052854e-24, 2.052853e-24, 2.052854e-24, 
    2.052852e-24, 2.052855e-24, 2.052853e-24, 2.052855e-24, 2.052855e-24, 
    2.052855e-24, 2.052853e-24, 2.052853e-24, 2.052852e-24, 2.052853e-24, 
    2.052854e-24, 2.052854e-24, 2.052855e-24, 2.052855e-24, 2.052855e-24, 
    2.052856e-24, 2.052855e-24, 2.052855e-24, 2.052854e-24, 2.052852e-24, 
    2.052851e-24, 2.052851e-24, 2.052849e-24, 2.052851e-24, 2.052848e-24, 
    2.05285e-24, 2.052847e-24, 2.052853e-24, 2.05285e-24, 2.052855e-24, 
    2.052854e-24, 2.052853e-24, 2.052851e-24, 2.052852e-24, 2.052851e-24, 
    2.052854e-24, 2.052855e-24, 2.052855e-24, 2.052856e-24, 2.052855e-24, 
    2.052855e-24, 2.052855e-24, 2.052855e-24, 2.052854e-24, 2.052855e-24, 
    2.052852e-24, 2.052851e-24, 2.052849e-24, 2.052847e-24, 2.052846e-24, 
    2.052845e-24, 2.052845e-24, 2.052845e-24 ;

 CONC_CH4_SAT =
  7.839918e-08, 7.851e-08, 7.848841e-08, 7.857779e-08, 7.852815e-08, 
    7.858671e-08, 7.842156e-08, 7.851449e-08, 7.845512e-08, 7.840902e-08, 
    7.875109e-08, 7.858175e-08, 7.892534e-08, 7.881798e-08, 7.908691e-08, 
    7.890878e-08, 7.91227e-08, 7.908154e-08, 7.920473e-08, 7.916946e-08, 
    7.932718e-08, 7.9221e-08, 7.940834e-08, 7.930171e-08, 7.93185e-08, 
    7.921754e-08, 7.861564e-08, 7.873011e-08, 7.860891e-08, 7.862523e-08, 
    7.861786e-08, 7.852925e-08, 7.84847e-08, 7.839053e-08, 7.84076e-08, 
    7.847666e-08, 7.863257e-08, 7.857955e-08, 7.871261e-08, 7.87096e-08, 
    7.885748e-08, 7.879087e-08, 7.903854e-08, 7.896822e-08, 7.917092e-08, 
    7.912006e-08, 7.916858e-08, 7.915384e-08, 7.916877e-08, 7.909414e-08, 
    7.912615e-08, 7.906034e-08, 7.88034e-08, 7.887913e-08, 7.865301e-08, 
    7.851689e-08, 7.842568e-08, 7.836104e-08, 7.837019e-08, 7.838766e-08, 
    7.847707e-08, 7.85608e-08, 7.862457e-08, 7.866722e-08, 7.870917e-08, 
    7.883656e-08, 7.890332e-08, 7.905286e-08, 7.90257e-08, 7.907154e-08, 
    7.911499e-08, 7.918813e-08, 7.917608e-08, 7.920832e-08, 7.907018e-08, 
    7.916211e-08, 7.901028e-08, 7.905188e-08, 7.872138e-08, 7.859382e-08, 
    7.85402e-08, 7.84926e-08, 7.837723e-08, 7.845697e-08, 7.842556e-08, 
    7.850007e-08, 7.854747e-08, 7.8524e-08, 7.866839e-08, 7.861233e-08, 
    7.890728e-08, 7.878045e-08, 7.910992e-08, 7.903126e-08, 7.912873e-08, 
    7.907898e-08, 7.916426e-08, 7.908751e-08, 7.922025e-08, 7.92492e-08, 
    7.922943e-08, 7.930502e-08, 7.908328e-08, 7.916866e-08, 7.852338e-08, 
    7.852721e-08, 7.854498e-08, 7.846687e-08, 7.846204e-08, 7.83901e-08, 
    7.845404e-08, 7.848131e-08, 7.855015e-08, 7.859098e-08, 7.86297e-08, 
    7.871472e-08, 7.880963e-08, 7.894178e-08, 7.903638e-08, 7.909971e-08, 
    7.906083e-08, 7.909517e-08, 7.905681e-08, 7.903879e-08, 7.92384e-08, 
    7.912649e-08, 7.929416e-08, 7.928487e-08, 7.920912e-08, 7.928592e-08, 
    7.852989e-08, 7.850785e-08, 7.843153e-08, 7.849127e-08, 7.838226e-08, 
    7.844341e-08, 7.847859e-08, 7.861368e-08, 7.864312e-08, 7.867065e-08, 
    7.872479e-08, 7.879428e-08, 7.891598e-08, 7.902149e-08, 7.911748e-08, 
    7.911044e-08, 7.911293e-08, 7.913443e-08, 7.908126e-08, 7.914315e-08, 
    7.915361e-08, 7.912638e-08, 7.928363e-08, 7.923875e-08, 7.928467e-08, 
    7.925544e-08, 7.8515e-08, 7.855203e-08, 7.853204e-08, 7.856968e-08, 
    7.854322e-08, 7.866095e-08, 7.86962e-08, 7.886053e-08, 7.879296e-08, 
    7.890024e-08, 7.880381e-08, 7.882095e-08, 7.890407e-08, 7.880897e-08, 
    7.901583e-08, 7.887598e-08, 7.913527e-08, 7.899629e-08, 7.914398e-08, 
    7.911707e-08, 7.916154e-08, 7.920141e-08, 7.925138e-08, 7.934367e-08, 
    7.932228e-08, 7.939923e-08, 7.860712e-08, 7.865513e-08, 7.865075e-08, 
    7.870084e-08, 7.873789e-08, 7.88179e-08, 7.894611e-08, 7.889788e-08, 
    7.89862e-08, 7.900397e-08, 7.886968e-08, 7.895233e-08, 7.868712e-08, 
    7.873023e-08, 7.870445e-08, 7.8611e-08, 7.890921e-08, 7.875649e-08, 
    7.903796e-08, 7.895549e-08, 7.919575e-08, 7.907657e-08, 7.931054e-08, 
    7.941059e-08, 7.950385e-08, 7.961341e-08, 7.868115e-08, 7.864856e-08, 
    7.870675e-08, 7.878743e-08, 7.886172e-08, 7.896055e-08, 7.897057e-08, 
    7.89891e-08, 7.903688e-08, 7.90771e-08, 7.899511e-08, 7.908716e-08, 
    7.874053e-08, 7.892238e-08, 7.863638e-08, 7.872288e-08, 7.878261e-08, 
    7.875627e-08, 7.889233e-08, 7.89244e-08, 7.905454e-08, 7.898722e-08, 
    7.938606e-08, 7.921005e-08, 7.969614e-08, 7.956093e-08, 7.863721e-08, 
    7.868096e-08, 7.883315e-08, 7.876078e-08, 7.896706e-08, 7.901777e-08, 
    7.905881e-08, 7.911148e-08, 7.911705e-08, 7.914821e-08, 7.909716e-08, 
    7.914613e-08, 7.896076e-08, 7.904367e-08, 7.88156e-08, 7.88713e-08, 
    7.884562e-08, 7.881757e-08, 7.890413e-08, 7.899644e-08, 7.899816e-08, 
    7.902776e-08, 7.911151e-08, 7.896789e-08, 7.940917e-08, 7.913756e-08, 
    7.872864e-08, 7.881306e-08, 7.88248e-08, 7.879218e-08, 7.901269e-08, 
    7.893294e-08, 7.914741e-08, 7.90895e-08, 7.91843e-08, 7.913723e-08, 
    7.913032e-08, 7.906974e-08, 7.903205e-08, 7.893665e-08, 7.885882e-08, 
    7.879689e-08, 7.881128e-08, 7.887927e-08, 7.900202e-08, 7.911767e-08, 
    7.909239e-08, 7.917709e-08, 7.895214e-08, 7.904673e-08, 7.901027e-08, 
    7.910522e-08, 7.889665e-08, 7.907506e-08, 7.885104e-08, 7.887067e-08, 
    7.893136e-08, 7.90533e-08, 7.907987e-08, 7.910867e-08, 7.909085e-08, 
    7.900508e-08, 7.899091e-08, 7.892982e-08, 7.891307e-08, 7.886638e-08, 
    7.88278e-08, 7.886311e-08, 7.890021e-08, 7.900502e-08, 7.909941e-08, 
    7.920202e-08, 7.9227e-08, 7.934715e-08, 7.92497e-08, 7.941073e-08, 
    7.927436e-08, 7.95099e-08, 7.908502e-08, 7.926986e-08, 7.893404e-08, 
    7.897027e-08, 7.9036e-08, 7.918589e-08, 7.910477e-08, 7.91995e-08, 
    7.899033e-08, 7.888174e-08, 7.88533e-08, 7.88007e-08, 7.885451e-08, 
    7.885012e-08, 7.890157e-08, 7.888503e-08, 7.900849e-08, 7.89422e-08, 
    7.913021e-08, 7.919869e-08, 7.939126e-08, 7.950906e-08, 7.962825e-08, 
    7.96809e-08, 7.969689e-08, 7.970359e-08,
  2.100338e-10, 2.106256e-10, 2.105103e-10, 2.109883e-10, 2.107226e-10, 
    2.110363e-10, 2.101533e-10, 2.106495e-10, 2.103325e-10, 2.100864e-10, 
    2.119223e-10, 2.110096e-10, 2.128642e-10, 2.122838e-10, 2.137394e-10, 
    2.127746e-10, 2.139335e-10, 2.137104e-10, 2.143788e-10, 2.141873e-10, 
    2.150441e-10, 2.144672e-10, 2.154858e-10, 2.149057e-10, 2.149969e-10, 
    2.144483e-10, 2.111923e-10, 2.118091e-10, 2.11156e-10, 2.112439e-10, 
    2.112042e-10, 2.107285e-10, 2.104903e-10, 2.099878e-10, 2.100788e-10, 
    2.104475e-10, 2.112834e-10, 2.109979e-10, 2.117151e-10, 2.116989e-10, 
    2.124973e-10, 2.121374e-10, 2.134773e-10, 2.130965e-10, 2.141953e-10, 
    2.139193e-10, 2.141825e-10, 2.141026e-10, 2.141836e-10, 2.137787e-10, 
    2.139523e-10, 2.135955e-10, 2.122051e-10, 2.126144e-10, 2.113936e-10, 
    2.106622e-10, 2.101753e-10, 2.098304e-10, 2.098792e-10, 2.099724e-10, 
    2.104496e-10, 2.108971e-10, 2.112404e-10, 2.114703e-10, 2.116965e-10, 
    2.12384e-10, 2.127451e-10, 2.135548e-10, 2.134078e-10, 2.136561e-10, 
    2.138918e-10, 2.142887e-10, 2.142232e-10, 2.143983e-10, 2.136488e-10, 
    2.141474e-10, 2.133242e-10, 2.135496e-10, 2.11762e-10, 2.110747e-10, 
    2.107868e-10, 2.105326e-10, 2.099168e-10, 2.103423e-10, 2.101747e-10, 
    2.105726e-10, 2.108259e-10, 2.107005e-10, 2.114766e-10, 2.111745e-10, 
    2.127665e-10, 2.120811e-10, 2.138643e-10, 2.134379e-10, 2.139663e-10, 
    2.136965e-10, 2.141591e-10, 2.137428e-10, 2.144631e-10, 2.146203e-10, 
    2.145129e-10, 2.149238e-10, 2.137198e-10, 2.141829e-10, 2.106971e-10, 
    2.107176e-10, 2.108126e-10, 2.103951e-10, 2.103694e-10, 2.099855e-10, 
    2.103267e-10, 2.104723e-10, 2.108403e-10, 2.110594e-10, 2.11268e-10, 
    2.117264e-10, 2.122387e-10, 2.129533e-10, 2.134656e-10, 2.138089e-10, 
    2.135982e-10, 2.137843e-10, 2.135764e-10, 2.134787e-10, 2.145616e-10, 
    2.139541e-10, 2.148647e-10, 2.148142e-10, 2.144026e-10, 2.148199e-10, 
    2.107319e-10, 2.106142e-10, 2.102065e-10, 2.105256e-10, 2.099436e-10, 
    2.102699e-10, 2.104577e-10, 2.111816e-10, 2.113404e-10, 2.114887e-10, 
    2.117808e-10, 2.121559e-10, 2.128137e-10, 2.133849e-10, 2.139054e-10, 
    2.138672e-10, 2.138806e-10, 2.139973e-10, 2.137089e-10, 2.140446e-10, 
    2.141012e-10, 2.139536e-10, 2.148075e-10, 2.145636e-10, 2.148132e-10, 
    2.146543e-10, 2.106524e-10, 2.108503e-10, 2.107434e-10, 2.109447e-10, 
    2.108032e-10, 2.114364e-10, 2.116264e-10, 2.125137e-10, 2.121487e-10, 
    2.127285e-10, 2.122073e-10, 2.122999e-10, 2.12749e-10, 2.122352e-10, 
    2.133542e-10, 2.125972e-10, 2.140018e-10, 2.132482e-10, 2.140491e-10, 
    2.139031e-10, 2.141444e-10, 2.143608e-10, 2.146322e-10, 2.151339e-10, 
    2.150176e-10, 2.154363e-10, 2.111464e-10, 2.11405e-10, 2.113815e-10, 
    2.116516e-10, 2.118514e-10, 2.122835e-10, 2.129767e-10, 2.127159e-10, 
    2.131939e-10, 2.1329e-10, 2.125634e-10, 2.130103e-10, 2.115775e-10, 
    2.1181e-10, 2.11671e-10, 2.111672e-10, 2.12777e-10, 2.119517e-10, 
    2.134742e-10, 2.130275e-10, 2.1433e-10, 2.136833e-10, 2.149537e-10, 
    2.15498e-10, 2.160063e-10, 2.166037e-10, 2.115454e-10, 2.113697e-10, 
    2.116835e-10, 2.121188e-10, 2.125203e-10, 2.130549e-10, 2.131092e-10, 
    2.132095e-10, 2.134684e-10, 2.136863e-10, 2.132419e-10, 2.137409e-10, 
    2.118653e-10, 2.128483e-10, 2.11304e-10, 2.117703e-10, 2.120928e-10, 
    2.119506e-10, 2.126859e-10, 2.128593e-10, 2.135639e-10, 2.131993e-10, 
    2.153644e-10, 2.144075e-10, 2.170557e-10, 2.163174e-10, 2.113085e-10, 
    2.115444e-10, 2.123658e-10, 2.11975e-10, 2.130902e-10, 2.133648e-10, 
    2.135872e-10, 2.138727e-10, 2.13903e-10, 2.14072e-10, 2.137951e-10, 
    2.140608e-10, 2.13056e-10, 2.135051e-10, 2.122711e-10, 2.125721e-10, 
    2.124333e-10, 2.122817e-10, 2.127497e-10, 2.132491e-10, 2.132586e-10, 
    2.134189e-10, 2.138724e-10, 2.130947e-10, 2.154899e-10, 2.140138e-10, 
    2.118016e-10, 2.122572e-10, 2.123208e-10, 2.121446e-10, 2.133373e-10, 
    2.129055e-10, 2.140677e-10, 2.137536e-10, 2.142679e-10, 2.140124e-10, 
    2.139749e-10, 2.136464e-10, 2.134422e-10, 2.129255e-10, 2.125046e-10, 
    2.1217e-10, 2.122477e-10, 2.126152e-10, 2.132794e-10, 2.139063e-10, 
    2.137692e-10, 2.142288e-10, 2.130094e-10, 2.135216e-10, 2.133241e-10, 
    2.138388e-10, 2.127092e-10, 2.136748e-10, 2.124626e-10, 2.125687e-10, 
    2.128969e-10, 2.135572e-10, 2.137014e-10, 2.138574e-10, 2.137609e-10, 
    2.13296e-10, 2.132193e-10, 2.128887e-10, 2.127979e-10, 2.125455e-10, 
    2.12337e-10, 2.125278e-10, 2.127284e-10, 2.132957e-10, 2.138072e-10, 
    2.143641e-10, 2.144998e-10, 2.151525e-10, 2.146228e-10, 2.154984e-10, 
    2.147565e-10, 2.160389e-10, 2.13729e-10, 2.147323e-10, 2.129115e-10, 
    2.131076e-10, 2.134634e-10, 2.142763e-10, 2.138364e-10, 2.143503e-10, 
    2.132162e-10, 2.126284e-10, 2.124748e-10, 2.121906e-10, 2.124813e-10, 
    2.124576e-10, 2.127358e-10, 2.126464e-10, 2.133145e-10, 2.129557e-10, 
    2.139743e-10, 2.143459e-10, 2.153928e-10, 2.160345e-10, 2.16685e-10, 
    2.169725e-10, 2.170599e-10, 2.170965e-10,
  1.163728e-13, 1.168086e-13, 1.167237e-13, 1.170758e-13, 1.168801e-13, 
    1.171111e-13, 1.164608e-13, 1.168262e-13, 1.165927e-13, 1.164116e-13, 
    1.177633e-13, 1.170915e-13, 1.184582e-13, 1.180301e-13, 1.191076e-13, 
    1.18392e-13, 1.192548e-13, 1.190857e-13, 1.195928e-13, 1.194475e-13, 
    1.200977e-13, 1.196598e-13, 1.204336e-13, 1.199927e-13, 1.20062e-13, 
    1.196455e-13, 1.17226e-13, 1.176799e-13, 1.171992e-13, 1.172639e-13, 
    1.172347e-13, 1.168844e-13, 1.167088e-13, 1.16339e-13, 1.16406e-13, 
    1.166774e-13, 1.17293e-13, 1.170829e-13, 1.17611e-13, 1.17599e-13, 
    1.181876e-13, 1.179222e-13, 1.189111e-13, 1.186298e-13, 1.194535e-13, 
    1.192441e-13, 1.194438e-13, 1.193832e-13, 1.194446e-13, 1.191375e-13, 
    1.192691e-13, 1.189987e-13, 1.179721e-13, 1.182739e-13, 1.173742e-13, 
    1.168354e-13, 1.16477e-13, 1.162232e-13, 1.162591e-13, 1.163276e-13, 
    1.16679e-13, 1.170087e-13, 1.172614e-13, 1.174307e-13, 1.175973e-13, 
    1.181038e-13, 1.183703e-13, 1.189683e-13, 1.188597e-13, 1.190445e-13, 
    1.192233e-13, 1.195243e-13, 1.194747e-13, 1.196075e-13, 1.190391e-13, 
    1.194171e-13, 1.187981e-13, 1.189645e-13, 1.176452e-13, 1.171395e-13, 
    1.169272e-13, 1.167401e-13, 1.162867e-13, 1.165999e-13, 1.164765e-13, 
    1.167696e-13, 1.169562e-13, 1.168638e-13, 1.174353e-13, 1.172129e-13, 
    1.183861e-13, 1.178807e-13, 1.192024e-13, 1.18882e-13, 1.192798e-13, 
    1.190753e-13, 1.19426e-13, 1.191103e-13, 1.196567e-13, 1.19776e-13, 
    1.196945e-13, 1.200066e-13, 1.190929e-13, 1.194441e-13, 1.168614e-13, 
    1.168764e-13, 1.169464e-13, 1.166388e-13, 1.166199e-13, 1.163373e-13, 
    1.165885e-13, 1.166957e-13, 1.169668e-13, 1.171282e-13, 1.172817e-13, 
    1.176193e-13, 1.179968e-13, 1.18524e-13, 1.189024e-13, 1.191605e-13, 
    1.190007e-13, 1.191418e-13, 1.189843e-13, 1.189122e-13, 1.197315e-13, 
    1.192705e-13, 1.199617e-13, 1.199233e-13, 1.196107e-13, 1.199277e-13, 
    1.16887e-13, 1.168003e-13, 1.165e-13, 1.16735e-13, 1.163065e-13, 
    1.165467e-13, 1.166849e-13, 1.172181e-13, 1.17335e-13, 1.174442e-13, 
    1.176594e-13, 1.179358e-13, 1.18421e-13, 1.188428e-13, 1.192336e-13, 
    1.192046e-13, 1.192148e-13, 1.193033e-13, 1.190846e-13, 1.193391e-13, 
    1.193821e-13, 1.192701e-13, 1.199182e-13, 1.19733e-13, 1.199225e-13, 
    1.198019e-13, 1.168284e-13, 1.169742e-13, 1.168955e-13, 1.170437e-13, 
    1.169395e-13, 1.174056e-13, 1.175455e-13, 1.181996e-13, 1.179305e-13, 
    1.183581e-13, 1.179737e-13, 1.18042e-13, 1.183731e-13, 1.179943e-13, 
    1.1882e-13, 1.182612e-13, 1.193067e-13, 1.187417e-13, 1.193426e-13, 
    1.192319e-13, 1.194149e-13, 1.19579e-13, 1.197851e-13, 1.201661e-13, 
    1.200778e-13, 1.20396e-13, 1.171922e-13, 1.173825e-13, 1.173653e-13, 
    1.175642e-13, 1.177114e-13, 1.180299e-13, 1.185414e-13, 1.183489e-13, 
    1.187017e-13, 1.187728e-13, 1.182364e-13, 1.185662e-13, 1.175096e-13, 
    1.176808e-13, 1.175785e-13, 1.172075e-13, 1.183939e-13, 1.177852e-13, 
    1.189088e-13, 1.185789e-13, 1.195557e-13, 1.190652e-13, 1.200293e-13, 
    1.204428e-13, 1.208297e-13, 1.212845e-13, 1.174859e-13, 1.173566e-13, 
    1.175877e-13, 1.179084e-13, 1.182045e-13, 1.185991e-13, 1.186392e-13, 
    1.187133e-13, 1.189045e-13, 1.190675e-13, 1.187371e-13, 1.191089e-13, 
    1.177214e-13, 1.184465e-13, 1.173082e-13, 1.176515e-13, 1.178892e-13, 
    1.177845e-13, 1.183267e-13, 1.184547e-13, 1.18975e-13, 1.187058e-13, 
    1.203411e-13, 1.196144e-13, 1.216292e-13, 1.210664e-13, 1.173116e-13, 
    1.174852e-13, 1.180905e-13, 1.178024e-13, 1.186252e-13, 1.188279e-13, 
    1.189924e-13, 1.192088e-13, 1.192318e-13, 1.193599e-13, 1.1915e-13, 
    1.193514e-13, 1.185999e-13, 1.189317e-13, 1.180208e-13, 1.182427e-13, 
    1.181405e-13, 1.180286e-13, 1.183738e-13, 1.187424e-13, 1.187495e-13, 
    1.188679e-13, 1.192081e-13, 1.186285e-13, 1.204364e-13, 1.193154e-13, 
    1.176747e-13, 1.180104e-13, 1.180574e-13, 1.179275e-13, 1.188076e-13, 
    1.184888e-13, 1.193567e-13, 1.191185e-13, 1.195086e-13, 1.193148e-13, 
    1.192863e-13, 1.190373e-13, 1.188851e-13, 1.185036e-13, 1.181929e-13, 
    1.179463e-13, 1.180036e-13, 1.182745e-13, 1.187648e-13, 1.192342e-13, 
    1.191302e-13, 1.194789e-13, 1.185655e-13, 1.189438e-13, 1.187978e-13, 
    1.191831e-13, 1.183439e-13, 1.190584e-13, 1.18162e-13, 1.182403e-13, 
    1.184825e-13, 1.1897e-13, 1.190789e-13, 1.191972e-13, 1.191241e-13, 
    1.187771e-13, 1.187205e-13, 1.184764e-13, 1.184094e-13, 1.182232e-13, 
    1.180694e-13, 1.182101e-13, 1.18358e-13, 1.187769e-13, 1.191591e-13, 
    1.195815e-13, 1.196846e-13, 1.201801e-13, 1.197778e-13, 1.204428e-13, 
    1.19879e-13, 1.208541e-13, 1.190996e-13, 1.198609e-13, 1.184932e-13, 
    1.18638e-13, 1.189008e-13, 1.195148e-13, 1.191812e-13, 1.19571e-13, 
    1.187182e-13, 1.182843e-13, 1.18171e-13, 1.179614e-13, 1.181758e-13, 
    1.181584e-13, 1.183636e-13, 1.182976e-13, 1.187908e-13, 1.185259e-13, 
    1.192858e-13, 1.195677e-13, 1.203629e-13, 1.20851e-13, 1.213466e-13, 
    1.215658e-13, 1.216324e-13, 1.216603e-13,
  1.68729e-17, 1.69449e-17, 1.693087e-17, 1.698905e-17, 1.695673e-17, 
    1.699488e-17, 1.688745e-17, 1.69478e-17, 1.690924e-17, 1.687932e-17, 
    1.710239e-17, 1.699164e-17, 1.721719e-17, 1.714649e-17, 1.732473e-17, 
    1.720624e-17, 1.734995e-17, 1.732101e-17, 1.74079e-17, 1.738299e-17, 
    1.749447e-17, 1.741939e-17, 1.755216e-17, 1.747647e-17, 1.748835e-17, 
    1.741694e-17, 1.701382e-17, 1.708862e-17, 1.700941e-17, 1.702006e-17, 
    1.701526e-17, 1.695743e-17, 1.69284e-17, 1.686734e-17, 1.68784e-17, 
    1.692321e-17, 1.702486e-17, 1.699024e-17, 1.707732e-17, 1.707535e-17, 
    1.717249e-17, 1.712868e-17, 1.729208e-17, 1.724558e-17, 1.738402e-17, 
    1.734814e-17, 1.738236e-17, 1.737197e-17, 1.738249e-17, 1.732987e-17, 
    1.735242e-17, 1.730658e-17, 1.71369e-17, 1.718675e-17, 1.703824e-17, 
    1.694931e-17, 1.689011e-17, 1.684821e-17, 1.685414e-17, 1.686545e-17, 
    1.692348e-17, 1.6978e-17, 1.701967e-17, 1.704757e-17, 1.707507e-17, 
    1.715862e-17, 1.720266e-17, 1.730154e-17, 1.728359e-17, 1.731416e-17, 
    1.734457e-17, 1.739616e-17, 1.738765e-17, 1.741041e-17, 1.731327e-17, 
    1.737776e-17, 1.72734e-17, 1.730093e-17, 1.708289e-17, 1.699956e-17, 
    1.696449e-17, 1.693358e-17, 1.68587e-17, 1.691042e-17, 1.689003e-17, 
    1.693847e-17, 1.696932e-17, 1.695405e-17, 1.704834e-17, 1.701166e-17, 
    1.720527e-17, 1.712181e-17, 1.7341e-17, 1.728727e-17, 1.735426e-17, 
    1.731927e-17, 1.737929e-17, 1.732523e-17, 1.741885e-17, 1.743929e-17, 
    1.742533e-17, 1.747886e-17, 1.732224e-17, 1.738239e-17, 1.695364e-17, 
    1.695613e-17, 1.69677e-17, 1.691685e-17, 1.691372e-17, 1.686705e-17, 
    1.690854e-17, 1.692625e-17, 1.697108e-17, 1.69977e-17, 1.702301e-17, 
    1.707869e-17, 1.714097e-17, 1.722807e-17, 1.729065e-17, 1.733382e-17, 
    1.730692e-17, 1.733062e-17, 1.73042e-17, 1.729227e-17, 1.743166e-17, 
    1.735265e-17, 1.747116e-17, 1.746458e-17, 1.741096e-17, 1.746532e-17, 
    1.695787e-17, 1.694354e-17, 1.689391e-17, 1.693275e-17, 1.686196e-17, 
    1.690162e-17, 1.692446e-17, 1.70125e-17, 1.70318e-17, 1.70498e-17, 
    1.70853e-17, 1.713092e-17, 1.721105e-17, 1.728078e-17, 1.734634e-17, 
    1.734138e-17, 1.734313e-17, 1.735827e-17, 1.732082e-17, 1.736442e-17, 
    1.737177e-17, 1.73526e-17, 1.746371e-17, 1.743194e-17, 1.746444e-17, 
    1.744375e-17, 1.694819e-17, 1.69723e-17, 1.695927e-17, 1.698378e-17, 
    1.696654e-17, 1.704342e-17, 1.706649e-17, 1.717446e-17, 1.713004e-17, 
    1.720065e-17, 1.713718e-17, 1.714845e-17, 1.720311e-17, 1.714059e-17, 
    1.7277e-17, 1.718462e-17, 1.735886e-17, 1.726403e-17, 1.7365e-17, 
    1.734605e-17, 1.73774e-17, 1.740553e-17, 1.744087e-17, 1.750623e-17, 
    1.749107e-17, 1.754571e-17, 1.700825e-17, 1.703962e-17, 1.70368e-17, 
    1.70696e-17, 1.709388e-17, 1.714646e-17, 1.723095e-17, 1.719914e-17, 
    1.725747e-17, 1.726921e-17, 1.718056e-17, 1.723504e-17, 1.706058e-17, 
    1.70888e-17, 1.707195e-17, 1.701076e-17, 1.720656e-17, 1.710605e-17, 
    1.72917e-17, 1.723715e-17, 1.740153e-17, 1.731758e-17, 1.748275e-17, 
    1.75537e-17, 1.762023e-17, 1.769841e-17, 1.705668e-17, 1.703536e-17, 
    1.707348e-17, 1.712637e-17, 1.717529e-17, 1.724049e-17, 1.724713e-17, 
    1.725937e-17, 1.729101e-17, 1.731799e-17, 1.72633e-17, 1.732498e-17, 
    1.709548e-17, 1.721526e-17, 1.702737e-17, 1.708398e-17, 1.712322e-17, 
    1.710594e-17, 1.719549e-17, 1.721664e-17, 1.730266e-17, 1.725814e-17, 
    1.753625e-17, 1.741157e-17, 1.775777e-17, 1.76609e-17, 1.702793e-17, 
    1.705658e-17, 1.715646e-17, 1.710891e-17, 1.724481e-17, 1.727833e-17, 
    1.730555e-17, 1.734208e-17, 1.734603e-17, 1.736797e-17, 1.733202e-17, 
    1.736653e-17, 1.724063e-17, 1.729549e-17, 1.714495e-17, 1.71816e-17, 
    1.716472e-17, 1.714625e-17, 1.720327e-17, 1.726418e-17, 1.726537e-17, 
    1.728493e-17, 1.734189e-17, 1.724536e-17, 1.755256e-17, 1.736028e-17, 
    1.708783e-17, 1.714321e-17, 1.715099e-17, 1.712956e-17, 1.727498e-17, 
    1.722226e-17, 1.736742e-17, 1.732662e-17, 1.739346e-17, 1.736025e-17, 
    1.735537e-17, 1.731298e-17, 1.728779e-17, 1.72247e-17, 1.717338e-17, 
    1.713265e-17, 1.714211e-17, 1.718685e-17, 1.726788e-17, 1.734644e-17, 
    1.732862e-17, 1.738838e-17, 1.723495e-17, 1.729749e-17, 1.727335e-17, 
    1.733769e-17, 1.719832e-17, 1.731641e-17, 1.716828e-17, 1.718121e-17, 
    1.722122e-17, 1.730181e-17, 1.731987e-17, 1.73401e-17, 1.732758e-17, 
    1.726992e-17, 1.726056e-17, 1.722022e-17, 1.720914e-17, 1.717839e-17, 
    1.715299e-17, 1.717622e-17, 1.720065e-17, 1.72699e-17, 1.733357e-17, 
    1.740595e-17, 1.742363e-17, 1.750859e-17, 1.743957e-17, 1.755365e-17, 
    1.745687e-17, 1.762436e-17, 1.732335e-17, 1.745381e-17, 1.7223e-17, 
    1.724694e-17, 1.729036e-17, 1.73945e-17, 1.733737e-17, 1.740413e-17, 
    1.726019e-17, 1.718845e-17, 1.716977e-17, 1.713515e-17, 1.717056e-17, 
    1.716768e-17, 1.720158e-17, 1.719068e-17, 1.72722e-17, 1.722839e-17, 
    1.735527e-17, 1.740358e-17, 1.754002e-17, 1.762387e-17, 1.770913e-17, 
    1.774687e-17, 1.775835e-17, 1.776315e-17,
  7.06754e-22, 7.101483e-22, 7.094869e-22, 7.122311e-22, 7.107067e-22, 
    7.125057e-22, 7.074399e-22, 7.102848e-22, 7.08467e-22, 7.07057e-22, 
    7.175772e-22, 7.123532e-22, 7.230047e-22, 7.196627e-22, 7.280869e-22, 
    7.224865e-22, 7.292798e-22, 7.27912e-22, 7.32022e-22, 7.308433e-22, 
    7.361396e-22, 7.325662e-22, 7.389559e-22, 7.352682e-22, 7.358417e-22, 
    7.324498e-22, 7.133993e-22, 7.169271e-22, 7.131914e-22, 7.136937e-22, 
    7.134675e-22, 7.107395e-22, 7.093695e-22, 7.064923e-22, 7.070135e-22, 
    7.091255e-22, 7.139196e-22, 7.122876e-22, 7.163962e-22, 7.163032e-22, 
    7.20892e-22, 7.188215e-22, 7.265503e-22, 7.243491e-22, 7.308924e-22, 
    7.291952e-22, 7.308133e-22, 7.30322e-22, 7.308197e-22, 7.283311e-22, 
    7.293972e-22, 7.272362e-22, 7.192098e-22, 7.215657e-22, 7.145515e-22, 
    7.103552e-22, 7.075653e-22, 7.055914e-22, 7.058704e-22, 7.06403e-22, 
    7.091379e-22, 7.117104e-22, 7.136756e-22, 7.149922e-22, 7.162898e-22, 
    7.202347e-22, 7.223176e-22, 7.269978e-22, 7.261488e-22, 7.275909e-22, 
    7.290263e-22, 7.314662e-22, 7.310638e-22, 7.321404e-22, 7.275498e-22, 
    7.305956e-22, 7.256662e-22, 7.269695e-22, 7.166563e-22, 7.127271e-22, 
    7.110718e-22, 7.096145e-22, 7.060851e-22, 7.085224e-22, 7.075614e-22, 
    7.098457e-22, 7.113008e-22, 7.105804e-22, 7.150281e-22, 7.132978e-22, 
    7.224412e-22, 7.184964e-22, 7.288573e-22, 7.263227e-22, 7.294844e-22, 
    7.278308e-22, 7.306681e-22, 7.281119e-22, 7.325402e-22, 7.335076e-22, 
    7.328467e-22, 7.353819e-22, 7.279706e-22, 7.308147e-22, 7.105608e-22, 
    7.106784e-22, 7.112246e-22, 7.088253e-22, 7.086779e-22, 7.064786e-22, 
    7.084342e-22, 7.092688e-22, 7.113841e-22, 7.126395e-22, 7.13833e-22, 
    7.164604e-22, 7.194019e-22, 7.235201e-22, 7.264829e-22, 7.285179e-22, 
    7.272526e-22, 7.283665e-22, 7.271247e-22, 7.265598e-22, 7.33146e-22, 
    7.294079e-22, 7.350171e-22, 7.347057e-22, 7.321666e-22, 7.347408e-22, 
    7.107607e-22, 7.100847e-22, 7.077445e-22, 7.095756e-22, 7.062392e-22, 
    7.081075e-22, 7.091838e-22, 7.133369e-22, 7.142478e-22, 7.150971e-22, 
    7.167728e-22, 7.189275e-22, 7.227149e-22, 7.260152e-22, 7.2911e-22, 
    7.288755e-22, 7.289582e-22, 7.29674e-22, 7.279034e-22, 7.299648e-22, 
    7.303123e-22, 7.294058e-22, 7.346641e-22, 7.3316e-22, 7.346991e-22, 
    7.337193e-22, 7.103041e-22, 7.114412e-22, 7.108268e-22, 7.11983e-22, 
    7.111694e-22, 7.147951e-22, 7.158838e-22, 7.209843e-22, 7.188857e-22, 
    7.222231e-22, 7.192234e-22, 7.197553e-22, 7.223378e-22, 7.193845e-22, 
    7.258356e-22, 7.214643e-22, 7.297018e-22, 7.252209e-22, 7.299925e-22, 
    7.290962e-22, 7.305791e-22, 7.319098e-22, 7.335828e-22, 7.367145e-22, 
    7.359754e-22, 7.386419e-22, 7.131371e-22, 7.146165e-22, 7.144837e-22, 
    7.160315e-22, 7.171778e-22, 7.196618e-22, 7.236566e-22, 7.221525e-22, 
    7.249121e-22, 7.254675e-22, 7.212738e-22, 7.238499e-22, 7.156055e-22, 
    7.169373e-22, 7.161424e-22, 7.132552e-22, 7.225025e-22, 7.177517e-22, 
    7.265324e-22, 7.239504e-22, 7.317204e-22, 7.277506e-22, 7.355692e-22, 
    7.390306e-22, 7.422822e-22, 7.461044e-22, 7.154218e-22, 7.144162e-22, 
    7.16215e-22, 7.187117e-22, 7.210245e-22, 7.241082e-22, 7.244226e-22, 
    7.250018e-22, 7.264998e-22, 7.277706e-22, 7.251874e-22, 7.281001e-22, 
    7.172514e-22, 7.229143e-22, 7.140384e-22, 7.167095e-22, 7.185633e-22, 
    7.177473e-22, 7.2198e-22, 7.2298e-22, 7.27051e-22, 7.249439e-22, 
    7.38178e-22, 7.321947e-22, 7.490114e-22, 7.442699e-22, 7.140655e-22, 
    7.154171e-22, 7.201337e-22, 7.178875e-22, 7.243129e-22, 7.258995e-22, 
    7.271884e-22, 7.289081e-22, 7.290952e-22, 7.301328e-22, 7.284331e-22, 
    7.300647e-22, 7.241148e-22, 7.26712e-22, 7.195908e-22, 7.213228e-22, 
    7.20525e-22, 7.196521e-22, 7.223477e-22, 7.252286e-22, 7.252861e-22, 
    7.262117e-22, 7.288959e-22, 7.243388e-22, 7.389722e-22, 7.297662e-22, 
    7.168925e-22, 7.195071e-22, 7.198759e-22, 7.188633e-22, 7.257405e-22, 
    7.232459e-22, 7.30107e-22, 7.281779e-22, 7.313387e-22, 7.297677e-22, 
    7.295368e-22, 7.27536e-22, 7.263474e-22, 7.233609e-22, 7.209338e-22, 
    7.190096e-22, 7.194565e-22, 7.215708e-22, 7.25404e-22, 7.291141e-22, 
    7.282715e-22, 7.310983e-22, 7.238463e-22, 7.268064e-22, 7.25663e-22, 
    7.287007e-22, 7.221134e-22, 7.276941e-22, 7.206933e-22, 7.213044e-22, 
    7.231963e-22, 7.270101e-22, 7.27859e-22, 7.288143e-22, 7.28223e-22, 
    7.255007e-22, 7.25058e-22, 7.231493e-22, 7.226248e-22, 7.21171e-22, 
    7.199704e-22, 7.210684e-22, 7.22223e-22, 7.255002e-22, 7.285058e-22, 
    7.319294e-22, 7.327666e-22, 7.368276e-22, 7.335195e-22, 7.390254e-22, 
    7.343367e-22, 7.424813e-22, 7.280213e-22, 7.341935e-22, 7.232811e-22, 
    7.244136e-22, 7.264682e-22, 7.313866e-22, 7.286857e-22, 7.318428e-22, 
    7.250404e-22, 7.216458e-22, 7.207636e-22, 7.191272e-22, 7.208011e-22, 
    7.206646e-22, 7.22268e-22, 7.217524e-22, 7.25609e-22, 7.235361e-22, 
    7.295322e-22, 7.318167e-22, 7.383638e-22, 7.42459e-22, 7.466307e-22, 
    7.484779e-22, 7.490401e-22, 7.492754e-22,
  9.115915e-27, 9.165612e-27, 9.155926e-27, 9.196131e-27, 9.173797e-27, 
    9.200157e-27, 9.125956e-27, 9.167606e-27, 9.140992e-27, 9.120354e-27, 
    9.274538e-27, 9.197922e-27, 9.354338e-27, 9.305204e-27, 9.429055e-27, 
    9.346709e-27, 9.446325e-27, 9.426534e-27, 9.486053e-27, 9.468976e-27, 
    9.545846e-27, 9.493939e-27, 9.587188e-27, 9.533106e-27, 9.541481e-27, 
    9.492252e-27, 9.213264e-27, 9.264992e-27, 9.210216e-27, 9.217577e-27, 
    9.214264e-27, 9.174274e-27, 9.154195e-27, 9.112092e-27, 9.119718e-27, 
    9.150629e-27, 9.220887e-27, 9.196968e-27, 9.257233e-27, 9.255869e-27, 
    9.323274e-27, 9.292846e-27, 9.406552e-27, 9.374138e-27, 9.469688e-27, 
    9.44511e-27, 9.468541e-27, 9.461426e-27, 9.468634e-27, 9.432599e-27, 
    9.448031e-27, 9.416652e-27, 9.298549e-27, 9.333177e-27, 9.230159e-27, 
    9.168628e-27, 9.127789e-27, 9.098914e-27, 9.102993e-27, 9.11078e-27, 
    9.15081e-27, 9.188509e-27, 9.217318e-27, 9.236629e-27, 9.255673e-27, 
    9.31359e-27, 9.34423e-27, 9.413138e-27, 9.400639e-27, 9.421834e-27, 
    9.442665e-27, 9.477997e-27, 9.47217e-27, 9.487764e-27, 9.421241e-27, 
    9.465383e-27, 9.393534e-27, 9.412729e-27, 9.261014e-27, 9.20341e-27, 
    9.17913e-27, 9.157793e-27, 9.106132e-27, 9.141797e-27, 9.127731e-27, 
    9.161184e-27, 9.182503e-27, 9.171949e-27, 9.237157e-27, 9.211777e-27, 
    9.346049e-27, 9.288065e-27, 9.440218e-27, 9.4032e-27, 9.449297e-27, 
    9.425354e-27, 9.466435e-27, 9.42943e-27, 9.493559e-27, 9.507576e-27, 
    9.497999e-27, 9.534761e-27, 9.427385e-27, 9.468556e-27, 9.17166e-27, 
    9.173382e-27, 9.181389e-27, 9.146233e-27, 9.144077e-27, 9.111891e-27, 
    9.140511e-27, 9.152729e-27, 9.183728e-27, 9.202125e-27, 9.219625e-27, 
    9.258173e-27, 9.301366e-27, 9.361929e-27, 9.405559e-27, 9.435307e-27, 
    9.416895e-27, 9.433116e-27, 9.415019e-27, 9.406697e-27, 9.502333e-27, 
    9.448185e-27, 9.529469e-27, 9.524955e-27, 9.488142e-27, 9.525463e-27, 
    9.174589e-27, 9.164688e-27, 9.130414e-27, 9.157229e-27, 9.108388e-27, 
    9.135726e-27, 9.151481e-27, 9.212342e-27, 9.225709e-27, 9.238166e-27, 
    9.262761e-27, 9.294403e-27, 9.350082e-27, 9.398666e-27, 9.443879e-27, 
    9.440485e-27, 9.441681e-27, 9.452041e-27, 9.426412e-27, 9.456251e-27, 
    9.46128e-27, 9.448159e-27, 9.524351e-27, 9.502545e-27, 9.524859e-27, 
    9.510653e-27, 9.167901e-27, 9.184562e-27, 9.175559e-27, 9.192501e-27, 
    9.180575e-27, 9.233726e-27, 9.249698e-27, 9.324622e-27, 9.293788e-27, 
    9.342846e-27, 9.298752e-27, 9.306565e-27, 9.344516e-27, 9.301121e-27, 
    9.396014e-27, 9.331675e-27, 9.452445e-27, 9.386951e-27, 9.456654e-27, 
    9.443679e-27, 9.465151e-27, 9.484424e-27, 9.508672e-27, 9.554292e-27, 
    9.543451e-27, 9.582583e-27, 9.209421e-27, 9.231112e-27, 9.229171e-27, 
    9.25188e-27, 9.268704e-27, 9.305195e-27, 9.363941e-27, 9.341814e-27, 
    9.382427e-27, 9.390604e-27, 9.328894e-27, 9.366783e-27, 9.245623e-27, 
    9.265164e-27, 9.253504e-27, 9.211147e-27, 9.346952e-27, 9.277122e-27, 
    9.406287e-27, 9.368266e-27, 9.481679e-27, 9.424168e-27, 9.537495e-27, 
    9.588273e-27, 9.637233e-27, 9.695018e-27, 9.242931e-27, 9.22818e-27, 
    9.254574e-27, 9.291225e-27, 9.325223e-27, 9.370589e-27, 9.375221e-27, 
    9.383746e-27, 9.405813e-27, 9.424472e-27, 9.386472e-27, 9.429261e-27, 
    9.269758e-27, 9.353015e-27, 9.222634e-27, 9.261817e-27, 9.289048e-27, 
    9.277066e-27, 9.33928e-27, 9.353991e-27, 9.413925e-27, 9.382896e-27, 
    9.575753e-27, 9.488541e-27, 9.739049e-27, 9.667269e-27, 9.223037e-27, 
    9.242865e-27, 9.312123e-27, 9.279126e-27, 9.373606e-27, 9.396965e-27, 
    9.415956e-27, 9.440949e-27, 9.443663e-27, 9.458684e-27, 9.43408e-27, 
    9.4577e-27, 9.370685e-27, 9.408936e-27, 9.304154e-27, 9.32961e-27, 
    9.317884e-27, 9.305054e-27, 9.344688e-27, 9.387077e-27, 9.387934e-27, 
    9.40156e-27, 9.440734e-27, 9.373989e-27, 9.587389e-27, 9.45334e-27, 
    9.26452e-27, 9.302908e-27, 9.30834e-27, 9.293463e-27, 9.394623e-27, 
    9.357898e-27, 9.458311e-27, 9.430386e-27, 9.476153e-27, 9.453399e-27, 
    9.450056e-27, 9.42104e-27, 9.403563e-27, 9.35959e-27, 9.323889e-27, 
    9.295614e-27, 9.30218e-27, 9.333254e-27, 9.389661e-27, 9.443932e-27, 
    9.431733e-27, 9.472669e-27, 9.366737e-27, 9.410321e-27, 9.393477e-27, 
    9.437951e-27, 9.341237e-27, 9.423315e-27, 9.32036e-27, 9.329344e-27, 
    9.35717e-27, 9.413315e-27, 9.425766e-27, 9.439592e-27, 9.431039e-27, 
    9.391086e-27, 9.384572e-27, 9.356481e-27, 9.348758e-27, 9.327383e-27, 
    9.309733e-27, 9.325871e-27, 9.342847e-27, 9.391084e-27, 9.435126e-27, 
    9.484707e-27, 9.496843e-27, 9.555931e-27, 9.507735e-27, 9.588168e-27, 
    9.519554e-27, 9.640204e-27, 9.428098e-27, 9.517502e-27, 9.358421e-27, 
    9.375089e-27, 9.405334e-27, 9.476832e-27, 9.437735e-27, 9.483443e-27, 
    9.384313e-27, 9.334352e-27, 9.321392e-27, 9.29734e-27, 9.321942e-27, 
    9.319938e-27, 9.343517e-27, 9.335932e-27, 9.392687e-27, 9.362173e-27, 
    9.449985e-27, 9.483069e-27, 9.578495e-27, 9.639889e-27, 9.703003e-27, 
    9.730972e-27, 9.739491e-27, 9.743055e-27,
  3.689617e-32, 3.713573e-32, 3.708902e-32, 3.728303e-32, 3.717524e-32, 
    3.730248e-32, 3.694456e-32, 3.714533e-32, 3.701702e-32, 3.691758e-32, 
    3.766635e-32, 3.729168e-32, 3.806428e-32, 3.781924e-32, 3.843745e-32, 
    3.802617e-32, 3.852255e-32, 3.84251e-32, 3.871856e-32, 3.86343e-32, 
    3.901339e-32, 3.875749e-32, 3.9216e-32, 3.895095e-32, 3.899206e-32, 
    3.874915e-32, 3.736582e-32, 3.761885e-32, 3.735109e-32, 3.738664e-32, 
    3.737065e-32, 3.717753e-32, 3.708062e-32, 3.68778e-32, 3.691452e-32, 
    3.706346e-32, 3.740263e-32, 3.728711e-32, 3.758045e-32, 3.757367e-32, 
    3.790933e-32, 3.775769e-32, 3.832532e-32, 3.816326e-32, 3.863781e-32, 
    3.851662e-32, 3.863214e-32, 3.859706e-32, 3.86326e-32, 3.845497e-32, 
    3.853101e-32, 3.837586e-32, 3.778609e-32, 3.795871e-32, 3.744747e-32, 
    3.715021e-32, 3.695338e-32, 3.681434e-32, 3.683397e-32, 3.687145e-32, 
    3.706433e-32, 3.724626e-32, 3.738543e-32, 3.747878e-32, 3.757269e-32, 
    3.786093e-32, 3.801382e-32, 3.835825e-32, 3.829576e-32, 3.840165e-32, 
    3.850457e-32, 3.867878e-32, 3.865004e-32, 3.872698e-32, 3.839874e-32, 
    3.861654e-32, 3.826023e-32, 3.835625e-32, 3.759905e-32, 3.731822e-32, 
    3.72009e-32, 3.709801e-32, 3.684908e-32, 3.702088e-32, 3.695309e-32, 
    3.71144e-32, 3.721727e-32, 3.716634e-32, 3.748134e-32, 3.735864e-32, 
    3.80229e-32, 3.773385e-32, 3.849251e-32, 3.830856e-32, 3.853726e-32, 
    3.841925e-32, 3.862174e-32, 3.843938e-32, 3.87556e-32, 3.882479e-32, 
    3.877751e-32, 3.895917e-32, 3.842931e-32, 3.86322e-32, 3.716494e-32, 
    3.717325e-32, 3.721189e-32, 3.704226e-32, 3.703187e-32, 3.687682e-32, 
    3.701471e-32, 3.70736e-32, 3.722319e-32, 3.731201e-32, 3.739656e-32, 
    3.75851e-32, 3.78001e-32, 3.810222e-32, 3.832037e-32, 3.846833e-32, 
    3.837708e-32, 3.845753e-32, 3.836772e-32, 3.832608e-32, 3.879889e-32, 
    3.853175e-32, 3.8933e-32, 3.891069e-32, 3.872883e-32, 3.891321e-32, 
    3.717907e-32, 3.713131e-32, 3.696604e-32, 3.709533e-32, 3.685996e-32, 
    3.699163e-32, 3.706755e-32, 3.736133e-32, 3.742599e-32, 3.74862e-32, 
    3.760793e-32, 3.776544e-32, 3.804307e-32, 3.828586e-32, 3.851057e-32, 
    3.849384e-32, 3.849973e-32, 3.855078e-32, 3.842451e-32, 3.857154e-32, 
    3.859631e-32, 3.853165e-32, 3.890771e-32, 3.879997e-32, 3.891022e-32, 
    3.884003e-32, 3.714681e-32, 3.722721e-32, 3.718376e-32, 3.726553e-32, 
    3.720795e-32, 3.746469e-32, 3.75429e-32, 3.7916e-32, 3.776237e-32, 
    3.800694e-32, 3.778711e-32, 3.782602e-32, 3.801519e-32, 3.779893e-32, 
    3.827255e-32, 3.795116e-32, 3.855277e-32, 3.822719e-32, 3.857352e-32, 
    3.850958e-32, 3.861543e-32, 3.87105e-32, 3.883024e-32, 3.905481e-32, 
    3.900174e-32, 3.919346e-32, 3.734727e-32, 3.745207e-32, 3.744272e-32, 
    3.755382e-32, 3.763749e-32, 3.781922e-32, 3.81123e-32, 3.800184e-32, 
    3.82047e-32, 3.824556e-32, 3.793739e-32, 3.812647e-32, 3.752268e-32, 
    3.761982e-32, 3.756188e-32, 3.735559e-32, 3.802743e-32, 3.767934e-32, 
    3.8324e-32, 3.813391e-32, 3.869695e-32, 3.841328e-32, 3.897258e-32, 
    3.922127e-32, 3.946371e-32, 3.975052e-32, 3.750931e-32, 3.743793e-32, 
    3.756723e-32, 3.774956e-32, 3.791905e-32, 3.814551e-32, 3.816867e-32, 
    3.821127e-32, 3.832165e-32, 3.841485e-32, 3.822486e-32, 3.843855e-32, 
    3.76426e-32, 3.805771e-32, 3.74111e-32, 3.760316e-32, 3.773874e-32, 
    3.767911e-32, 3.798921e-32, 3.806263e-32, 3.83622e-32, 3.820704e-32, 
    3.915988e-32, 3.873076e-32, 3.997301e-32, 3.961269e-32, 3.741307e-32, 
    3.7509e-32, 3.785371e-32, 3.768937e-32, 3.816061e-32, 3.827737e-32, 
    3.837241e-32, 3.84961e-32, 3.850949e-32, 3.858352e-32, 3.846229e-32, 
    3.857868e-32, 3.814599e-32, 3.833726e-32, 3.781405e-32, 3.794093e-32, 
    3.788248e-32, 3.781853e-32, 3.801619e-32, 3.822787e-32, 3.823222e-32, 
    3.830033e-32, 3.849483e-32, 3.816252e-32, 3.92168e-32, 3.855699e-32, 
    3.761669e-32, 3.780775e-32, 3.783489e-32, 3.776078e-32, 3.826565e-32, 
    3.808212e-32, 3.858169e-32, 3.844409e-32, 3.86697e-32, 3.855748e-32, 
    3.8541e-32, 3.839774e-32, 3.831038e-32, 3.809056e-32, 3.791239e-32, 
    3.77715e-32, 3.780421e-32, 3.79591e-32, 3.824081e-32, 3.851079e-32, 
    3.845068e-32, 3.865252e-32, 3.812628e-32, 3.834417e-32, 3.82599e-32, 
    3.848134e-32, 3.799895e-32, 3.840888e-32, 3.789483e-32, 3.793963e-32, 
    3.807848e-32, 3.83591e-32, 3.84213e-32, 3.848941e-32, 3.844731e-32, 
    3.824794e-32, 3.821539e-32, 3.807506e-32, 3.803648e-32, 3.792986e-32, 
    3.784185e-32, 3.79223e-32, 3.800696e-32, 3.824796e-32, 3.84674e-32, 
    3.871188e-32, 3.877182e-32, 3.906273e-32, 3.88255e-32, 3.922061e-32, 
    3.888374e-32, 3.947826e-32, 3.84327e-32, 3.887372e-32, 3.808475e-32, 
    3.816802e-32, 3.831918e-32, 3.867296e-32, 3.848028e-32, 3.870561e-32, 
    3.821411e-32, 3.796455e-32, 3.789997e-32, 3.778009e-32, 3.790271e-32, 
    3.789272e-32, 3.801035e-32, 3.797251e-32, 3.825598e-32, 3.810349e-32, 
    3.854063e-32, 3.870377e-32, 3.91734e-32, 3.947681e-32, 3.979031e-32, 
    3.993183e-32, 3.997529e-32, 3.999348e-32,
  4.88359e-38, 4.92606e-38, 4.917768e-38, 4.952258e-38, 4.933086e-38, 
    4.955722e-38, 4.89216e-38, 4.927762e-38, 4.904998e-38, 4.887385e-38, 
    5.020904e-38, 4.953801e-38, 5.092952e-38, 5.048544e-38, 5.162525e-38, 
    5.086026e-38, 5.178355e-38, 5.160242e-38, 5.214921e-38, 5.199188e-38, 
    5.270044e-38, 5.2222e-38, 5.307725e-38, 5.258445e-38, 5.266093e-38, 
    5.220639e-38, 4.96702e-38, 5.012339e-38, 4.964392e-38, 4.970729e-38, 
    4.96788e-38, 4.933489e-38, 4.916268e-38, 4.880346e-38, 4.886843e-38, 
    4.913229e-38, 4.973581e-38, 4.952992e-38, 5.005453e-38, 5.00423e-38, 
    5.064852e-38, 5.037421e-38, 5.141523e-38, 5.111166e-38, 5.199844e-38, 
    5.17726e-38, 5.198784e-38, 5.192244e-38, 5.198869e-38, 5.165792e-38, 
    5.179936e-38, 5.15101e-38, 5.042551e-38, 5.073799e-38, 4.981589e-38, 
    4.928619e-38, 4.893719e-38, 4.869128e-38, 4.872597e-38, 4.87922e-38, 
    4.913384e-38, 4.945719e-38, 4.97052e-38, 4.987187e-38, 5.004055e-38, 
    5.056069e-38, 5.08379e-38, 5.147697e-38, 5.135979e-38, 5.15584e-38, 
    5.175018e-38, 5.207488e-38, 5.202125e-38, 5.21649e-38, 5.155301e-38, 
    5.19587e-38, 5.129322e-38, 5.147329e-38, 5.008769e-38, 4.958534e-38, 
    4.937634e-38, 4.919364e-38, 4.875267e-38, 4.905678e-38, 4.893667e-38, 
    4.922278e-38, 4.94056e-38, 4.931506e-38, 4.987644e-38, 4.96574e-38, 
    5.085438e-38, 5.033109e-38, 5.172773e-38, 5.13838e-38, 5.181103e-38, 
    5.15915e-38, 5.19684e-38, 5.162898e-38, 5.221843e-38, 5.234788e-38, 
    5.225939e-38, 5.259996e-38, 5.161026e-38, 5.198792e-38, 4.931256e-38, 
    4.932731e-38, 4.939605e-38, 4.909469e-38, 4.907627e-38, 4.880172e-38, 
    4.904588e-38, 4.91503e-38, 4.941616e-38, 4.957428e-38, 4.972504e-38, 
    5.006286e-38, 5.045078e-38, 5.099851e-38, 5.140593e-38, 5.168279e-38, 
    5.151243e-38, 5.166271e-38, 5.149484e-38, 5.141669e-38, 5.229938e-38, 
    5.180072e-38, 5.255082e-38, 5.250897e-38, 5.216836e-38, 5.251368e-38, 
    4.933767e-38, 4.925282e-38, 4.895962e-38, 4.918891e-38, 4.877191e-38, 
    4.900495e-38, 4.913953e-38, 4.966213e-38, 4.977757e-38, 4.98851e-38, 
    5.010402e-38, 5.038822e-38, 5.089106e-38, 5.134117e-38, 5.176136e-38, 
    5.173024e-38, 5.17412e-38, 5.18362e-38, 5.160134e-38, 5.187486e-38, 
    5.1921e-38, 5.180058e-38, 5.250337e-38, 5.230148e-38, 5.250808e-38, 
    5.23765e-38, 4.928036e-38, 4.942329e-38, 4.934601e-38, 4.949147e-38, 
    4.9389e-38, 4.984659e-38, 4.998678e-38, 5.066051e-38, 5.038264e-38, 
    5.082546e-38, 5.042738e-38, 5.049771e-38, 5.084028e-38, 5.044876e-38, 
    5.131616e-38, 5.072419e-38, 5.183989e-38, 5.123107e-38, 5.187856e-38, 
    5.175952e-38, 5.195671e-38, 5.213412e-38, 5.235814e-38, 5.277743e-38, 
    5.267897e-38, 5.30353e-38, 4.963712e-38, 4.982409e-38, 4.980747e-38, 
    5.000655e-38, 5.015726e-38, 5.048545e-38, 5.101688e-38, 5.081628e-38, 
    5.118919e-38, 5.12657e-38, 5.069941e-38, 5.10428e-38, 4.995047e-38, 
    5.012533e-38, 5.002104e-38, 4.965192e-38, 5.086262e-38, 5.023266e-38, 
    5.141274e-38, 5.105675e-38, 5.21088e-38, 5.158019e-38, 5.26249e-38, 
    5.308695e-38, 5.353543e-38, 5.407339e-38, 4.992644e-38, 4.979891e-38, 
    5.003071e-38, 5.035943e-38, 5.066614e-38, 5.107842e-38, 5.112178e-38, 
    5.120147e-38, 5.140838e-38, 5.158324e-38, 5.122683e-38, 5.162743e-38, 
    5.016624e-38, 5.091764e-38, 4.975097e-38, 5.009529e-38, 5.033993e-38, 
    5.023232e-38, 5.079338e-38, 5.092666e-38, 5.148441e-38, 5.119358e-38, 
    5.297261e-38, 5.217187e-38, 5.450065e-38, 5.381144e-38, 4.975452e-38, 
    4.992593e-38, 5.054778e-38, 5.025084e-38, 5.110668e-38, 5.132529e-38, 
    5.150366e-38, 5.173438e-38, 5.175935e-38, 5.189718e-38, 5.167156e-38, 
    5.188819e-38, 5.107932e-38, 5.143765e-38, 5.047612e-38, 5.070579e-38, 
    5.059995e-38, 5.048422e-38, 5.084234e-38, 5.123246e-38, 5.124072e-38, 
    5.136832e-38, 5.173165e-38, 5.111027e-38, 5.307838e-38, 5.184741e-38, 
    5.011982e-38, 5.046458e-38, 5.051377e-38, 5.037982e-38, 5.130333e-38, 
    5.096204e-38, 5.189378e-38, 5.163773e-38, 5.205795e-38, 5.184868e-38, 
    5.181798e-38, 5.155115e-38, 5.138721e-38, 5.097735e-38, 5.065407e-38, 
    5.03992e-38, 5.045832e-38, 5.073872e-38, 5.125671e-38, 5.176172e-38, 
    5.16499e-38, 5.202588e-38, 5.104251e-38, 5.145057e-38, 5.129249e-38, 
    5.170697e-38, 5.081102e-38, 5.157166e-38, 5.06223e-38, 5.070347e-38, 
    5.095543e-38, 5.147853e-38, 5.159534e-38, 5.172194e-38, 5.164371e-38, 
    5.12701e-38, 5.120917e-38, 5.094924e-38, 5.087911e-38, 5.068577e-38, 
    5.052641e-38, 5.067204e-38, 5.082553e-38, 5.127016e-38, 5.168101e-38, 
    5.213668e-38, 5.224879e-38, 5.279195e-38, 5.234906e-38, 5.308545e-38, 
    5.245793e-38, 5.356204e-38, 5.161636e-38, 5.243937e-38, 5.096686e-38, 
    5.112056e-38, 5.140362e-38, 5.206388e-38, 5.170499e-38, 5.212488e-38, 
    5.120677e-38, 5.074853e-38, 5.063161e-38, 5.041469e-38, 5.063658e-38, 
    5.061848e-38, 5.083174e-38, 5.076309e-38, 5.12852e-38, 5.100091e-38, 
    5.181727e-38, 5.212149e-38, 5.299792e-38, 5.355955e-38, 5.414963e-38, 
    5.44214e-38, 5.450512e-38, 5.454017e-38,
  2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.522337e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.382207e-44, 2.522337e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.662467e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.522337e-44, 2.522337e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.662467e-44, 
    2.522337e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.522337e-44, 2.382207e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.662467e-44, 2.662467e-44, 2.802597e-44, 2.662467e-44, 2.382207e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 2.662467e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 2.802597e-44, 
    2.802597e-44, 2.802597e-44, 2.802597e-44,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_CH4_UNSAT =
  6.778707e-06, 7.045752e-06, 6.99349e-06, 7.211447e-06, 7.090201e-06, 
    7.233422e-06, 6.832496e-06, 7.056428e-06, 6.913117e-06, 6.802588e-06, 
    7.642347e-06, 7.221242e-06, 8.085404e-06, 7.810525e-06, 8.507648e-06, 
    8.042357e-06, 8.602514e-06, 8.494157e-06, 8.821607e-06, 8.727447e-06, 
    9.149589e-06, 8.865151e-06, 9.370066e-06, 9.081518e-06, 9.126532e-06, 
    8.855794e-06, 7.305245e-06, 7.589379e-06, 7.28854e-06, 7.328749e-06, 
    7.310707e-06, 7.092679e-06, 6.983857e-06, 6.758521e-06, 6.799192e-06, 
    6.964834e-06, 7.346861e-06, 7.216233e-06, 7.5474e-06, 7.539856e-06, 
    7.911418e-06, 7.741883e-06, 8.380981e-06, 8.197454e-06, 8.731374e-06, 
    8.596113e-06, 8.724997e-06, 8.685865e-06, 8.725508e-06, 8.527384e-06, 
    8.612105e-06, 8.438396e-06, 7.77351e-06, 7.966776e-06, 7.397875e-06, 
    7.06167e-06, 6.842241e-06, 6.688384e-06, 6.710038e-06, 6.751397e-06, 
    6.965807e-06, 7.170143e-06, 7.32755e-06, 7.433632e-06, 7.53877e-06, 
    7.856732e-06, 8.02858e-06, 8.418232e-06, 8.347484e-06, 8.467484e-06, 
    8.582691e-06, 8.777074e-06, 8.745003e-06, 8.830922e-06, 8.464343e-06, 
    8.707468e-06, 8.307265e-06, 8.41613e-06, 7.567282e-06, 7.251385e-06, 
    7.118678e-06, 7.003517e-06, 6.726706e-06, 6.917323e-06, 6.841889e-06, 
    7.021989e-06, 7.137473e-06, 7.080261e-06, 7.436542e-06, 7.297147e-06, 
    8.038812e-06, 7.715173e-06, 8.569231e-06, 8.361993e-06, 8.619141e-06, 
    8.487629e-06, 8.713312e-06, 8.51012e-06, 8.862968e-06, 8.940277e-06, 
    8.887425e-06, 9.090892e-06, 8.498893e-06, 8.724979e-06, 7.078653e-06, 
    7.087968e-06, 7.131457e-06, 6.941159e-06, 6.929601e-06, 6.757399e-06, 
    6.910544e-06, 6.976211e-06, 7.144206e-06, 7.244355e-06, 7.340116e-06, 
    7.552489e-06, 7.789039e-06, 8.128316e-06, 8.375375e-06, 8.542354e-06, 
    8.439853e-06, 8.530326e-06, 8.429201e-06, 8.381943e-06, 8.911279e-06, 
    8.612885e-06, 9.061566e-06, 9.036604e-06, 8.83296e-06, 9.039416e-06, 
    7.094515e-06, 7.040956e-06, 6.856337e-06, 7.000634e-06, 6.738767e-06, 
    6.884775e-06, 6.969351e-06, 7.300012e-06, 7.373575e-06, 7.442006e-06, 
    7.577951e-06, 7.750523e-06, 8.061662e-06, 8.336137e-06, 8.589417e-06, 
    8.570782e-06, 8.57734e-06, 8.634195e-06, 8.493542e-06, 8.657354e-06, 
    8.684918e-06, 8.612872e-06, 9.033261e-06, 8.912655e-06, 9.036073e-06, 
    8.957503e-06, 7.058351e-06, 7.148677e-06, 7.099803e-06, 7.191818e-06, 
    7.126926e-06, 7.417328e-06, 7.50533e-06, 7.918684e-06, 7.747049e-06, 
    8.020955e-06, 7.774712e-06, 7.818112e-06, 8.029877e-06, 7.787952e-06, 
    8.320885e-06, 7.958044e-06, 8.636408e-06, 8.26929e-06, 8.659571e-06, 
    8.588316e-06, 8.706401e-06, 8.812515e-06, 8.946509e-06, 9.194863e-06, 
    9.13724e-06, 9.345686e-06, 7.284266e-06, 7.403077e-06, 7.392617e-06, 
    7.517747e-06, 7.610824e-06, 7.810617e-06, 8.139795e-06, 8.015409e-06, 
    8.244335e-06, 8.290557e-06, 7.943013e-06, 8.155724e-06, 7.483057e-06, 
    7.590919e-06, 7.526648e-06, 7.293591e-06, 8.043963e-06, 7.657317e-06, 
    8.379473e-06, 8.16424e-06, 8.79736e-06, 8.480611e-06, 9.105541e-06, 
    9.375552e-06, 9.630785e-06, 9.929371e-06, 7.468288e-06, 7.387176e-06, 
    7.532694e-06, 7.732599e-06, 7.922341e-06, 8.177306e-06, 8.203579e-06, 
    8.251718e-06, 8.376906e-06, 8.482627e-06, 8.266928e-06, 8.5092e-06, 
    7.615955e-06, 8.078148e-06, 7.356574e-06, 7.57233e-06, 7.720629e-06, 
    7.657247e-06, 8.001247e-06, 8.083875e-06, 8.422764e-06, 8.246992e-06, 
    9.308763e-06, 8.834923e-06, 1.01567e-05, 9.78599e-06, 7.358913e-06, 
    7.468024e-06, 7.849024e-06, 7.668727e-06, 8.19445e-06, 8.326583e-06, 
    8.434554e-06, 8.573163e-06, 8.588193e-06, 8.670686e-06, 8.535625e-06, 
    8.665353e-06, 8.177852e-06, 8.39458e-06, 7.804877e-06, 7.946897e-06, 
    7.881448e-06, 7.809878e-06, 8.031585e-06, 8.270301e-06, 8.275482e-06, 
    8.352556e-06, 8.570895e-06, 8.19662e-06, 9.37014e-06, 8.640316e-06, 
    7.587739e-06, 7.79749e-06, 7.828085e-06, 7.745388e-06, 8.313302e-06, 
    8.105779e-06, 8.66868e-06, 8.515363e-06, 8.766991e-06, 8.641685e-06, 
    8.62329e-06, 8.463236e-06, 8.36405e-06, 8.115242e-06, 7.914849e-06, 
    7.757366e-06, 7.793874e-06, 7.967259e-06, 8.284996e-06, 8.589531e-06, 
    8.522517e-06, 8.747797e-06, 8.155663e-06, 8.402307e-06, 8.306661e-06, 
    8.556801e-06, 8.012101e-06, 8.475025e-06, 7.895287e-06, 7.94552e-06, 
    8.101679e-06, 8.419089e-06, 8.489946e-06, 8.565708e-06, 8.518946e-06, 
    8.293129e-06, 8.256351e-06, 8.097883e-06, 8.0543e-06, 7.934577e-06, 
    7.835962e-06, 7.926031e-06, 8.02104e-06, 8.293247e-06, 8.541183e-06, 
    8.81402e-06, 8.881159e-06, 9.203038e-06, 8.940749e-06, 9.374225e-06, 
    9.005317e-06, 9.645272e-06, 8.502197e-06, 8.994626e-06, 8.10883e-06, 
    8.202852e-06, 8.37382e-06, 8.770279e-06, 8.555619e-06, 8.806834e-06, 
    8.254916e-06, 7.973241e-06, 7.901031e-06, 7.766894e-06, 7.904107e-06, 
    7.892914e-06, 8.025023e-06, 7.98248e-06, 8.302341e-06, 8.129959e-06, 
    8.622813e-06, 8.804855e-06, 9.323785e-06, 9.644187e-06, 9.971066e-06, 
    1.011527e-05, 1.015913e-05, 1.017745e-05,
  7.386523e-06, 7.258159e-06, 7.282782e-06, 7.181714e-06, 7.237423e-06, 
    7.171761e-06, 7.360163e-06, 7.25315e-06, 7.321124e-06, 7.374798e-06, 
    6.994268e-06, 7.177274e-06, 6.519998e-06, 6.592286e-06, 6.419202e-06, 
    6.53096e-06, 6.398232e-06, 6.422246e-06, 6.352116e-06, 6.371545e-06, 
    6.289024e-06, 6.34333e-06, 6.250636e-06, 6.301538e-06, 6.293231e-06, 
    6.345206e-06, 7.139539e-06, 7.01642e-06, 7.146995e-06, 7.12908e-06, 
    7.137106e-06, 7.236262e-06, 7.287321e-06, 7.396505e-06, 7.376465e-06, 
    7.296377e-06, 7.121057e-06, 7.179561e-06, 7.034228e-06, 7.037432e-06, 
    6.565139e-06, 6.611176e-06, 6.448169e-06, 6.492071e-06, 6.370723e-06, 
    6.399637e-06, 6.372057e-06, 6.380315e-06, 6.37195e-06, 6.414799e-06, 
    6.396152e-06, 6.434911e-06, 6.602429e-06, 6.550546e-06, 7.098635e-06, 
    7.250674e-06, 7.355407e-06, 7.431411e-06, 7.420584e-06, 7.400018e-06, 
    7.295913e-06, 7.200558e-06, 7.129629e-06, 7.083062e-06, 7.037893e-06, 
    6.579739e-06, 6.534503e-06, 6.439534e-06, 6.456011e-06, 6.428272e-06, 
    6.402574e-06, 6.361228e-06, 6.367876e-06, 6.350221e-06, 6.428992e-06, 
    6.375738e-06, 6.465529e-06, 6.440026e-06, 7.025729e-06, 7.163673e-06, 
    7.224186e-06, 7.278036e-06, 7.412278e-06, 7.319092e-06, 7.355575e-06, 
    7.269337e-06, 7.215555e-06, 7.242054e-06, 7.0818e-06, 7.143155e-06, 
    6.531876e-06, 6.618609e-06, 6.40553e-06, 6.452605e-06, 6.394629e-06, 
    6.423721e-06, 6.374509e-06, 6.418663e-06, 6.343765e-06, 6.328462e-06, 
    6.33888e-06, 6.299804e-06, 6.421183e-06, 6.372057e-06, 7.242799e-06, 
    7.238463e-06, 7.218331e-06, 7.30767e-06, 7.313205e-06, 7.397055e-06, 
    7.322361e-06, 7.290972e-06, 7.212463e-06, 7.166841e-06, 7.124055e-06, 
    7.032063e-06, 6.598156e-06, 6.5092e-06, 6.449477e-06, 6.411473e-06, 
    6.43458e-06, 6.414148e-06, 6.437021e-06, 6.44795e-06, 6.334154e-06, 
    6.395981e-06, 6.305267e-06, 6.309963e-06, 6.349807e-06, 6.309432e-06, 
    7.235421e-06, 7.260425e-06, 7.348555e-06, 7.279413e-06, 7.40629e-06, 
    7.334775e-06, 7.294221e-06, 7.141858e-06, 7.109303e-06, 7.079422e-06, 
    7.021305e-06, 6.60878e-06, 6.52604e-06, 6.458679e-06, 6.401103e-06, 
    6.405191e-06, 6.40375e-06, 6.391372e-06, 6.422386e-06, 6.386393e-06, 
    6.380511e-06, 6.395988e-06, 6.310595e-06, 6.333889e-06, 6.310063e-06, 
    6.325115e-06, 7.252278e-06, 7.210402e-06, 7.232969e-06, 7.190654e-06, 
    7.22041e-06, 7.090129e-06, 7.052121e-06, 6.5632e-06, 6.60974e-06, 
    6.536474e-06, 6.602102e-06, 6.59022e-06, 6.534157e-06, 6.598466e-06, 
    6.462278e-06, 6.552819e-06, 6.390894e-06, 6.474588e-06, 6.385918e-06, 
    6.401344e-06, 6.37597e-06, 6.353962e-06, 6.327252e-06, 6.280887e-06, 
    6.291282e-06, 6.254729e-06, 7.148913e-06, 7.096357e-06, 7.10095e-06, 
    7.046844e-06, 7.007488e-06, 6.592267e-06, 6.506337e-06, 6.537914e-06, 
    6.480638e-06, 6.46951e-06, 6.556792e-06, 6.502368e-06, 7.061693e-06, 
    7.015818e-06, 7.043041e-06, 7.144733e-06, 6.530558e-06, 6.988099e-06, 
    6.44852e-06, 6.500261e-06, 6.357058e-06, 6.425295e-06, 6.297093e-06, 
    6.249713e-06, 6.209385e-06, 6.167667e-06, 7.068059e-06, 7.103335e-06, 
    7.040477e-06, 6.613744e-06, 6.562243e-06, 6.497027e-06, 6.490569e-06, 
    6.478848e-06, 6.449123e-06, 6.42485e-06, 6.47517e-06, 6.41887e-06, 
    7.005285e-06, 6.521846e-06, 7.116779e-06, 7.023645e-06, 6.617085e-06, 
    6.988147e-06, 6.541581e-06, 6.520403e-06, 6.438492e-06, 6.479995e-06, 
    6.260979e-06, 6.349401e-06, 6.139932e-06, 6.186955e-06, 7.115758e-06, 
    7.068181e-06, 6.581838e-06, 6.983395e-06, 6.492809e-06, 6.46094e-06, 
    6.435794e-06, 6.404662e-06, 6.401369e-06, 6.383541e-06, 6.412969e-06, 
    6.384683e-06, 6.496893e-06, 6.44501e-06, 6.593836e-06, 6.555764e-06, 
    6.573135e-06, 6.592471e-06, 6.533749e-06, 6.474357e-06, 6.473124e-06, 
    6.454814e-06, 6.405121e-06, 6.492276e-06, 6.250595e-06, 6.390015e-06, 
    7.017185e-06, 6.595835e-06, 6.587512e-06, 6.610207e-06, 6.464089e-06, 
    6.514866e-06, 6.383971e-06, 6.417489e-06, 6.363313e-06, 6.389758e-06, 
    6.393729e-06, 6.429245e-06, 6.452124e-06, 6.512483e-06, 6.564228e-06, 
    6.606891e-06, 6.596844e-06, 6.550421e-06, 6.470832e-06, 6.401072e-06, 
    6.415881e-06, 6.367296e-06, 6.502391e-06, 6.443214e-06, 6.465662e-06, 
    6.408272e-06, 6.538766e-06, 6.426531e-06, 6.569438e-06, 6.556131e-06, 
    6.515899e-06, 6.439331e-06, 6.423198e-06, 6.406303e-06, 6.416687e-06, 
    6.468889e-06, 6.477727e-06, 6.51686e-06, 6.527922e-06, 6.559016e-06, 
    6.585381e-06, 6.56127e-06, 6.536455e-06, 6.468867e-06, 6.411727e-06, 
    6.353654e-06, 6.340131e-06, 6.279414e-06, 6.328357e-06, 6.249913e-06, 
    6.315861e-06, 6.2072e-06, 6.420417e-06, 6.317928e-06, 6.514102e-06, 
    6.490748e-06, 6.449829e-06, 6.362618e-06, 6.408533e-06, 6.355112e-06, 
    6.478075e-06, 6.548851e-06, 6.567906e-06, 6.604257e-06, 6.567087e-06, 
    6.57007e-06, 6.535438e-06, 6.546457e-06, 6.466697e-06, 6.5088e-06, 
    6.393829e-06, 6.355519e-06, 6.258431e-06, 6.207376e-06, 6.162328e-06, 
    6.144731e-06, 6.139659e-06, 6.137578e-06,
  9.864346e-06, 9.872007e-06, 9.870747e-06, 9.875229e-06, 9.872987e-06, 
    9.875568e-06, 9.866133e-06, 9.872249e-06, 9.868581e-06, 9.865154e-06, 
    9.878062e-06, 9.875383e-06, 1.019394e-05, 1.024211e-05, 1.011908e-05, 
    1.02015e-05, 1.01021e-05, 1.012151e-05, 1.00626e-05, 1.007963e-05, 
    1.000262e-05, 1.00547e-05, 9.961702e-06, 1.001516e-05, 1.000688e-05, 
    1.00564e-05, 9.876531e-06, 9.878147e-06, 9.876328e-06, 9.876797e-06, 
    9.876595e-06, 9.873039e-06, 9.870501e-06, 9.863644e-06, 9.865041e-06, 
    9.870007e-06, 9.876986e-06, 9.875305e-06, 9.878137e-06, 9.878125e-06, 
    1.022448e-05, 1.025408e-05, 1.014168e-05, 1.017421e-05, 1.007893e-05, 
    1.010326e-05, 1.008007e-05, 1.008713e-05, 1.007998e-05, 1.011557e-05, 
    1.010039e-05, 1.013146e-05, 1.024856e-05, 1.021478e-05, 9.877444e-06, 
    9.872366e-06, 9.866444e-06, 9.861068e-06, 9.861886e-06, 9.863391e-06, 
    9.870032e-06, 9.874537e-06, 9.876786e-06, 9.877698e-06, 9.878123e-06, 
    1.023401e-05, 1.020393e-05, 1.013504e-05, 1.014764e-05, 1.012627e-05, 
    1.010567e-05, 1.007066e-05, 1.007646e-05, 1.006091e-05, 1.012684e-05, 
    1.008323e-05, 1.015478e-05, 1.013543e-05, 9.878146e-06, 9.87583e-06, 
    9.873568e-06, 9.870998e-06, 9.862501e-06, 9.868701e-06, 9.866432e-06, 
    9.871449e-06, 9.873937e-06, 9.872776e-06, 9.877716e-06, 9.876434e-06, 
    1.020213e-05, 1.025872e-05, 1.010808e-05, 1.014506e-05, 1.009913e-05, 
    1.012268e-05, 1.008218e-05, 1.011866e-05, 1.005509e-05, 1.004102e-05, 
    1.005065e-05, 1.001345e-05, 1.012067e-05, 1.008007e-05, 9.872741e-06, 
    9.872941e-06, 9.873822e-06, 9.869368e-06, 9.869048e-06, 9.863604e-06, 
    9.868508e-06, 9.870305e-06, 9.874065e-06, 9.87573e-06, 9.876919e-06, 
    9.878142e-06, 1.024585e-05, 1.018639e-05, 1.014268e-05, 1.01129e-05, 
    1.013121e-05, 1.011505e-05, 1.01331e-05, 1.014152e-05, 1.00463e-05, 
    1.010025e-05, 1.001884e-05, 1.002342e-05, 1.006054e-05, 1.00229e-05, 
    9.873078e-06, 9.871897e-06, 9.866886e-06, 9.870927e-06, 9.862939e-06, 
    9.867752e-06, 9.870125e-06, 9.876468e-06, 9.877242e-06, 9.877749e-06, 
    9.878157e-06, 1.025257e-05, 1.019812e-05, 1.014964e-05, 1.010447e-05, 
    1.010781e-05, 1.010663e-05, 1.009642e-05, 1.012162e-05, 1.009226e-05, 
    1.008729e-05, 1.010025e-05, 1.002403e-05, 1.004606e-05, 1.002351e-05, 
    1.003789e-05, 9.872294e-06, 9.874148e-06, 9.873188e-06, 9.87491e-06, 
    9.873733e-06, 9.877587e-06, 9.878037e-06, 1.022319e-05, 1.025317e-05, 
    1.020527e-05, 1.024836e-05, 1.024078e-05, 1.020368e-05, 1.024605e-05, 
    1.015234e-05, 1.021629e-05, 1.009603e-05, 1.016147e-05, 1.009186e-05, 
    1.010466e-05, 1.008343e-05, 1.006425e-05, 1.003989e-05, 9.994272e-06, 
    1.000491e-05, 9.966263e-06, 9.876274e-06, 9.877484e-06, 9.877403e-06, 
    9.878076e-06, 9.878136e-06, 1.02421e-05, 1.018437e-05, 1.020626e-05, 
    1.016592e-05, 1.015773e-05, 1.021896e-05, 1.018156e-05, 9.877956e-06, 
    9.878151e-06, 9.878097e-06, 9.876389e-06, 1.020123e-05, 9.878021e-06, 
    1.014195e-05, 1.018007e-05, 1.006699e-05, 1.012392e-05, 1.001075e-05, 
    9.96066e-06, 9.912575e-06, 9.855148e-06, 9.877891e-06, 9.877359e-06, 
    9.878111e-06, 1.025568e-05, 1.022257e-05, 1.017776e-05, 1.017313e-05, 
    1.016461e-05, 1.014241e-05, 1.012357e-05, 1.016191e-05, 1.011883e-05, 
    9.878121e-06, 1.019522e-05, 9.877082e-06, 9.878153e-06, 1.025777e-05, 
    9.878024e-06, 1.020875e-05, 1.019423e-05, 1.013424e-05, 1.016545e-05, 
    9.973116e-06, 1.006017e-05, 9.810544e-06, 9.882879e-06, 9.877106e-06, 
    9.87789e-06, 1.023538e-05, 9.877983e-06, 1.017474e-05, 1.015134e-05, 
    1.013215e-05, 1.010737e-05, 1.010468e-05, 1.008986e-05, 1.01141e-05, 
    1.009082e-05, 1.017766e-05, 1.013927e-05, 1.02431e-05, 1.021827e-05, 
    1.022973e-05, 1.024223e-05, 1.020342e-05, 1.016131e-05, 1.016041e-05, 
    1.014673e-05, 1.010772e-05, 1.017435e-05, 9.961633e-06, 1.009527e-05, 
    9.878157e-06, 1.024437e-05, 1.023905e-05, 1.025347e-05, 1.01537e-05, 
    1.019037e-05, 1.009022e-05, 1.011773e-05, 1.007249e-05, 1.009508e-05, 
    1.009838e-05, 1.012704e-05, 1.014469e-05, 1.01887e-05, 1.022388e-05, 
    1.025138e-05, 1.024502e-05, 1.02147e-05, 1.015871e-05, 1.010444e-05, 
    1.011644e-05, 1.007596e-05, 1.018158e-05, 1.013788e-05, 1.015487e-05, 
    1.011031e-05, 1.020684e-05, 1.012488e-05, 1.022731e-05, 1.021852e-05, 
    1.019109e-05, 1.013488e-05, 1.012227e-05, 1.010871e-05, 1.011709e-05, 
    1.015727e-05, 1.016379e-05, 1.019176e-05, 1.019942e-05, 1.022043e-05, 
    1.023768e-05, 1.022193e-05, 1.020526e-05, 1.015726e-05, 1.01131e-05, 
    1.006397e-05, 1.005179e-05, 9.99273e-06, 1.004091e-05, 9.960866e-06, 
    1.002907e-05, 9.909768e-06, 1.012005e-05, 1.003106e-05, 1.018984e-05, 
    1.017325e-05, 1.014294e-05, 1.007187e-05, 1.011052e-05, 1.006526e-05, 
    1.016404e-05, 1.021364e-05, 1.02263e-05, 1.024972e-05, 1.022577e-05, 
    1.022772e-05, 1.020457e-05, 1.021204e-05, 1.015564e-05, 1.018611e-05, 
    1.009846e-05, 1.006562e-05, 9.97034e-06, 9.910005e-06, 9.847054e-06, 
    9.818749e-06, 9.810073e-06, 9.806437e-06,
  4.318993e-06, 4.232694e-06, 4.249457e-06, 4.179964e-06, 4.218499e-06, 
    4.173017e-06, 4.301485e-06, 4.229268e-06, 4.275356e-06, 4.311221e-06, 
    4.045519e-06, 4.176868e-06, 3.910047e-06, 3.993352e-06, 3.784661e-06, 
    3.922987e-06, 3.756878e-06, 3.788648e-06, 3.693203e-06, 3.7205e-06, 
    3.598924e-06, 3.680618e-06, 3.536246e-06, 3.618404e-06, 3.605522e-06, 
    3.683318e-06, 4.150398e-06, 4.061837e-06, 4.15565e-06, 4.143004e-06, 
    4.148681e-06, 4.217699e-06, 4.252528e-06, 4.325603e-06, 4.312328e-06, 
    4.258664e-06, 4.13732e-06, 4.178467e-06, 4.074887e-06, 4.077223e-06, 
    3.962622e-06, 4.014381e-06, 3.821999e-06, 3.87652e-06, 3.71936e-06, 
    3.75877e-06, 3.721208e-06, 3.732591e-06, 3.721059e-06, 3.778891e-06, 
    3.754092e-06, 3.805058e-06, 4.004678e-06, 3.945835e-06, 4.121362e-06, 
    4.227568e-06, 4.298313e-06, 4.348586e-06, 4.341475e-06, 4.327921e-06, 
    4.258351e-06, 4.193068e-06, 4.143399e-06, 4.110217e-06, 4.077559e-06, 
    3.97921e-06, 3.927151e-06, 3.810986e-06, 3.831913e-06, 3.79648e-06, 
    3.762696e-06, 3.706092e-06, 3.715398e-06, 3.690499e-06, 3.797419e-06, 
    3.726293e-06, 3.843841e-06, 3.811623e-06, 4.068656e-06, 4.167363e-06, 
    4.209385e-06, 4.246233e-06, 4.336008e-06, 4.273987e-06, 4.298424e-06, 
    4.240319e-06, 4.203443e-06, 4.221678e-06, 4.10931e-06, 4.152948e-06, 
    3.924069e-06, 4.022573e-06, 3.766633e-06, 3.827617e-06, 3.752044e-06, 
    3.790574e-06, 3.724597e-06, 3.783966e-06, 3.681243e-06, 3.658944e-06, 
    3.674179e-06, 3.615738e-06, 3.787262e-06, 3.721205e-06, 4.222188e-06, 
    4.219213e-06, 4.205361e-06, 4.266292e-06, 4.270024e-06, 4.325965e-06, 
    4.276188e-06, 4.255008e-06, 4.201309e-06, 4.16958e-06, 4.13945e-06, 
    4.073305e-06, 3.999912e-06, 3.897183e-06, 3.823658e-06, 3.774511e-06, 
    3.804636e-06, 3.778037e-06, 3.807772e-06, 3.821725e-06, 3.667294e-06, 
    3.753859e-06, 3.624132e-06, 3.631287e-06, 3.689906e-06, 3.630481e-06, 
    4.217125e-06, 4.234245e-06, 4.293739e-06, 4.247172e-06, 4.332062e-06, 
    4.284518e-06, 4.257204e-06, 4.152028e-06, 4.128973e-06, 4.1076e-06, 
    4.065439e-06, 4.011729e-06, 3.917202e-06, 3.835263e-06, 3.760733e-06, 
    3.766185e-06, 3.764265e-06, 3.747647e-06, 3.788833e-06, 3.740893e-06, 
    3.732856e-06, 3.753873e-06, 3.632246e-06, 3.666913e-06, 3.63144e-06, 
    3.654004e-06, 4.22868e-06, 4.199883e-06, 4.21544e-06, 4.18619e-06, 
    4.206792e-06, 4.115275e-06, 4.087889e-06, 3.960395e-06, 4.01279e-06, 
    3.929462e-06, 4.004316e-06, 3.991035e-06, 3.926736e-06, 4.000267e-06, 
    3.839767e-06, 3.948453e-06, 3.747001e-06, 3.855067e-06, 3.740247e-06, 
    3.761055e-06, 3.726619e-06, 3.695826e-06, 3.657164e-06, 3.586034e-06, 
    3.602481e-06, 3.543169e-06, 4.157002e-06, 4.119735e-06, 4.123019e-06, 
    4.084067e-06, 4.055292e-06, 3.993335e-06, 3.893753e-06, 3.931154e-06, 
    3.862544e-06, 3.848792e-06, 3.953049e-06, 3.888977e-06, 4.094823e-06, 
    4.061409e-06, 4.081303e-06, 4.154057e-06, 3.922522e-06, 4.040965e-06, 
    3.822444e-06, 3.88644e-06, 3.700213e-06, 3.792613e-06, 3.611539e-06, 
    3.534669e-06, 3.462681e-06, 3.378955e-06, 4.09942e-06, 4.12472e-06, 
    4.07944e-06, 4.017209e-06, 3.959308e-06, 3.88253e-06, 3.874692e-06, 
    3.860339e-06, 3.823213e-06, 3.792043e-06, 3.855798e-06, 3.784238e-06, 
    4.053653e-06, 3.912243e-06, 4.134286e-06, 4.067144e-06, 4.020896e-06, 
    4.041005e-06, 3.935435e-06, 3.91054e-06, 3.809654e-06, 3.861753e-06, 
    3.553603e-06, 3.68932e-06, 3.315555e-06, 3.419086e-06, 4.133564e-06, 
    4.099511e-06, 3.981596e-06, 4.037481e-06, 3.877417e-06, 3.838101e-06, 
    3.806197e-06, 3.765475e-06, 3.761088e-06, 3.737005e-06, 3.776484e-06, 
    3.738565e-06, 3.882367e-06, 3.817986e-06, 3.995094e-06, 3.951863e-06, 
    3.971743e-06, 3.993564e-06, 3.926279e-06, 3.854791e-06, 3.853275e-06, 
    3.8304e-06, 3.766055e-06, 3.876769e-06, 3.536148e-06, 3.745781e-06, 
    4.062421e-06, 3.997317e-06, 3.987996e-06, 4.013311e-06, 3.842039e-06, 
    3.903955e-06, 3.737592e-06, 3.782427e-06, 3.709021e-06, 3.745464e-06, 
    3.75083e-06, 3.797747e-06, 3.827009e-06, 3.901111e-06, 3.96158e-06, 
    4.00964e-06, 3.998457e-06, 3.945693e-06, 3.850428e-06, 3.760686e-06, 
    3.78031e-06, 3.714591e-06, 3.88901e-06, 3.815692e-06, 3.843998e-06, 
    3.770273e-06, 3.932147e-06, 3.794198e-06, 3.967536e-06, 3.952289e-06, 
    3.905186e-06, 3.810722e-06, 3.789892e-06, 3.767657e-06, 3.781377e-06, 
    3.848016e-06, 3.858957e-06, 3.906332e-06, 3.919424e-06, 3.955608e-06, 
    3.985601e-06, 3.958194e-06, 3.929442e-06, 3.847992e-06, 3.77484e-06, 
    3.695387e-06, 3.675996e-06, 3.583662e-06, 3.658777e-06, 3.534986e-06, 
    3.640156e-06, 3.458536e-06, 3.786245e-06, 3.643277e-06, 3.903047e-06, 
    3.87491e-06, 3.824097e-06, 3.708033e-06, 3.77062e-06, 3.69745e-06, 
    3.859387e-06, 3.94387e-06, 3.965788e-06, 4.006713e-06, 3.964853e-06, 
    3.968256e-06, 3.928259e-06, 3.941105e-06, 3.845293e-06, 3.89671e-06, 
    3.750963e-06, 3.698029e-06, 3.549372e-06, 3.458884e-06, 3.367343e-06, 
    3.327112e-06, 3.314892e-06, 3.309786e-06,
  4.42685e-07, 4.259929e-07, 4.292083e-07, 4.159626e-07, 4.232802e-07, 
    4.146509e-07, 4.392707e-07, 4.253374e-07, 4.342017e-07, 4.411676e-07, 
    3.909649e-07, 4.153777e-07, 3.665589e-07, 3.814325e-07, 3.447602e-07, 
    3.688487e-07, 3.400254e-07, 3.454425e-07, 3.293033e-07, 3.338776e-07, 
    3.137583e-07, 3.272055e-07, 3.036412e-07, 3.169381e-07, 3.148335e-07, 
    3.27655e-07, 4.103944e-07, 3.93955e-07, 4.113809e-07, 4.090084e-07, 
    4.100723e-07, 4.231277e-07, 4.297989e-07, 4.439777e-07, 4.413835e-07, 
    4.3098e-07, 4.079443e-07, 4.156799e-07, 3.963551e-07, 3.967854e-07, 
    3.759094e-07, 3.852367e-07, 3.511778e-07, 3.606609e-07, 3.336859e-07, 
    3.403467e-07, 3.339967e-07, 3.359145e-07, 3.339718e-07, 3.437741e-07, 
    3.395525e-07, 3.482584e-07, 3.834789e-07, 3.729102e-07, 4.049652e-07, 
    4.250123e-07, 4.386537e-07, 4.484883e-07, 4.470901e-07, 4.444315e-07, 
    4.309196e-07, 4.184433e-07, 4.090822e-07, 4.028913e-07, 3.968472e-07, 
    3.788854e-07, 3.695871e-07, 3.492785e-07, 3.528924e-07, 3.467849e-07, 
    3.410139e-07, 3.314591e-07, 3.330202e-07, 3.28852e-07, 3.469461e-07, 
    3.348526e-07, 3.549609e-07, 3.493882e-07, 3.952081e-07, 4.135846e-07, 
    4.215434e-07, 4.285889e-07, 4.460167e-07, 4.339369e-07, 4.386752e-07, 
    4.27454e-07, 4.204131e-07, 4.238869e-07, 4.027228e-07, 4.108732e-07, 
    3.690404e-07, 3.867241e-07, 3.416839e-07, 3.521489e-07, 3.39205e-07, 
    3.457725e-07, 3.345671e-07, 3.446414e-07, 3.273095e-07, 3.236091e-07, 
    3.261348e-07, 3.165018e-07, 3.452053e-07, 3.339962e-07, 4.239843e-07, 
    4.234164e-07, 4.207776e-07, 4.324507e-07, 4.331713e-07, 4.440486e-07, 
    4.343626e-07, 4.30276e-07, 4.200076e-07, 4.140026e-07, 4.083427e-07, 
    3.960636e-07, 3.826171e-07, 3.642898e-07, 3.514645e-07, 3.430265e-07, 
    3.481858e-07, 3.436283e-07, 3.487253e-07, 3.511306e-07, 3.249922e-07, 
    3.39513e-07, 3.178761e-07, 3.190501e-07, 3.28753e-07, 3.189177e-07, 
    4.230181e-07, 4.262899e-07, 4.377649e-07, 4.287693e-07, 4.452429e-07, 
    4.359755e-07, 4.306988e-07, 4.107006e-07, 4.063845e-07, 4.024052e-07, 
    3.946168e-07, 3.847559e-07, 3.678241e-07, 3.534726e-07, 3.406803e-07, 
    3.416077e-07, 3.41281e-07, 3.384597e-07, 3.454742e-07, 3.373168e-07, 
    3.359591e-07, 3.395153e-07, 3.192075e-07, 3.24929e-07, 3.190751e-07, 
    3.227923e-07, 4.252249e-07, 4.197367e-07, 4.226969e-07, 4.171404e-07, 
    4.210499e-07, 4.038318e-07, 3.987538e-07, 3.755108e-07, 3.849482e-07, 
    3.699973e-07, 3.834134e-07, 3.810145e-07, 3.695135e-07, 3.826813e-07, 
    3.542537e-07, 3.733772e-07, 3.383504e-07, 3.569138e-07, 3.372075e-07, 
    3.40735e-07, 3.349076e-07, 3.297414e-07, 3.233145e-07, 3.116635e-07, 
    3.143376e-07, 3.047501e-07, 4.116347e-07, 4.046619e-07, 4.05274e-07, 
    3.98048e-07, 3.927543e-07, 3.814294e-07, 3.636862e-07, 3.702978e-07, 
    3.582173e-07, 3.558216e-07, 3.741976e-07, 3.628464e-07, 4.000363e-07, 
    3.938763e-07, 3.975377e-07, 4.110815e-07, 3.687663e-07, 3.901324e-07, 
    3.512547e-07, 3.624008e-07, 3.304748e-07, 3.461218e-07, 3.158156e-07, 
    3.033889e-07, 2.91987e-07, 2.790114e-07, 4.008879e-07, 4.055912e-07, 
    3.971942e-07, 3.857499e-07, 3.753163e-07, 3.617145e-07, 3.603409e-07, 
    3.578327e-07, 3.513875e-07, 3.460242e-07, 3.57041e-07, 3.446879e-07, 
    3.924539e-07, 3.669469e-07, 4.07377e-07, 3.949301e-07, 3.864193e-07, 
    3.901399e-07, 3.710584e-07, 3.666459e-07, 3.490491e-07, 3.580793e-07, 
    3.064256e-07, 3.286553e-07, 2.693892e-07, 2.851926e-07, 4.07242e-07, 
    4.009045e-07, 3.793146e-07, 3.894965e-07, 3.608181e-07, 3.539647e-07, 
    3.484543e-07, 3.414868e-07, 3.407406e-07, 3.366595e-07, 3.433631e-07, 
    3.369231e-07, 3.616859e-07, 3.50485e-07, 3.817468e-07, 3.739856e-07, 
    3.775443e-07, 3.814708e-07, 3.694323e-07, 3.568656e-07, 3.566016e-07, 
    3.526305e-07, 3.415855e-07, 3.607047e-07, 3.036255e-07, 3.381438e-07, 
    3.940622e-07, 3.821482e-07, 3.804667e-07, 3.850428e-07, 3.546481e-07, 
    3.654834e-07, 3.367589e-07, 3.443783e-07, 3.319501e-07, 3.3809e-07, 
    3.389992e-07, 3.470025e-07, 3.520436e-07, 3.649818e-07, 3.757228e-07, 
    3.843772e-07, 3.823542e-07, 3.728849e-07, 3.56106e-07, 3.406723e-07, 
    3.440165e-07, 3.328846e-07, 3.628522e-07, 3.500895e-07, 3.549883e-07, 
    3.423039e-07, 3.704741e-07, 3.463936e-07, 3.767896e-07, 3.740617e-07, 
    3.657005e-07, 3.492331e-07, 3.456556e-07, 3.418583e-07, 3.441987e-07, 
    3.556866e-07, 3.575917e-07, 3.659027e-07, 3.682174e-07, 3.746547e-07, 
    3.800353e-07, 3.75117e-07, 3.699938e-07, 3.556823e-07, 3.430827e-07, 
    3.29668e-07, 3.264367e-07, 3.112788e-07, 3.235814e-07, 3.034395e-07, 
    3.205083e-07, 2.913375e-07, 3.450312e-07, 3.210224e-07, 3.653234e-07, 
    3.603791e-07, 3.515403e-07, 3.317844e-07, 3.423629e-07, 3.300128e-07, 
    3.576666e-07, 3.725599e-07, 3.764764e-07, 3.838473e-07, 3.763089e-07, 
    3.769187e-07, 3.697837e-07, 3.720675e-07, 3.552132e-07, 3.642067e-07, 
    3.390217e-07, 3.301096e-07, 3.057455e-07, 2.91392e-07, 2.77236e-07, 
    2.711303e-07, 2.692895e-07, 2.685223e-07,
  1.244382e-08, 1.172625e-08, 1.186334e-08, 1.13022e-08, 1.161104e-08, 
    1.124714e-08, 1.229585e-08, 1.169838e-08, 1.20773e-08, 1.237798e-08, 
    1.026909e-08, 1.127763e-08, 9.293927e-09, 9.884218e-09, 8.45179e-09, 
    9.383982e-09, 8.272557e-09, 8.47773e-09, 7.871628e-09, 8.041829e-09, 
    7.30274e-09, 7.793995e-09, 6.945613e-09, 7.417901e-09, 7.341609e-09, 
    7.810605e-09, 1.106912e-08, 1.039086e-08, 1.111029e-08, 1.101137e-08, 
    1.105569e-08, 1.160457e-08, 1.188857e-08, 1.25e-08, 1.238734e-08, 
    1.19391e-08, 1.09671e-08, 1.129032e-08, 1.048896e-08, 1.050658e-08, 
    9.663556e-09, 1.00372e-08, 8.69684e-09, 9.063351e-09, 8.034672e-09, 
    8.284679e-09, 8.046277e-09, 8.118023e-09, 8.045346e-09, 8.414353e-09, 
    8.254728e-09, 8.585064e-09, 9.966413e-09, 9.544456e-09, 1.084349e-08, 
    1.168456e-08, 1.226917e-08, 1.269672e-08, 1.263563e-08, 1.251974e-08, 
    1.193651e-08, 1.140657e-08, 1.101444e-08, 1.075772e-08, 1.050911e-08, 
    9.782241e-09, 9.413085e-09, 8.624066e-09, 8.762718e-09, 8.528838e-09, 
    8.309868e-09, 7.951682e-09, 8.009832e-09, 7.854902e-09, 8.534985e-09, 
    8.07827e-09, 8.842425e-09, 8.628263e-09, 1.044204e-08, 1.120245e-08, 
    1.153748e-08, 1.183689e-08, 1.25888e-08, 1.206592e-08, 1.227011e-08, 
    1.178848e-08, 1.148969e-08, 1.163677e-08, 1.075076e-08, 1.10891e-08, 
    9.391536e-09, 1.009724e-08, 8.335189e-09, 8.734129e-09, 8.241637e-09, 
    8.490281e-09, 8.067595e-09, 8.447279e-09, 7.797835e-09, 7.661525e-09, 
    7.754475e-09, 7.402064e-09, 8.468707e-09, 8.04626e-09, 1.16409e-08, 
    1.161681e-08, 1.150509e-08, 1.200212e-08, 1.203304e-08, 1.250308e-08, 
    1.208422e-08, 1.190897e-08, 1.147256e-08, 1.121996e-08, 1.098367e-08, 
    1.047703e-08, 9.93177e-09, 9.204981e-09, 8.707842e-09, 8.386007e-09, 
    8.58229e-09, 8.408821e-09, 8.602906e-09, 8.695026e-09, 7.712376e-09, 
    8.25324e-09, 7.451992e-09, 7.494736e-09, 7.851238e-09, 7.489911e-09, 
    1.159992e-08, 1.17389e-08, 1.223078e-08, 1.184458e-08, 1.255507e-08, 
    1.215362e-08, 1.192706e-08, 1.108189e-08, 1.090232e-08, 1.073765e-08, 
    1.041787e-08, 1.001782e-08, 9.343648e-09, 8.78505e-09, 8.297268e-09, 
    8.332306e-09, 8.319957e-09, 8.213583e-09, 8.478933e-09, 8.170623e-09, 
    8.119696e-09, 8.253329e-09, 7.500474e-09, 7.710051e-09, 7.495647e-09, 
    7.631548e-09, 1.16936e-08, 1.146112e-08, 1.158631e-08, 1.135171e-08, 
    1.15166e-08, 1.079659e-08, 1.058732e-08, 9.647697e-09, 1.002558e-08, 
    9.429271e-09, 9.963778e-09, 9.867457e-09, 9.410184e-09, 9.934348e-09, 
    8.815145e-09, 9.562966e-09, 8.209469e-09, 8.917902e-09, 8.166521e-09, 
    8.299333e-09, 8.080328e-09, 7.887873e-09, 7.65071e-09, 7.227217e-09, 
    7.323673e-09, 6.979911e-09, 1.11209e-08, 1.083093e-08, 1.085628e-08, 
    1.055834e-08, 1.03419e-08, 9.884094e-09, 9.18137e-09, 9.441131e-09, 
    8.968407e-09, 8.875661e-09, 9.595515e-09, 9.148556e-09, 1.064004e-08, 
    1.038765e-08, 1.053741e-08, 1.109779e-08, 9.380738e-09, 1.023528e-08, 
    8.699791e-09, 9.13116e-09, 7.915095e-09, 8.50358e-09, 7.377177e-09, 
    6.936631e-09, 6.535179e-09, 6.088717e-09, 1.067509e-08, 1.086942e-08, 
    1.052333e-08, 1.00579e-08, 9.639963e-09, 9.104394e-09, 9.050896e-09, 
    8.953497e-09, 8.704887e-09, 8.499862e-09, 8.922826e-09, 8.449041e-09, 
    1.032967e-08, 9.309167e-09, 1.094352e-08, 1.043067e-08, 1.008493e-08, 
    1.023558e-08, 9.471173e-09, 9.297344e-09, 8.615288e-09, 8.963056e-09, 
    7.039572e-09, 7.847617e-09, 5.764934e-09, 6.300001e-09, 1.093792e-08, 
    1.067578e-08, 9.7994e-09, 1.020947e-08, 9.069469e-09, 8.804007e-09, 
    8.592549e-09, 8.327738e-09, 8.299545e-09, 8.145956e-09, 8.398764e-09, 
    8.155846e-09, 9.103278e-09, 8.67027e-09, 9.896827e-09, 9.587104e-09, 
    9.728696e-09, 9.885754e-09, 9.406985e-09, 8.916038e-09, 8.905824e-09, 
    8.752642e-09, 8.331465e-09, 9.065054e-09, 6.945051e-09, 8.201702e-09, 
    1.039523e-08, 9.91294e-09, 9.84551e-09, 1.002939e-08, 8.830354e-09, 
    9.251731e-09, 8.149682e-09, 8.437286e-09, 7.969954e-09, 8.199678e-09, 
    8.233888e-09, 8.537133e-09, 8.730084e-09, 9.232076e-09, 9.656132e-09, 
    1.000257e-08, 9.921211e-09, 9.543451e-09, 8.886655e-09, 8.296968e-09, 
    8.423551e-09, 8.004773e-09, 9.148784e-09, 8.655114e-09, 8.843479e-09, 
    8.358644e-09, 9.448092e-09, 8.513928e-09, 9.698608e-09, 9.590122e-09, 
    9.260244e-09, 8.622325e-09, 8.485836e-09, 8.341784e-09, 8.430467e-09, 
    8.870444e-09, 8.944157e-09, 9.268176e-09, 9.359124e-09, 9.61367e-09, 
    9.828235e-09, 9.63204e-09, 9.42913e-09, 8.870281e-09, 8.388136e-09, 
    7.885149e-09, 7.765612e-09, 7.213376e-09, 7.660507e-09, 6.938432e-09, 
    7.547944e-09, 6.512565e-09, 8.462089e-09, 7.566734e-09, 9.245459e-09, 
    9.052385e-09, 8.710752e-09, 7.963789e-09, 8.360877e-09, 7.897942e-09, 
    8.947058e-09, 9.530578e-09, 9.686132e-09, 9.981235e-09, 9.679462e-09, 
    9.703752e-09, 9.420841e-09, 9.511082e-09, 8.852161e-09, 9.201728e-09, 
    8.234734e-09, 7.901535e-09, 7.015334e-09, 6.514461e-09, 6.028502e-09, 
    5.823052e-09, 5.761612e-09, 5.736073e-09,
  8.583546e-11, 7.828845e-11, 7.971288e-11, 7.393521e-11, 7.709768e-11, 
    7.337598e-11, 8.426102e-11, 7.799981e-11, 8.195267e-11, 8.513381e-11, 
    6.367942e-11, 7.368555e-11, 5.448361e-11, 5.999168e-11, 4.695276e-11, 
    5.531204e-11, 4.540215e-11, 4.717873e-11, 4.200308e-11, 4.343415e-11, 
    3.73516e-11, 4.135626e-11, 3.139945e-11, 3.827646e-11, 3.766279e-11, 
    4.149434e-11, 7.157744e-11, 6.486158e-11, 7.199205e-11, 7.099707e-11, 
    7.144231e-11, 7.703103e-11, 7.997599e-11, 8.643568e-11, 8.523344e-11, 
    8.050371e-11, 7.055328e-11, 7.38145e-11, 6.581923e-11, 6.599175e-11, 
    5.791134e-11, 6.144864e-11, 4.910298e-11, 5.238247e-11, 4.337361e-11, 
    4.550643e-11, 4.347179e-11, 4.408051e-11, 4.34639e-11, 4.662732e-11, 
    4.524895e-11, 4.811791e-11, 6.077298e-11, 5.679899e-11, 6.931895e-11, 
    7.785685e-11, 8.397818e-11, 8.854785e-11, 8.789017e-11, 8.664695e-11, 
    8.047665e-11, 7.499915e-11, 7.102791e-11, 6.846679e-11, 6.601658e-11, 
    5.902714e-11, 5.558071e-11, 4.846081e-11, 4.968689e-11, 4.76251e-11, 
    4.572339e-11, 4.267397e-11, 4.316376e-11, 4.18634e-11, 4.767889e-11, 
    4.374285e-11, 5.039665e-11, 4.849778e-11, 6.536061e-11, 7.292315e-11, 
    7.63405e-11, 7.943739e-11, 8.738708e-11, 8.183308e-11, 8.398805e-11, 
    7.893401e-11, 7.584995e-11, 7.736314e-11, 6.839782e-11, 7.177849e-11, 
    5.538173e-11, 6.202359e-11, 4.594186e-11, 4.943319e-11, 4.513658e-11, 
    4.728822e-11, 4.365233e-11, 4.691351e-11, 4.138816e-11, 4.026124e-11, 
    4.102842e-11, 3.814876e-11, 4.710008e-11, 4.347164e-11, 7.740577e-11, 
    7.715723e-11, 7.600796e-11, 8.11634e-11, 8.148771e-11, 8.64687e-11, 
    8.202544e-11, 8.018895e-11, 7.567436e-11, 7.310048e-11, 7.071928e-11, 
    6.570251e-11, 6.044326e-11, 5.366967e-11, 4.920033e-11, 4.638146e-11, 
    4.809355e-11, 4.657931e-11, 4.827466e-11, 4.908694e-11, 4.068027e-11, 
    4.523617e-11, 3.85519e-11, 3.889832e-11, 4.183283e-11, 3.885916e-11, 
    7.698313e-11, 7.841947e-11, 8.357165e-11, 7.951755e-11, 8.702537e-11, 
    8.275648e-11, 8.03779e-11, 7.170597e-11, 6.990551e-11, 6.82679e-11, 
    6.512486e-11, 6.12634e-11, 5.494047e-11, 4.98854e-11, 4.561482e-11, 
    4.591697e-11, 4.581039e-11, 4.48961e-11, 4.718923e-11, 4.452877e-11, 
    4.409475e-11, 4.523693e-11, 3.894491e-11, 4.066108e-11, 3.890571e-11, 
    4.001497e-11, 7.795032e-11, 7.555719e-11, 7.684292e-11, 7.44393e-11, 
    7.612612e-11, 6.885254e-11, 6.678415e-11, 5.776278e-11, 6.133746e-11, 
    5.573031e-11, 6.074789e-11, 5.983278e-11, 5.55539e-11, 6.046778e-11, 
    5.015334e-11, 5.697137e-11, 4.486087e-11, 5.107204e-11, 4.449375e-11, 
    4.56326e-11, 4.37603e-11, 4.21389e-11, 4.017232e-11, 3.67498e-11, 
    3.751907e-11, 3.480581e-11, 7.209899e-11, 6.919398e-11, 6.944635e-11, 
    6.64994e-11, 6.438542e-11, 5.999051e-11, 5.345433e-11, 5.584002e-11, 
    5.152575e-11, 5.069366e-11, 5.727495e-11, 5.315554e-11, 6.730323e-11, 
    6.483033e-11, 6.629399e-11, 7.186608e-11, 5.528213e-11, 6.335249e-11, 
    4.912908e-11, 5.299738e-11, 4.236687e-11, 4.740431e-11, 3.794842e-11, 
    3.134702e-11, 2.901615e-11, 2.6454e-11, 6.764914e-11, 6.957732e-11, 
    6.615589e-11, 6.164669e-11, 5.769039e-11, 5.275436e-11, 5.22698e-11, 
    5.139165e-11, 4.917418e-11, 4.737185e-11, 5.111621e-11, 4.692884e-11, 
    6.426661e-11, 5.462351e-11, 7.03173e-11, 6.524972e-11, 6.190556e-11, 
    6.335543e-11, 5.611826e-11, 5.451498e-11, 4.838356e-11, 5.147761e-11, 
    3.527101e-11, 4.180262e-11, 2.461713e-11, 2.766242e-11, 7.026123e-11, 
    6.765591e-11, 5.918906e-11, 6.310335e-11, 5.243785e-11, 5.005412e-11, 
    4.818364e-11, 4.587753e-11, 4.563443e-11, 4.431834e-11, 4.649206e-11, 
    4.440267e-11, 5.274424e-11, 4.886818e-11, 6.011131e-11, 5.719645e-11, 
    5.852284e-11, 6.000624e-11, 5.552436e-11, 5.105532e-11, 5.096375e-11, 
    4.959743e-11, 4.590971e-11, 5.239788e-11, 3.139617e-11, 4.47944e-11, 
    6.490419e-11, 6.02643e-11, 5.962494e-11, 6.137389e-11, 5.028894e-11, 
    5.409694e-11, 4.435011e-11, 4.682658e-11, 4.282766e-11, 4.477709e-11, 
    4.507011e-11, 4.769769e-11, 4.939734e-11, 5.391717e-11, 5.784178e-11, 
    6.111775e-11, 6.034289e-11, 5.678964e-11, 5.079205e-11, 4.561223e-11, 
    4.67072e-11, 4.312107e-11, 5.315761e-11, 4.873442e-11, 5.040607e-11, 
    4.614457e-11, 5.590445e-11, 4.749472e-11, 5.824011e-11, 5.722462e-11, 
    5.417488e-11, 4.844549e-11, 4.724943e-11, 4.599882e-11, 4.67673e-11, 
    5.0647e-11, 5.130772e-11, 5.424753e-11, 5.508295e-11, 5.744451e-11, 
    5.946151e-11, 5.761627e-11, 5.572901e-11, 5.064555e-11, 4.63999e-11, 
    4.211612e-11, 4.112071e-11, 3.663992e-11, 4.025286e-11, 3.135753e-11, 
    3.933117e-11, 2.888559e-11, 4.704243e-11, 3.948447e-11, 5.403955e-11, 
    5.228327e-11, 4.922609e-11, 4.277577e-11, 4.616388e-11, 4.222317e-11, 
    5.133379e-11, 5.666986e-11, 5.812301e-11, 6.091425e-11, 5.806045e-11, 
    5.828842e-11, 5.565238e-11, 5.648863e-11, 5.04836e-11, 5.363998e-11, 
    4.507736e-11, 4.225326e-11, 3.508172e-11, 2.889654e-11, 2.6111e-11, 
    2.494547e-11, 2.459838e-11, 2.445431e-11,
  8.27314e-14, 7.055169e-14, 7.281933e-14, 6.371829e-14, 6.866776e-14, 
    6.285148e-14, 8.01578e-14, 7.009404e-14, 7.641503e-14, 8.158243e-14, 
    4.826444e-14, 6.3331e-14, 3.533273e-14, 4.296112e-14, 2.556761e-14, 
    3.645593e-14, 2.366757e-14, 2.584792e-14, 1.965447e-14, 2.131752e-14, 
    1.454472e-14, 1.891611e-14, 1.164471e-14, 1.552212e-14, 1.487132e-14, 
    1.907302e-14, 6.008155e-14, 4.999491e-14, 6.071765e-14, 5.919363e-14, 
    5.987454e-14, 6.856263e-14, 7.323985e-14, 8.371683e-14, 8.174537e-14, 
    7.408477e-14, 5.851666e-14, 6.353097e-14, 5.140706e-14, 5.166242e-14, 
    4.003661e-14, 4.50387e-14, 2.826855e-14, 3.252511e-14, 2.124637e-14, 
    2.379404e-14, 2.136179e-14, 2.208151e-14, 2.135252e-14, 2.516543e-14, 
    2.348211e-14, 2.702193e-14, 4.40723e-14, 3.849403e-14, 5.6643e-14, 
    6.98676e-14, 7.969724e-14, 8.720311e-14, 8.611451e-14, 8.406426e-14, 
    7.40414e-14, 6.53745e-14, 5.924075e-14, 5.53575e-14, 5.16992e-14, 
    4.159891e-14, 3.68221e-14, 2.745413e-14, 2.901466e-14, 2.64041e-14, 
    2.405779e-14, 2.042915e-14, 2.100026e-14, 1.949431e-14, 2.647134e-14, 
    2.168142e-14, 2.992859e-14, 2.750083e-14, 5.072963e-14, 6.215151e-14, 
    6.747551e-14, 7.237958e-14, 8.528364e-14, 7.622214e-14, 7.971331e-14, 
    7.157752e-14, 6.670548e-14, 6.908682e-14, 5.525375e-14, 6.038982e-14, 
    3.655082e-14, 4.5865e-14, 2.43242e-14, 2.868984e-14, 2.334633e-14, 
    2.598403e-14, 2.157453e-14, 2.551901e-14, 1.895233e-14, 1.768581e-14, 
    1.854515e-14, 1.538597e-14, 2.575026e-14, 2.136162e-14, 6.915416e-14, 
    6.876171e-14, 6.695331e-14, 7.514385e-14, 7.566564e-14, 8.37711e-14, 
    7.653245e-14, 7.358057e-14, 6.643033e-14, 6.242541e-14, 5.876967e-14, 
    5.123446e-14, 4.360253e-14, 3.423799e-14, 2.839257e-14, 2.486277e-14, 
    2.699129e-14, 2.510624e-14, 2.721927e-14, 2.824813e-14, 1.815364e-14, 
    2.346665e-14, 1.581709e-14, 1.619054e-14, 1.94593e-14, 1.614818e-14, 
    6.84871e-14, 7.075963e-14, 7.90362e-14, 7.250748e-14, 8.468728e-14, 
    7.771415e-14, 7.388315e-14, 6.027858e-14, 5.753168e-14, 5.505843e-14, 
    5.038223e-14, 4.477326e-14, 3.595104e-14, 2.92695e-14, 2.392569e-14, 
    2.42938e-14, 2.416378e-14, 2.305654e-14, 2.586096e-14, 2.261591e-14, 
    2.209843e-14, 2.346757e-14, 1.624097e-14, 1.813214e-14, 1.619853e-14, 
    1.741262e-14, 7.001563e-14, 6.624685e-14, 6.826612e-14, 6.450186e-14, 
    6.713876e-14, 5.593858e-14, 5.283905e-14, 3.982974e-14, 4.487934e-14, 
    3.70264e-14, 4.403649e-14, 4.273598e-14, 3.678552e-14, 4.363741e-14, 
    2.961443e-14, 3.873209e-14, 2.301419e-14, 3.080525e-14, 2.257402e-14, 
    2.394732e-14, 2.170205e-14, 1.981058e-14, 1.758702e-14, 1.391978e-14, 
    1.472019e-14, 1.196371e-14, 6.088196e-14, 5.645406e-14, 5.683574e-14, 
    5.241554e-14, 4.929618e-14, 4.295946e-14, 3.394985e-14, 3.71764e-14, 
    3.139792e-14, 3.031329e-14, 3.915223e-14, 3.355109e-14, 5.361311e-14, 
    4.994897e-14, 5.21105e-14, 6.052422e-14, 3.641522e-14, 4.77884e-14, 
    2.830179e-14, 3.334053e-14, 2.007343e-14, 2.612858e-14, 1.517312e-14, 
    1.157743e-14, 8.761244e-15, 6.081587e-15, 5.413036e-14, 5.703406e-14, 
    5.190565e-14, 4.532292e-14, 3.972902e-14, 3.301764e-14, 3.237628e-14, 
    3.122244e-14, 2.835925e-14, 2.608814e-14, 3.086281e-14, 2.5538e-14, 
    4.912218e-14, 3.552177e-14, 5.81574e-14, 5.056616e-14, 4.569508e-14, 
    4.779267e-14, 3.755752e-14, 3.537509e-14, 2.73566e-14, 3.133489e-14, 
    1.242281e-14, 1.942474e-14, 4.446713e-15, 7.289163e-15, 5.80721e-14, 
    5.414051e-14, 4.182684e-14, 4.742639e-14, 3.259833e-14, 2.948657e-14, 
    2.710464e-14, 2.424567e-14, 2.394955e-14, 2.236459e-14, 2.499879e-14, 
    2.24652e-14, 3.300421e-14, 2.797001e-14, 4.313082e-14, 3.904348e-14, 
    4.089099e-14, 4.298177e-14, 3.674522e-14, 3.078346e-14, 3.066424e-14, 
    2.890001e-14, 2.428493e-14, 3.254549e-14, 1.16405e-14, 2.293431e-14, 
    5.005755e-14, 4.334806e-14, 4.244192e-14, 4.493153e-14, 2.978941e-14, 
    3.481156e-14, 2.240247e-14, 2.541147e-14, 2.060785e-14, 2.291352e-14, 
    2.326613e-14, 2.649486e-14, 2.864402e-14, 3.456993e-14, 3.993971e-14, 
    4.456479e-14, 4.345977e-14, 3.848112e-14, 3.0441e-14, 2.392256e-14, 
    2.526398e-14, 2.09503e-14, 3.355386e-14, 2.780033e-14, 2.994077e-14, 
    2.457213e-14, 3.726457e-14, 2.62413e-14, 4.049542e-14, 3.90825e-14, 
    3.491645e-14, 2.743478e-14, 2.593579e-14, 2.43938e-14, 2.53382e-14, 
    3.025276e-14, 3.111274e-14, 3.501429e-14, 3.614442e-14, 3.93874e-14, 
    4.221105e-14, 3.962595e-14, 3.702463e-14, 3.025087e-14, 2.488544e-14, 
    1.978437e-14, 1.864935e-14, 1.380664e-14, 1.767649e-14, 1.15909e-14, 
    1.666097e-14, 8.61391e-15, 2.567874e-14, 1.682858e-14, 3.473437e-14, 
    3.239406e-14, 2.842541e-14, 2.054747e-14, 2.45958e-14, 1.990762e-14, 
    3.114681e-14, 3.831594e-14, 4.033186e-14, 4.427393e-14, 4.024454e-14, 
    4.056295e-14, 3.691994e-14, 3.806633e-14, 3.004107e-14, 3.419823e-14, 
    2.327487e-14, 1.994231e-14, 1.223531e-14, 8.626219e-15, 5.757653e-15, 
    4.720723e-15, 4.431308e-15, 4.313832e-15,
  2.796268e-19, 2.389788e-19, 2.465546e-19, 2.161257e-19, 2.32682e-19, 
    2.132241e-19, 2.710463e-19, 2.374494e-19, 2.585597e-19, 2.757966e-19, 
    1.642947e-19, 2.148294e-19, 1.20729e-19, 1.464527e-19, 8.76823e-20, 
    1.245213e-19, 8.123272e-20, 8.863317e-20, 6.758499e-20, 7.324514e-20, 
    5.014851e-20, 6.506983e-20, 4.025421e-20, 5.348965e-20, 5.12653e-20, 
    6.560445e-20, 2.039479e-19, 1.7011e-19, 2.060787e-19, 2.009729e-19, 
    2.032544e-19, 2.323305e-19, 2.479591e-19, 2.829111e-19, 2.763398e-19, 
    2.507807e-19, 1.987042e-19, 2.154987e-19, 1.748532e-19, 1.757108e-19, 
    1.365997e-19, 1.53446e-19, 9.683848e-20, 1.112424e-19, 7.30031e-20, 
    8.166224e-20, 7.339572e-20, 7.58432e-20, 7.336417e-20, 8.631771e-20, 
    8.06028e-20, 9.261411e-20, 1.501936e-19, 1.313983e-19, 1.924231e-19, 
    2.366926e-19, 2.695102e-19, 2.945256e-19, 2.908998e-19, 2.840689e-19, 
    2.506359e-19, 2.21668e-19, 2.011308e-19, 1.881119e-19, 1.758342e-19, 
    1.418645e-19, 1.257573e-19, 9.407902e-20, 9.93655e-20, 9.051945e-20, 
    8.255788e-20, 7.02224e-20, 7.216587e-20, 6.703952e-20, 9.074747e-20, 
    7.448281e-20, 1.024595e-19, 9.423729e-20, 1.725781e-19, 2.108806e-19, 
    2.286956e-19, 2.450858e-19, 2.881319e-19, 2.579159e-19, 2.695638e-19, 
    2.424064e-19, 2.261204e-19, 2.340829e-19, 1.877638e-19, 2.049805e-19, 
    1.248416e-19, 1.562261e-19, 8.346243e-20, 9.826548e-20, 8.014157e-20, 
    8.909485e-20, 7.411928e-20, 8.751741e-20, 6.519326e-20, 6.087579e-20, 
    6.380566e-20, 5.302441e-20, 8.830192e-20, 7.339513e-20, 2.34308e-19, 
    2.329961e-19, 2.269492e-19, 2.543166e-19, 2.560585e-19, 2.83092e-19, 
    2.589516e-19, 2.49097e-19, 2.252e-19, 2.117977e-19, 1.995522e-19, 
    1.742736e-19, 1.486122e-19, 1.17031e-19, 9.725862e-20, 8.529059e-20, 
    9.251027e-20, 8.611687e-20, 9.328304e-20, 9.67693e-20, 6.247106e-20, 
    8.055028e-20, 5.449741e-20, 5.577288e-20, 6.692031e-20, 5.562823e-20, 
    2.32078e-19, 2.396736e-19, 2.673054e-19, 2.45513e-19, 2.86145e-19, 
    2.628949e-19, 2.501074e-19, 2.046079e-19, 1.954027e-19, 1.871086e-19, 
    1.714111e-19, 1.525528e-19, 1.228168e-19, 1.002284e-19, 8.210934e-20, 
    8.335924e-20, 8.291778e-20, 7.915706e-20, 8.867741e-20, 7.765971e-20, 
    7.590071e-20, 8.055341e-20, 5.59451e-20, 6.239776e-20, 5.58002e-20, 
    5.994394e-20, 2.371873e-19, 2.245863e-19, 2.313392e-19, 2.187481e-19, 
    2.275694e-19, 1.900609e-19, 1.796611e-19, 1.359023e-19, 1.529098e-19, 
    1.264467e-19, 1.500731e-19, 1.456945e-19, 1.256338e-19, 1.487297e-19, 
    1.013961e-19, 1.322012e-19, 7.901314e-20, 1.054261e-19, 7.751737e-20, 
    8.218277e-20, 7.455295e-20, 6.811659e-20, 6.053887e-20, 4.80106e-20, 
    5.074858e-20, 4.130997e-20, 2.06629e-19, 1.917896e-19, 1.930694e-19, 
    1.782394e-19, 1.677623e-19, 1.464471e-19, 1.160574e-19, 1.26953e-19, 
    1.07431e-19, 1.037615e-19, 1.336181e-19, 1.147099e-19, 1.822591e-19, 
    1.699556e-19, 1.772153e-19, 2.054308e-19, 1.243839e-19, 1.626944e-19, 
    9.695109e-20, 1.139984e-19, 6.901154e-20, 8.958512e-20, 5.2297e-20, 
    4.002319e-20, 3.033592e-20, 2.10797e-20, 1.839949e-19, 1.937343e-19, 
    1.765275e-19, 1.544024e-19, 1.355628e-19, 1.129072e-19, 1.107393e-19, 
    1.068374e-19, 9.714572e-20, 8.944796e-20, 1.056209e-19, 8.758183e-20, 
    1.671776e-19, 1.213674e-19, 1.975002e-19, 1.72029e-19, 1.556545e-19, 
    1.627088e-19, 1.28239e-19, 1.20872e-19, 9.374848e-20, 1.072178e-19, 
    4.288393e-20, 6.680258e-20, 1.540766e-20, 2.525624e-20, 1.972142e-19, 
    1.840289e-19, 1.426324e-19, 1.614773e-19, 1.114899e-19, 1.009633e-19, 
    9.289447e-20, 8.31958e-20, 8.219033e-20, 7.68055e-20, 8.575222e-20, 
    7.71475e-20, 1.128618e-19, 9.58271e-20, 1.470241e-19, 1.332514e-19, 
    1.394793e-19, 1.465222e-19, 1.254978e-19, 1.053524e-19, 1.04949e-19, 
    9.897724e-20, 8.332912e-20, 1.113113e-19, 4.023975e-20, 7.874172e-20, 
    1.703204e-19, 1.477555e-19, 1.447042e-19, 1.530854e-19, 1.019885e-19, 
    1.189687e-19, 7.693427e-20, 8.715256e-20, 7.08306e-20, 7.867108e-20, 
    7.986912e-20, 9.082718e-20, 9.811028e-20, 1.181525e-19, 1.362731e-19, 
    1.518512e-19, 1.481316e-19, 1.313548e-19, 1.041937e-19, 8.209868e-20, 
    8.665213e-20, 7.199587e-20, 1.147193e-19, 9.525219e-20, 1.025008e-19, 
    8.430412e-20, 1.272505e-19, 8.996738e-20, 1.381462e-19, 1.333829e-19, 
    1.19323e-19, 9.401344e-20, 8.893123e-20, 8.369872e-20, 8.690394e-20, 
    1.035567e-19, 1.064663e-19, 1.196535e-19, 1.234697e-19, 1.34411e-19, 
    1.439266e-19, 1.352153e-19, 1.264408e-19, 1.035503e-19, 8.536755e-20, 
    6.802735e-20, 6.416081e-20, 4.762339e-20, 6.084401e-20, 4.006946e-20, 
    5.737902e-20, 2.982806e-20, 8.805928e-20, 5.795112e-20, 1.18708e-19, 
    1.107994e-19, 9.736985e-20, 7.06251e-20, 8.438443e-20, 6.844702e-20, 
    1.065816e-19, 1.307976e-19, 1.375949e-19, 1.508723e-19, 1.373006e-19, 
    1.383737e-19, 1.260875e-19, 1.299556e-19, 1.028402e-19, 1.168967e-19, 
    7.989882e-20, 6.856511e-20, 4.22412e-20, 2.987049e-20, 1.995759e-20, 
    1.635994e-20, 1.535411e-20, 1.494559e-20,
  2.052501e-25, 1.7556e-25, 1.810952e-25, 1.588576e-25, 1.709587e-25, 
    1.567364e-25, 1.989845e-25, 1.744425e-25, 1.898649e-25, 2.024533e-25, 
    1.209434e-25, 1.5791e-25, 8.902828e-26, 1.078789e-25, 6.47751e-26, 
    9.180861e-26, 6.003617e-26, 6.547359e-26, 5.000089e-26, 5.416417e-26, 
    3.716151e-26, 4.815025e-26, 2.987375e-26, 3.962365e-26, 3.79846e-26, 
    4.854365e-26, 1.49954e-25, 1.251999e-25, 1.515121e-25, 1.477785e-25, 
    1.494469e-25, 1.707018e-25, 1.821213e-25, 2.076482e-25, 2.0285e-25, 
    1.841825e-25, 1.461194e-25, 1.583993e-25, 1.286712e-25, 1.292987e-25, 
    1.006608e-25, 1.130006e-25, 7.149941e-26, 8.207072e-26, 5.398618e-26, 
    6.035183e-26, 5.42749e-26, 5.60745e-26, 5.42517e-26, 6.377262e-26, 
    5.957322e-26, 6.839749e-26, 1.106188e-25, 9.684927e-26, 1.415255e-25, 
    1.738895e-25, 1.978627e-25, 2.161276e-25, 2.134806e-25, 2.084935e-25, 
    1.840767e-25, 1.62909e-25, 1.47894e-25, 1.383719e-25, 1.293891e-25, 
    1.045181e-25, 9.271465e-26, 6.947325e-26, 7.335462e-26, 6.685911e-26, 
    6.101003e-26, 5.194106e-26, 5.337046e-26, 4.959958e-26, 6.702658e-26, 
    5.507426e-26, 7.562577e-26, 6.958947e-26, 1.270062e-25, 1.550231e-25, 
    1.680454e-25, 1.800221e-25, 2.114599e-25, 1.893947e-25, 1.979019e-25, 
    1.780644e-25, 1.661633e-25, 1.719824e-25, 1.381173e-25, 1.507091e-25, 
    9.204342e-26, 1.150363e-25, 6.167472e-26, 7.254708e-26, 5.923423e-26, 
    6.581273e-26, 5.480696e-26, 6.465398e-26, 4.824107e-26, 4.50633e-26, 
    4.72199e-26, 3.928087e-26, 6.523027e-26, 5.427446e-26, 1.721469e-25, 
    1.711882e-25, 1.667691e-25, 1.867656e-25, 1.880379e-25, 2.077803e-25, 
    1.901512e-25, 1.829525e-25, 1.654906e-25, 1.556936e-25, 1.467396e-25, 
    1.28247e-25, 1.094606e-25, 8.631669e-26, 7.180787e-26, 6.3018e-26, 
    6.832123e-26, 6.362507e-26, 6.888873e-26, 7.144862e-26, 4.623762e-26, 
    5.953462e-26, 4.036609e-26, 4.130564e-26, 4.951187e-26, 4.119909e-26, 
    1.705173e-25, 1.760677e-25, 1.962525e-25, 1.803342e-25, 2.100092e-25, 
    1.930313e-25, 1.836907e-25, 1.504366e-25, 1.437048e-25, 1.37638e-25, 
    1.261522e-25, 1.123465e-25, 9.055904e-26, 7.398803e-26, 6.068041e-26, 
    6.15989e-26, 6.12745e-26, 5.85106e-26, 6.55061e-26, 5.740994e-26, 
    5.611678e-26, 5.953692e-26, 4.143249e-26, 4.618366e-26, 4.132576e-26, 
    4.437726e-26, 1.74251e-25, 1.65042e-25, 1.699774e-25, 1.607746e-25, 
    1.672224e-25, 1.397976e-25, 1.321893e-25, 1.001498e-25, 1.126079e-25, 
    9.322006e-26, 1.105306e-25, 1.073236e-25, 9.262414e-26, 1.095467e-25, 
    7.484521e-26, 9.743769e-26, 5.840481e-26, 7.780298e-26, 5.73053e-26, 
    6.073437e-26, 5.512583e-26, 5.039199e-26, 4.481526e-26, 3.558551e-26, 
    3.760379e-26, 3.0643e-26, 1.519145e-25, 1.410621e-25, 1.419983e-25, 
    1.31149e-25, 1.234816e-25, 1.078748e-25, 8.56027e-26, 9.359113e-26, 
    7.927419e-26, 7.658133e-26, 9.8476e-26, 8.461443e-26, 1.340902e-25, 
    1.250869e-25, 1.303996e-25, 1.510383e-25, 9.170788e-26, 1.197719e-25, 
    7.15821e-26, 8.409251e-26, 5.105037e-26, 6.617285e-26, 3.874488e-26, 
    2.970317e-26, 2.254425e-26, 1.568876e-26, 1.353601e-25, 1.424846e-25, 
    1.298963e-25, 1.137009e-25, 9.990104e-26, 8.329203e-26, 8.170159e-26, 
    7.883865e-26, 7.172498e-26, 6.607209e-26, 7.79459e-26, 6.470129e-26, 
    1.230536e-25, 8.949636e-26, 1.452388e-25, 1.266043e-25, 1.146177e-25, 
    1.197824e-25, 9.453377e-26, 8.913318e-26, 6.923052e-26, 7.911776e-26, 
    3.180442e-26, 4.942524e-26, 1.147744e-26, 1.878435e-26, 1.450297e-25, 
    1.35385e-25, 1.050806e-25, 1.188809e-25, 8.225231e-26, 7.45275e-26, 
    6.860338e-26, 6.14788e-26, 6.073993e-26, 5.678198e-26, 6.335717e-26, 
    5.70334e-26, 8.325873e-26, 7.075683e-26, 1.082974e-25, 9.820727e-26, 
    1.027706e-25, 1.079298e-25, 9.252444e-26, 7.774889e-26, 7.745285e-26, 
    7.30696e-26, 6.157677e-26, 8.212125e-26, 2.986307e-26, 5.820531e-26, 
    1.253539e-25, 1.088332e-25, 1.065982e-25, 1.127365e-25, 7.527999e-26, 
    8.77376e-26, 5.687664e-26, 6.438595e-26, 5.238842e-26, 5.815339e-26, 
    5.903399e-26, 6.708513e-26, 7.243314e-26, 8.713907e-26, 1.004215e-25, 
    1.118327e-25, 1.091086e-25, 9.681737e-26, 7.68985e-26, 6.067257e-26, 
    6.401831e-26, 5.324544e-26, 8.462131e-26, 7.03347e-26, 7.565601e-26, 
    6.229319e-26, 9.380922e-26, 6.645362e-26, 1.017939e-25, 9.830369e-26, 
    8.799739e-26, 6.942509e-26, 6.569255e-26, 6.184836e-26, 6.42033e-26, 
    7.643101e-26, 7.856634e-26, 8.823971e-26, 9.103769e-26, 9.905707e-26, 
    1.060286e-25, 9.964643e-26, 9.321569e-26, 7.642631e-26, 6.307454e-26, 
    5.032634e-26, 4.748128e-26, 3.530002e-26, 4.503991e-26, 2.973734e-26, 
    4.248858e-26, 2.216855e-26, 6.505203e-26, 4.290989e-26, 8.754642e-26, 
    8.174567e-26, 7.188954e-26, 5.223727e-26, 6.23522e-26, 5.063508e-26, 
    7.865091e-26, 9.640903e-26, 1.0139e-25, 1.111158e-25, 1.011744e-25, 
    1.019607e-25, 9.295671e-26, 9.579195e-26, 7.590518e-26, 8.62182e-26, 
    5.905581e-26, 5.072196e-26, 3.133019e-26, 2.219994e-26, 1.485636e-26, 
    1.218517e-26, 1.143763e-26, 1.113392e-26,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_SAT =
  0.0104524, 0.01046719, 0.01046431, 0.01047624, 0.01046961, 0.01047743, 
    0.01045539, 0.01046779, 0.01045987, 0.01045371, 0.01049936, 0.01047676, 
    0.01052261, 0.01050829, 0.01054417, 0.0105204, 0.01054895, 0.01054346, 
    0.0105599, 0.01055519, 0.01057623, 0.01056207, 0.01058706, 0.01057284, 
    0.01057508, 0.0105616, 0.01048129, 0.01049656, 0.01048039, 0.01048257, 
    0.01048158, 0.01046976, 0.01046381, 0.01045125, 0.01045352, 0.01046274, 
    0.01048355, 0.01047647, 0.01049423, 0.01049383, 0.01051356, 0.01050467, 
    0.01053772, 0.01052834, 0.01055539, 0.0105486, 0.01055507, 0.01055311, 
    0.0105551, 0.01054514, 0.01054941, 0.01054063, 0.01050634, 0.01051645, 
    0.01048627, 0.01046811, 0.01045594, 0.01044731, 0.01044853, 0.01045086, 
    0.0104628, 0.01047397, 0.01048248, 0.01048817, 0.01049377, 0.01051077, 
    0.01051967, 0.01053963, 0.01053601, 0.01054212, 0.01054792, 0.01055768, 
    0.01055607, 0.01056037, 0.01054194, 0.01055421, 0.01053395, 0.0105395, 
    0.0104954, 0.01047838, 0.01047122, 0.01046487, 0.01044947, 0.01046011, 
    0.01045592, 0.01046587, 0.01047219, 0.01046906, 0.01048833, 0.01048085, 
    0.0105202, 0.01050328, 0.01054725, 0.01053675, 0.01054976, 0.01054312, 
    0.0105545, 0.01054426, 0.01056197, 0.01056583, 0.01056319, 0.01057328, 
    0.01054369, 0.01055508, 0.01046898, 0.01046949, 0.01047186, 0.01046143, 
    0.01046079, 0.01045119, 0.01045972, 0.01046336, 0.01047255, 0.010478, 
    0.01048316, 0.01049451, 0.01050717, 0.01052481, 0.01053743, 0.01054588, 
    0.01054069, 0.01054528, 0.01054016, 0.01053775, 0.01056439, 0.01054946, 
    0.01057183, 0.01057059, 0.01056048, 0.01057073, 0.01046984, 0.0104669, 
    0.01045672, 0.01046469, 0.01045014, 0.0104583, 0.010463, 0.01048103, 
    0.01048495, 0.01048863, 0.01049585, 0.01050513, 0.01052137, 0.01053545, 
    0.01054825, 0.01054731, 0.01054765, 0.01055052, 0.01054342, 0.01055168, 
    0.01055307, 0.01054944, 0.01057042, 0.01056444, 0.01057056, 0.01056666, 
    0.01046786, 0.0104728, 0.01047013, 0.01047515, 0.01047162, 0.01048733, 
    0.01049204, 0.01051397, 0.01050495, 0.01051926, 0.0105064, 0.01050868, 
    0.01051977, 0.01050709, 0.01053469, 0.01051603, 0.01055063, 0.01053208, 
    0.01055179, 0.0105482, 0.01055413, 0.01055945, 0.01056612, 0.01057844, 
    0.01057558, 0.01058585, 0.01048015, 0.01048656, 0.01048597, 0.01049266, 
    0.0104976, 0.01050828, 0.01052538, 0.01051895, 0.01053074, 0.01053311, 
    0.01051519, 0.01052621, 0.01049083, 0.01049658, 0.01049314, 0.01048067, 
    0.01052046, 0.01050008, 0.01053764, 0.01052664, 0.0105587, 0.01054279, 
    0.01057401, 0.01058736, 0.01059981, 0.01061443, 0.01049003, 0.01048568, 
    0.01049345, 0.01050421, 0.01051413, 0.01052731, 0.01052865, 0.01053112, 
    0.0105375, 0.01054286, 0.01053192, 0.01054421, 0.01049795, 0.01052222, 
    0.01048405, 0.0104956, 0.01050357, 0.01050005, 0.01051821, 0.01052249, 
    0.01053985, 0.01053087, 0.01058409, 0.0105606, 0.01062547, 0.01060742, 
    0.01048417, 0.01049, 0.01051031, 0.01050065, 0.01052818, 0.01053495, 
    0.01054043, 0.01054745, 0.0105482, 0.01055235, 0.01054554, 0.01055208, 
    0.01052734, 0.0105384, 0.01050797, 0.0105154, 0.01051198, 0.01050823, 
    0.01051978, 0.0105321, 0.01053233, 0.01053628, 0.01054745, 0.01052829, 
    0.01058717, 0.01055093, 0.01049637, 0.01050763, 0.0105092, 0.01050485, 
    0.01053427, 0.01052363, 0.01055225, 0.01054452, 0.01055717, 0.01055089, 
    0.01054997, 0.01054188, 0.01053685, 0.01052412, 0.01051374, 0.01050547, 
    0.01050739, 0.01051647, 0.01053285, 0.01054828, 0.01054491, 0.01055621, 
    0.01052619, 0.01053881, 0.01053395, 0.01054662, 0.01051879, 0.01054259, 
    0.0105127, 0.01051532, 0.01052342, 0.01053969, 0.01054324, 0.01054708, 
    0.0105447, 0.01053326, 0.01053136, 0.01052321, 0.01052098, 0.01051475, 
    0.0105096, 0.01051431, 0.01051926, 0.01053325, 0.01054584, 0.01055953, 
    0.01056287, 0.0105789, 0.0105659, 0.01058738, 0.01056918, 0.01060061, 
    0.01054392, 0.01056858, 0.01052377, 0.01052861, 0.01053738, 0.01055738, 
    0.01054656, 0.0105592, 0.01053129, 0.0105168, 0.010513, 0.01050598, 
    0.01051316, 0.01051258, 0.01051944, 0.01051724, 0.01053371, 0.01052487, 
    0.01054995, 0.01055909, 0.01058479, 0.0106005, 0.01061641, 0.01062343, 
    0.01062557, 0.01062646,
  3.328509e-05, 3.337547e-05, 3.335786e-05, 3.343088e-05, 3.339029e-05, 
    3.343821e-05, 3.330334e-05, 3.337913e-05, 3.333071e-05, 3.329312e-05, 
    3.357355e-05, 3.343413e-05, 3.371737e-05, 3.362875e-05, 3.385097e-05, 
    3.370369e-05, 3.388059e-05, 3.384654e-05, 3.394856e-05, 3.391933e-05, 
    3.405006e-05, 3.396203e-05, 3.411745e-05, 3.402895e-05, 3.404287e-05, 
    3.395916e-05, 3.346203e-05, 3.355626e-05, 3.345648e-05, 3.346992e-05, 
    3.346385e-05, 3.339118e-05, 3.335482e-05, 3.327806e-05, 3.329197e-05, 
    3.334827e-05, 3.347595e-05, 3.343233e-05, 3.354188e-05, 3.353941e-05, 
    3.366135e-05, 3.360639e-05, 3.381096e-05, 3.375282e-05, 3.392055e-05, 
    3.387843e-05, 3.39186e-05, 3.39064e-05, 3.391876e-05, 3.385697e-05, 
    3.388346e-05, 3.3829e-05, 3.361672e-05, 3.367922e-05, 3.349279e-05, 
    3.338107e-05, 3.33067e-05, 3.325403e-05, 3.326147e-05, 3.327571e-05, 
    3.334861e-05, 3.341694e-05, 3.346938e-05, 3.350449e-05, 3.353905e-05, 
    3.364406e-05, 3.369919e-05, 3.38228e-05, 3.380035e-05, 3.383826e-05, 
    3.387423e-05, 3.39348e-05, 3.392481e-05, 3.395152e-05, 3.383714e-05, 
    3.391323e-05, 3.378759e-05, 3.3822e-05, 3.354907e-05, 3.344407e-05, 
    3.34001e-05, 3.336127e-05, 3.326721e-05, 3.333221e-05, 3.330661e-05, 
    3.336738e-05, 3.340606e-05, 3.338691e-05, 3.350545e-05, 3.345931e-05, 
    3.370246e-05, 3.35978e-05, 3.387003e-05, 3.380494e-05, 3.38856e-05, 
    3.384442e-05, 3.391502e-05, 3.385148e-05, 3.396141e-05, 3.39854e-05, 
    3.396902e-05, 3.403171e-05, 3.384798e-05, 3.391866e-05, 3.33864e-05, 
    3.338953e-05, 3.340403e-05, 3.334028e-05, 3.333635e-05, 3.327771e-05, 
    3.332983e-05, 3.335207e-05, 3.340826e-05, 3.344173e-05, 3.34736e-05, 
    3.354362e-05, 3.362186e-05, 3.373097e-05, 3.380917e-05, 3.386158e-05, 
    3.38294e-05, 3.385782e-05, 3.382608e-05, 3.381117e-05, 3.397645e-05, 
    3.388374e-05, 3.402269e-05, 3.401499e-05, 3.395218e-05, 3.401585e-05, 
    3.339172e-05, 3.337373e-05, 3.331147e-05, 3.33602e-05, 3.327131e-05, 
    3.332115e-05, 3.334984e-05, 3.34604e-05, 3.348465e-05, 3.350731e-05, 
    3.355192e-05, 3.360921e-05, 3.370965e-05, 3.379686e-05, 3.387629e-05, 
    3.387047e-05, 3.387252e-05, 3.389032e-05, 3.384631e-05, 3.389754e-05, 
    3.390619e-05, 3.388366e-05, 3.401396e-05, 3.397675e-05, 3.401483e-05, 
    3.399058e-05, 3.337956e-05, 3.340979e-05, 3.339347e-05, 3.342421e-05, 
    3.340259e-05, 3.349932e-05, 3.352834e-05, 3.366386e-05, 3.360811e-05, 
    3.369665e-05, 3.361706e-05, 3.363121e-05, 3.369979e-05, 3.362133e-05, 
    3.379217e-05, 3.367661e-05, 3.389101e-05, 3.3776e-05, 3.389823e-05, 
    3.387595e-05, 3.391277e-05, 3.39458e-05, 3.398722e-05, 3.406376e-05, 
    3.404602e-05, 3.410989e-05, 3.345501e-05, 3.349453e-05, 3.349093e-05, 
    3.353219e-05, 3.356271e-05, 3.362869e-05, 3.373454e-05, 3.369472e-05, 
    3.376769e-05, 3.378238e-05, 3.367143e-05, 3.373968e-05, 3.352088e-05, 
    3.355639e-05, 3.353516e-05, 3.34582e-05, 3.370406e-05, 3.357804e-05, 
    3.381049e-05, 3.37423e-05, 3.394111e-05, 3.384242e-05, 3.403627e-05, 
    3.411931e-05, 3.419682e-05, 3.428794e-05, 3.351596e-05, 3.348913e-05, 
    3.353706e-05, 3.360354e-05, 3.366486e-05, 3.374648e-05, 3.375476e-05, 
    3.377008e-05, 3.38096e-05, 3.384287e-05, 3.377504e-05, 3.385119e-05, 
    3.356485e-05, 3.371494e-05, 3.347909e-05, 3.355033e-05, 3.359958e-05, 
    3.357786e-05, 3.369014e-05, 3.371662e-05, 3.382419e-05, 3.376853e-05, 
    3.409892e-05, 3.395294e-05, 3.435685e-05, 3.424428e-05, 3.347978e-05, 
    3.351581e-05, 3.364126e-05, 3.358158e-05, 3.375186e-05, 3.379378e-05, 
    3.382774e-05, 3.387132e-05, 3.387593e-05, 3.390173e-05, 3.385947e-05, 
    3.390001e-05, 3.374666e-05, 3.381521e-05, 3.362679e-05, 3.367276e-05, 
    3.365158e-05, 3.362842e-05, 3.369988e-05, 3.377613e-05, 3.377757e-05, 
    3.380204e-05, 3.387129e-05, 3.375255e-05, 3.41181e-05, 3.389287e-05, 
    3.355509e-05, 3.362468e-05, 3.363439e-05, 3.360748e-05, 3.378959e-05, 
    3.372367e-05, 3.390107e-05, 3.385312e-05, 3.393162e-05, 3.389264e-05, 
    3.388691e-05, 3.383678e-05, 3.380559e-05, 3.372673e-05, 3.366246e-05, 
    3.361136e-05, 3.362323e-05, 3.367935e-05, 3.378075e-05, 3.387644e-05, 
    3.385551e-05, 3.392565e-05, 3.373954e-05, 3.381773e-05, 3.378758e-05, 
    3.386614e-05, 3.36937e-05, 3.384113e-05, 3.365604e-05, 3.367224e-05, 
    3.372236e-05, 3.382316e-05, 3.384516e-05, 3.386899e-05, 3.385424e-05, 
    3.378329e-05, 3.377158e-05, 3.37211e-05, 3.370725e-05, 3.36687e-05, 
    3.363687e-05, 3.3666e-05, 3.369663e-05, 3.378324e-05, 3.386132e-05, 
    3.39463e-05, 3.3967e-05, 3.406662e-05, 3.39858e-05, 3.411938e-05, 
    3.400621e-05, 3.420181e-05, 3.384939e-05, 3.400251e-05, 3.372458e-05, 
    3.375452e-05, 3.380885e-05, 3.393292e-05, 3.386577e-05, 3.394421e-05, 
    3.37711e-05, 3.368138e-05, 3.365791e-05, 3.36145e-05, 3.36589e-05, 
    3.365528e-05, 3.369776e-05, 3.36841e-05, 3.378611e-05, 3.373132e-05, 
    3.388682e-05, 3.394354e-05, 3.410326e-05, 3.420113e-05, 3.430032e-05, 
    3.434416e-05, 3.435749e-05, 3.436307e-05,
  7.912032e-10, 7.938588e-10, 7.933413e-10, 7.954884e-10, 7.942945e-10, 
    7.957045e-10, 7.917394e-10, 7.939662e-10, 7.925434e-10, 7.914393e-10, 
    7.996949e-10, 7.955843e-10, 8.039432e-10, 8.013252e-10, 8.079161e-10, 
    8.035388e-10, 8.0882e-10, 8.077813e-10, 8.108947e-10, 8.100025e-10, 
    8.139955e-10, 8.113065e-10, 8.160567e-10, 8.133505e-10, 8.137759e-10, 
    8.112186e-10, 7.964067e-10, 7.991848e-10, 7.962432e-10, 7.966391e-10, 
    7.964604e-10, 7.943208e-10, 7.932515e-10, 7.909969e-10, 7.914053e-10, 
    7.930593e-10, 7.96817e-10, 7.955314e-10, 7.987616e-10, 7.986885e-10, 
    8.02288e-10, 8.006652e-10, 8.06711e-10, 8.049916e-10, 8.100396e-10, 
    8.087541e-10, 8.099801e-10, 8.096077e-10, 8.09985e-10, 8.080994e-10, 
    8.089076e-10, 8.072466e-10, 8.009701e-10, 8.02816e-10, 7.973133e-10, 
    7.940231e-10, 7.91838e-10, 7.902912e-10, 7.905099e-10, 7.909278e-10, 
    7.930691e-10, 7.950783e-10, 7.966234e-10, 7.976587e-10, 7.986781e-10, 
    8.017769e-10, 8.034057e-10, 8.070611e-10, 8.063971e-10, 8.075285e-10, 
    8.08626e-10, 8.104746e-10, 8.101697e-10, 8.109852e-10, 8.074948e-10, 
    8.098162e-10, 8.060199e-10, 8.070377e-10, 7.989725e-10, 7.958774e-10, 
    7.945826e-10, 7.934414e-10, 7.906784e-10, 7.925874e-10, 7.918352e-10, 
    7.936212e-10, 7.947584e-10, 7.941952e-10, 7.97687e-10, 7.963264e-10, 
    8.035024e-10, 8.004113e-10, 8.08498e-10, 8.06533e-10, 8.089732e-10, 
    8.077169e-10, 8.098707e-10, 8.079323e-10, 8.112873e-10, 8.120198e-10, 
    8.115196e-10, 8.13435e-10, 8.078253e-10, 8.099819e-10, 7.941802e-10, 
    7.942722e-10, 7.946987e-10, 7.928245e-10, 7.92709e-10, 7.909865e-10, 
    7.925176e-10, 7.93171e-10, 7.94823e-10, 7.958085e-10, 7.967478e-10, 
    7.988127e-10, 8.011217e-10, 8.043452e-10, 8.066581e-10, 8.082403e-10, 
    8.07259e-10, 8.081254e-10, 8.071585e-10, 8.067175e-10, 8.117465e-10, 
    8.089161e-10, 8.131595e-10, 8.129241e-10, 8.110052e-10, 8.129507e-10, 
    7.943365e-10, 7.938079e-10, 7.919781e-10, 7.934101e-10, 7.907987e-10, 
    7.922625e-10, 7.931054e-10, 7.963587e-10, 7.970735e-10, 7.977418e-10, 
    7.990577e-10, 8.007484e-10, 8.037153e-10, 8.062938e-10, 8.086891e-10, 
    8.085113e-10, 8.08574e-10, 8.091171e-10, 8.077744e-10, 8.093374e-10, 
    8.096013e-10, 8.089137e-10, 8.128927e-10, 8.117558e-10, 8.129192e-10, 
    8.121784e-10, 7.939793e-10, 7.948679e-10, 7.94388e-10, 7.95292e-10, 
    7.946563e-10, 7.975059e-10, 7.983618e-10, 8.023621e-10, 8.00716e-10, 
    8.033309e-10, 8.009803e-10, 8.013978e-10, 8.034235e-10, 8.011062e-10, 
    8.061549e-10, 8.027387e-10, 8.091382e-10, 8.056765e-10, 8.093584e-10, 
    8.086787e-10, 8.098023e-10, 8.108105e-10, 8.120755e-10, 8.144148e-10, 
    8.138724e-10, 8.158257e-10, 7.961999e-10, 7.973647e-10, 7.972589e-10, 
    7.984756e-10, 7.993761e-10, 8.013237e-10, 8.044511e-10, 8.03274e-10, 
    8.054313e-10, 8.058655e-10, 8.025861e-10, 8.046028e-10, 7.981417e-10, 
    7.99189e-10, 7.985631e-10, 7.962937e-10, 8.035498e-10, 7.99828e-10, 
    8.06697e-10, 8.046803e-10, 8.106672e-10, 8.076554e-10, 8.135746e-10, 
    8.161133e-10, 8.184868e-10, 8.212782e-10, 7.979968e-10, 7.972057e-10, 
    7.986193e-10, 8.005809e-10, 8.023917e-10, 8.04804e-10, 8.05049e-10, 
    8.055019e-10, 8.066708e-10, 8.076694e-10, 8.056482e-10, 8.079233e-10, 
    7.994384e-10, 8.038713e-10, 7.969096e-10, 7.990105e-10, 8.004639e-10, 
    7.99823e-10, 8.031387e-10, 8.039213e-10, 8.071023e-10, 8.05456e-10, 
    8.154897e-10, 8.110281e-10, 8.233921e-10, 8.199399e-10, 7.969302e-10, 
    7.979926e-10, 8.016948e-10, 7.999328e-10, 8.049633e-10, 8.062028e-10, 
    8.072082e-10, 8.085371e-10, 8.086781e-10, 8.094651e-10, 8.081759e-10, 
    8.094129e-10, 8.048091e-10, 8.068367e-10, 8.012677e-10, 8.026252e-10, 
    8.019996e-10, 8.013158e-10, 8.034266e-10, 8.056806e-10, 8.057235e-10, 
    8.064471e-10, 8.08535e-10, 8.049835e-10, 8.160754e-10, 8.091936e-10, 
    7.991514e-10, 8.012049e-10, 8.014918e-10, 8.006975e-10, 8.060788e-10, 
    8.041297e-10, 8.094451e-10, 8.079823e-10, 8.103777e-10, 8.091879e-10, 
    8.090131e-10, 8.074837e-10, 8.065523e-10, 8.042201e-10, 8.023208e-10, 
    8.00812e-10, 8.011625e-10, 8.028197e-10, 8.058172e-10, 8.086933e-10, 
    8.080549e-10, 8.101956e-10, 8.045987e-10, 8.069112e-10, 8.060191e-10, 
    8.083793e-10, 8.032439e-10, 8.076154e-10, 8.021314e-10, 8.026101e-10, 
    8.04091e-10, 8.070716e-10, 8.077394e-10, 8.08466e-10, 8.080165e-10, 
    8.058924e-10, 8.05546e-10, 8.040537e-10, 8.036443e-10, 8.025055e-10, 
    8.015651e-10, 8.024256e-10, 8.033303e-10, 8.058911e-10, 8.082322e-10, 
    8.108257e-10, 8.114582e-10, 8.145015e-10, 8.120315e-10, 8.161148e-10, 
    8.126543e-10, 8.186385e-10, 8.078677e-10, 8.125419e-10, 8.041566e-10, 
    8.050418e-10, 8.066484e-10, 8.104169e-10, 8.083679e-10, 8.107616e-10, 
    8.05532e-10, 8.028795e-10, 8.021867e-10, 8.009047e-10, 8.02216e-10, 
    8.021091e-10, 8.033641e-10, 8.029605e-10, 8.05976e-10, 8.04356e-10, 
    8.090101e-10, 8.107413e-10, 8.156229e-10, 8.186183e-10, 8.216583e-10, 
    8.23003e-10, 8.234118e-10, 8.23583e-10,
  4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13,
  4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13,
  3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13,
  3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13,
  3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_UNSAT =
  0.8203498, 0.8517787, 0.8456301, 0.8712655, 0.8570073, 0.8738492, 
    0.8266826, 0.8530346, 0.8361722, 0.8231615, 0.9218926, 0.8724172, 
    0.9737335, 0.9414821, 1.023219, 0.9686847, 1.034327, 1.021639, 1.059969, 
    1.048951, 1.098321, 1.065063, 1.124078, 1.090365, 1.095626, 1.063969, 
    0.8822922, 0.9156732, 0.8803285, 0.8850547, 0.8829342, 0.8572988, 
    0.8444967, 0.817973, 0.8227617, 0.8422583, 0.8871834, 0.8718283, 
    0.9107433, 0.9098573, 0.9533231, 0.9334239, 1.008381, 0.9868718, 
    1.049411, 1.033578, 1.048665, 1.044085, 1.048724, 1.02553, 1.03545, 
    1.015107, 0.9371371, 0.9598185, 0.8931782, 0.8536512, 0.8278298, 
    0.8097132, 0.8122635, 0.8171341, 0.8423728, 0.8664089, 0.8849137, 
    0.8973793, 0.9097298, 0.9469056, 0.9670687, 1.012745, 1.004456, 1.018515, 
    1.032006, 1.054759, 1.051006, 1.061059, 1.018147, 1.046613, 0.999743, 
    1.012499, 0.9130783, 0.8759609, 0.8603567, 0.8468098, 0.8142264, 
    0.8366672, 0.8277883, 0.8489832, 0.8625671, 0.8558381, 0.8977212, 
    0.8813403, 0.9682688, 0.9302878, 1.03043, 1.006156, 1.036274, 1.020874, 
    1.047297, 1.023508, 1.064808, 1.07385, 1.067669, 1.09146, 1.022193, 
    1.048662, 0.8556489, 0.8567446, 0.8618595, 0.8394723, 0.8381121, 
    0.8178409, 0.8358694, 0.8435971, 0.8633589, 0.8751345, 0.8863906, 
    0.911341, 0.93896, 0.9787657, 1.007724, 1.027283, 1.015278, 1.025875, 
    1.01403, 1.008494, 1.070459, 1.035541, 1.088032, 1.085114, 1.061298, 
    1.085443, 0.8575147, 0.8512145, 0.8294891, 0.8464706, 0.8156468, 
    0.8328364, 0.8427898, 0.8816771, 0.8903226, 0.8983632, 0.9143312, 
    0.9344383, 0.9709489, 1.003127, 1.032794, 1.030612, 1.03138, 1.038036, 
    1.021567, 1.040747, 1.043974, 1.03554, 1.084723, 1.07062, 1.085052, 
    1.075865, 0.8532608, 0.8638847, 0.8581367, 0.8689577, 0.8613268, 
    0.8954638, 0.9058021, 0.9541758, 0.9340304, 0.9661743, 0.9372782, 
    0.9423727, 0.9672208, 0.9388324, 1.001339, 0.9587939, 1.038295, 
    0.9952925, 1.041007, 1.032665, 1.046488, 1.058906, 1.074579, 1.103612, 
    1.096878, 1.121231, 0.8798263, 0.8937894, 0.8925602, 0.9072606, 
    0.9181913, 0.9414929, 0.9801116, 0.9655237, 0.9923674, 0.997785, 
    0.9570304, 0.9819793, 0.9031858, 0.915854, 0.9083061, 0.8809223, 
    0.968873, 0.9236501, 1.008204, 0.9829778, 1.057132, 1.020052, 1.093173, 
    1.124719, 1.154513, 1.189335, 0.9014509, 0.8919209, 0.9090161, 0.9323339, 
    0.9546049, 0.9845097, 0.9875898, 0.9932329, 1.007904, 1.020288, 
    0.9950155, 1.0234, 0.9187939, 0.9728824, 0.8883247, 0.9136711, 0.9309284, 
    0.923642, 0.9638624, 0.9735541, 1.013276, 0.9926789, 1.116919, 1.061527, 
    1.215823, 1.172618, 0.8885996, 0.9014198, 0.9460009, 0.9249896, 
    0.9865197, 1.002007, 1.014657, 1.030891, 1.032651, 1.042308, 1.026495, 
    1.041684, 0.9845737, 1.009974, 0.9408191, 0.9574862, 0.9498062, 
    0.9414062, 0.9674211, 0.9954109, 0.9960182, 1.00505, 1.030625, 0.986774, 
    1.124087, 1.038753, 0.9154806, 0.9399521, 0.9435433, 0.9338354, 1.00045, 
    0.9761227, 1.042073, 1.024122, 1.053579, 1.038913, 1.03676, 1.018017, 
    1.006397, 0.9772325, 0.9537258, 0.9352417, 0.9395276, 0.959875, 
    0.9971332, 1.032807, 1.02496, 1.051333, 0.9819722, 1.01088, 0.9996724, 
    1.028975, 0.9651356, 1.019398, 0.9514303, 0.9573246, 0.975642, 1.012846, 
    1.021145, 1.030018, 1.024542, 0.9980865, 0.9937759, 0.9751968, 0.9700856, 
    0.9560406, 0.9444678, 0.9550378, 0.9661843, 0.9981003, 1.027146, 
    1.059082, 1.066936, 1.104567, 1.073906, 1.124564, 1.081456, 1.156203, 
    1.02258, 1.080206, 0.9764806, 0.9875047, 1.007542, 1.053964, 1.028836, 
    1.058241, 0.9936077, 0.9605769, 0.9521042, 0.9363602, 0.9524653, 
    0.9511518, 0.9666514, 0.9616609, 0.999166, 0.9789582, 1.036704, 1.058009, 
    1.118673, 1.156077, 1.194195, 1.210997, 1.216105, 1.21824,
  0.8834646, 0.8687027, 0.8715314, 0.8599308, 0.8663218, 0.8587898, 
    0.8804301, 0.8681275, 0.8759388, 0.8821148, 0.838492, 0.8594217, 
    0.7817581, 0.7896651, 0.7708438, 0.7829533, 0.7685931, 0.7711711, 
    0.7636739, 0.7657411, 0.7570257, 0.7627419, 0.753041, 0.7583355, 
    0.7574655, 0.7629408, 0.8550981, 0.8410197, 0.855952, 0.8539003, 
    0.8548194, 0.8661885, 0.8720528, 0.8846142, 0.8823066, 0.8730937, 
    0.8529818, 0.8596839, 0.8430533, 0.8434192, 0.786689, 0.7917405, 
    0.7739649, 0.7787198, 0.7656535, 0.7687438, 0.7657956, 0.7666767, 
    0.7657843, 0.7703706, 0.7683704, 0.7725347, 0.7907791, 0.7850924, 
    0.8504156, 0.8678431, 0.8798828, 0.8886358, 0.8873882, 0.8850189, 
    0.8730403, 0.8620917, 0.8539633, 0.8486344, 0.8434718, 0.7882886, 
    0.78334, 0.7730331, 0.7748123, 0.7718196, 0.7690585, 0.7646424, 
    0.7653501, 0.7634727, 0.7718972, 0.7661883, 0.7758419, 0.7730862, 
    0.8420826, 0.8578629, 0.8648024, 0.870986, 0.8864312, 0.8757052, 
    0.8799021, 0.8699866, 0.8638121, 0.8668534, 0.84849, 0.8555121, 
    0.7830533, 0.792558, 0.7693756, 0.7744442, 0.7682073, 0.7713298, 
    0.7660571, 0.7707858, 0.7627881, 0.7611691, 0.7622706, 0.7581537, 
    0.7710568, 0.7657957, 0.8669389, 0.8664411, 0.8641306, 0.8743919, 
    0.8750283, 0.8846776, 0.8760812, 0.8724725, 0.8634573, 0.8582259, 
    0.853325, 0.8428059, 0.7903096, 0.7805822, 0.7741062, 0.7700135, 
    0.7724991, 0.7703006, 0.7727622, 0.7739413, 0.7617705, 0.768352, 
    0.7587267, 0.75922, 0.7634288, 0.7591642, 0.866092, 0.8689629, 0.8790943, 
    0.8711442, 0.8857413, 0.8775089, 0.8728459, 0.8553636, 0.8516364, 
    0.848218, 0.8415775, 0.791477, 0.7824166, 0.7751007, 0.7689009, 
    0.7693393, 0.7691846, 0.7678587, 0.7711862, 0.7673262, 0.7666977, 
    0.7683529, 0.7592864, 0.7617425, 0.7592305, 0.7608157, 0.8680274, 
    0.8632209, 0.8658105, 0.8609558, 0.8643692, 0.8494426, 0.8450973, 
    0.7864767, 0.7915826, 0.783555, 0.7907431, 0.7894383, 0.7833022, 
    0.7903438, 0.77549, 0.785341, 0.7678076, 0.776823, 0.7672755, 0.7689267, 
    0.7662131, 0.76387, 0.7610413, 0.7561767, 0.7572617, 0.7534631, 
    0.8561717, 0.8501551, 0.8506806, 0.8444943, 0.8400005, 0.7896631, 
    0.7802706, 0.7837123, 0.7774789, 0.7762729, 0.7857754, 0.7798389, 
    0.8461913, 0.8409511, 0.8440599, 0.8556929, 0.7829095, 0.8377883, 
    0.7740029, 0.7796097, 0.764199, 0.7714992, 0.7578697, 0.7529458, 
    0.7488283, 0.7446707, 0.8469189, 0.8509534, 0.843767, 0.7920228, 
    0.786372, 0.7792583, 0.7785566, 0.7772848, 0.774068, 0.7714513, 
    0.7768861, 0.770808, 0.8397489, 0.7819595, 0.852492, 0.8418446, 
    0.7923903, 0.8377938, 0.7841127, 0.7818022, 0.7729208, 0.7774091, 
    0.7541092, 0.7633858, 0.7419911, 0.7465773, 0.8523752, 0.8469328, 
    0.7885188, 0.8372519, 0.7787999, 0.7753453, 0.7726299, 0.7692825, 
    0.7689294, 0.7670214, 0.770174, 0.7671434, 0.7792436, 0.7736239, 
    0.7898353, 0.7856631, 0.7875648, 0.7896854, 0.7832576, 0.776798, 
    0.7766644, 0.7746828, 0.7693317, 0.7787421, 0.7530367, 0.7677136, 
    0.8411073, 0.7900548, 0.7891413, 0.7916339, 0.775686, 0.781199, 
    0.7670674, 0.7706596, 0.7648642, 0.7676861, 0.7681109, 0.7719244, 
    0.7743921, 0.7809395, 0.7865893, 0.7912694, 0.7901656, 0.7850788, 
    0.7764161, 0.7688975, 0.7704868, 0.7652883, 0.7798414, 0.7734301, 
    0.7758562, 0.7696698, 0.7838053, 0.7716322, 0.7871597, 0.7857032, 
    0.7813115, 0.7730112, 0.7712736, 0.7694585, 0.7705736, 0.7762057, 
    0.7771633, 0.7814162, 0.7826219, 0.7860188, 0.7889075, 0.7862655, 
    0.7835529, 0.7762032, 0.7700406, 0.7638372, 0.7624031, 0.7560232, 
    0.7611579, 0.7529663, 0.7598404, 0.7486077, 0.7709745, 0.7600581, 
    0.7811158, 0.7785761, 0.7741443, 0.7647902, 0.7696978, 0.7639921, 
    0.7772009, 0.7849071, 0.786992, 0.7909799, 0.7869024, 0.787229, 0.783442, 
    0.7846455, 0.7759683, 0.7805386, 0.7681217, 0.7640354, 0.7538456, 
    0.7486254, 0.7441486, 0.7424484, 0.7419651, 0.7417678,
  1.19218, 1.192447, 1.192423, 1.192433, 1.192456, 1.192421, 1.192263, 
    1.19245, 1.192359, 1.192219, 1.191749, 1.192428, 1.229152, 1.235591, 
    1.219169, 1.230162, 1.216908, 1.219492, 1.211657, 1.21392, 1.203696, 
    1.210607, 1.198278, 1.20536, 1.204261, 1.210833, 1.192364, 1.191884, 
    1.19238, 1.19234, 1.192359, 1.192457, 1.192416, 1.192146, 1.192214, 
    1.192403, 1.192319, 1.192431, 1.191982, 1.191998, 1.233233, 1.237194, 
    1.222179, 1.226517, 1.213826, 1.217063, 1.213979, 1.214917, 1.213966, 
    1.218701, 1.216681, 1.220818, 1.236455, 1.231936, 1.192253, 1.192451, 
    1.192276, 1.192011, 1.192055, 1.192133, 1.192404, 1.192449, 1.192342, 
    1.192199, 1.192001, 1.234508, 1.230486, 1.221295, 1.222973, 1.220126, 
    1.217383, 1.212728, 1.213499, 1.211432, 1.220202, 1.214398, 1.223925, 
    1.221346, 1.191936, 1.192409, 1.192457, 1.192428, 1.192088, 1.192363, 
    1.192275, 1.192438, 1.192456, 1.192455, 1.192194, 1.192372, 1.230246, 
    1.237815, 1.217704, 1.22263, 1.216513, 1.219648, 1.214258, 1.219113, 
    1.210659, 1.20879, 1.210069, 1.205133, 1.21938, 1.213978, 1.192455, 
    1.192456, 1.192457, 1.192385, 1.192374, 1.192144, 1.192356, 1.192411, 
    1.192455, 1.192414, 1.192327, 1.191971, 1.236092, 1.228144, 1.222312, 
    1.218346, 1.220784, 1.218632, 1.221036, 1.222158, 1.209491, 1.216662, 
    1.205847, 1.206455, 1.211382, 1.206386, 1.192457, 1.192445, 1.192294, 
    1.192427, 1.19211, 1.192329, 1.192407, 1.192369, 1.192286, 1.192185, 
    1.191913, 1.236992, 1.229711, 1.223241, 1.217223, 1.217668, 1.217511, 
    1.216153, 1.219507, 1.215599, 1.214939, 1.216663, 1.206536, 1.20946, 
    1.206467, 1.208374, 1.192451, 1.192454, 1.192457, 1.192442, 1.192457, 
    1.192224, 1.192069, 1.233061, 1.237073, 1.230666, 1.236428, 1.235414, 
    1.230453, 1.236119, 1.2236, 1.232139, 1.2161, 1.224818, 1.215546, 
    1.21725, 1.214425, 1.211875, 1.20864, 1.20259, 1.204001, 1.198881, 
    1.192384, 1.192245, 1.192261, 1.192045, 1.191833, 1.23559, 1.227875, 
    1.230798, 1.225412, 1.22432, 1.232495, 1.227499, 1.192112, 1.191881, 
    1.192026, 1.192375, 1.230126, 1.19171, 1.222215, 1.227299, 1.21224, 
    1.219813, 1.204775, 1.19814, 1.191782, 1.184205, 1.192139, 1.192268, 
    1.192014, 1.237408, 1.232978, 1.226991, 1.226373, 1.225237, 1.222277, 
    1.219767, 1.224876, 1.219135, 1.191818, 1.229323, 1.192308, 1.191925, 
    1.237688, 1.19171, 1.23113, 1.22919, 1.221188, 1.225349, 1.199788, 
    1.211333, 1.178331, 1.187862, 1.192305, 1.19214, 1.234692, 1.191678, 
    1.226588, 1.223468, 1.22091, 1.21761, 1.217252, 1.21528, 1.218506, 
    1.215408, 1.226979, 1.221857, 1.235724, 1.232403, 1.233935, 1.235608, 
    1.230418, 1.224796, 1.224676, 1.222852, 1.217657, 1.226537, 1.198269, 
    1.216, 1.191889, 1.235894, 1.235182, 1.237112, 1.223782, 1.228675, 
    1.215328, 1.218988, 1.212971, 1.215974, 1.216414, 1.220228, 1.222581, 
    1.228452, 1.233153, 1.236833, 1.235981, 1.231925, 1.22445, 1.217219, 
    1.218817, 1.213432, 1.227502, 1.221673, 1.223938, 1.218001, 1.230875, 
    1.219941, 1.233612, 1.232436, 1.228771, 1.221274, 1.219593, 1.217788, 
    1.218903, 1.224258, 1.225127, 1.228861, 1.229884, 1.232692, 1.234998, 
    1.232892, 1.230664, 1.224256, 1.218372, 1.211838, 1.210221, 1.202386, 
    1.208776, 1.198167, 1.207205, 1.191412, 1.219298, 1.207469, 1.228604, 
    1.22639, 1.222347, 1.212889, 1.218029, 1.21201, 1.225161, 1.231784, 
    1.233477, 1.236611, 1.233405, 1.233667, 1.230572, 1.23157, 1.224041, 
    1.228107, 1.216425, 1.212058, 1.199421, 1.191443, 1.183138, 1.179411, 
    1.178269, 1.177791,
  0.5002619, 0.4900357, 0.4920214, 0.4837911, 0.4883544, 0.4829688, 
    0.4981866, 0.4896299, 0.49509, 0.4993407, 0.4678833, 0.4834246, 
    0.4518843, 0.4617273, 0.4370832, 0.4534127, 0.433806, 0.4375536, 
    0.4262982, 0.4295161, 0.41519, 0.4248148, 0.4078108, 0.4174845, 
    0.4159672, 0.425133, 0.4802912, 0.4698131, 0.480913, 0.4794161, 
    0.4800879, 0.4882597, 0.4923853, 0.5010455, 0.4994718, 0.4931123, 
    0.4787433, 0.4836141, 0.4713566, 0.4716329, 0.4580955, 0.4642133, 
    0.4414889, 0.4479249, 0.4293817, 0.4340291, 0.4295996, 0.4309418, 
    0.4295821, 0.4364026, 0.4334774, 0.4394898, 0.4630661, 0.4561119, 
    0.4768549, 0.4894285, 0.4978107, 0.5037705, 0.5029273, 0.5013203, 
    0.4930751, 0.4853427, 0.4794628, 0.4755361, 0.4716726, 0.4600558, 
    0.4539045, 0.4401893, 0.442659, 0.4384776, 0.4344921, 0.4278175, 
    0.4289147, 0.4259794, 0.4385885, 0.4301991, 0.4440669, 0.4402645, 
    0.4706196, 0.4822994, 0.487275, 0.4916395, 0.5022791, 0.4949278, 
    0.4978238, 0.490939, 0.4865714, 0.4887309, 0.4754288, 0.480593, 
    0.4535404, 0.4651818, 0.4349566, 0.442152, 0.4332358, 0.4377809, 
    0.4299992, 0.4370013, 0.4248884, 0.4222606, 0.4240559, 0.4171704, 
    0.4373901, 0.4295993, 0.4887913, 0.4884389, 0.4867984, 0.4940161, 
    0.4944583, 0.5010884, 0.4951886, 0.4926791, 0.4863186, 0.4825619, 
    0.4789954, 0.4711694, 0.4625027, 0.4503648, 0.4416847, 0.4358858, 
    0.43944, 0.4363018, 0.4398101, 0.4414566, 0.4232446, 0.4334499, 
    0.4181591, 0.4190021, 0.4259095, 0.418907, 0.4881916, 0.4902194, 
    0.4972686, 0.4917507, 0.5018113, 0.4961757, 0.4929393, 0.4804842, 
    0.4777555, 0.4752265, 0.4702392, 0.4638997, 0.4527294, 0.4430543, 
    0.4342606, 0.4349037, 0.4346773, 0.4327172, 0.4375754, 0.4319208, 
    0.430973, 0.4334516, 0.4191149, 0.4231997, 0.41902, 0.4216785, 0.4895602, 
    0.4861498, 0.4879921, 0.4845284, 0.4869679, 0.4761346, 0.4728945, 
    0.4578323, 0.4640252, 0.4541776, 0.4630233, 0.4614534, 0.4538555, 
    0.4625447, 0.443586, 0.4564213, 0.4326411, 0.4453921, 0.4318446, 
    0.4342986, 0.4302376, 0.4266073, 0.4220508, 0.4136721, 0.4156089, 
    0.4086256, 0.4810729, 0.4766623, 0.477051, 0.4724425, 0.4690391, 
    0.4617253, 0.4499598, 0.4543775, 0.4462747, 0.4446514, 0.4569643, 
    0.4493958, 0.4737148, 0.4697624, 0.4721155, 0.4807243, 0.4533578, 
    0.4673448, 0.4415414, 0.4490962, 0.4271244, 0.4380214, 0.4166759, 
    0.4076252, 0.3991553, 0.3893117, 0.4742588, 0.4772523, 0.4718952, 
    0.4645476, 0.4577039, 0.4486346, 0.4477091, 0.4460145, 0.4416322, 
    0.4379542, 0.4454783, 0.4370333, 0.4688452, 0.4521436, 0.4783843, 
    0.4704408, 0.4649835, 0.4673496, 0.4548831, 0.4519425, 0.4400321, 
    0.4461814, 0.4098539, 0.4258404, 0.3818632, 0.3940289, 0.4782988, 
    0.4742694, 0.4603378, 0.4669329, 0.4480308, 0.4433894, 0.4396242, 
    0.43482, 0.4343025, 0.4314622, 0.4361185, 0.4316462, 0.4486153, 
    0.4410153, 0.4619332, 0.4568241, 0.4591734, 0.4617524, 0.4538015, 
    0.4453595, 0.4451806, 0.4424804, 0.4348883, 0.4479543, 0.4077992, 
    0.4324973, 0.4698821, 0.462196, 0.4610942, 0.4640868, 0.4438542, 
    0.4511647, 0.4315315, 0.4368197, 0.4281628, 0.4324598, 0.4330927, 
    0.4386272, 0.4420801, 0.4508288, 0.4579723, 0.4636527, 0.4623308, 
    0.4560951, 0.4448444, 0.4342551, 0.43657, 0.4288194, 0.4493997, 
    0.4407447, 0.4440854, 0.435386, 0.4544948, 0.4382084, 0.4586761, 
    0.4568745, 0.45131, 0.4401582, 0.4377004, 0.4350774, 0.4366958, 
    0.4445597, 0.4458514, 0.4514454, 0.4529918, 0.4572667, 0.4608111, 
    0.4575722, 0.4541752, 0.4445569, 0.4359247, 0.4265555, 0.42427, 
    0.4133928, 0.4222409, 0.4076624, 0.4200468, 0.3986678, 0.43727, 
    0.4204146, 0.4510575, 0.4477349, 0.4417365, 0.4280463, 0.4354268, 
    0.4267987, 0.445902, 0.4558797, 0.4584696, 0.4633068, 0.4583591, 
    0.4587612, 0.4540354, 0.4555531, 0.4442382, 0.4503091, 0.4331083, 
    0.426867, 0.4093557, 0.3987088, 0.3879471, 0.3832206, 0.3817853, 0.3811857,
  0.04899819, 0.04713374, 0.04749282, 0.04601381, 0.04683083, 0.04586738, 
    0.04861675, 0.04706054, 0.04805052, 0.04882867, 0.04322414, 0.04594852, 
    0.04050252, 0.0421609, 0.03807338, 0.04075778, 0.03754598, 0.03814939, 
    0.03635197, 0.03686131, 0.03462163, 0.03611841, 0.03349596, 0.0349755, 
    0.03474128, 0.03616845, 0.04539225, 0.04355772, 0.04550235, 0.04523754, 
    0.04535629, 0.0468138, 0.04755877, 0.04914261, 0.04885279, 0.04769069, 
    0.04511877, 0.04598226, 0.0438255, 0.04387351, 0.04154499, 0.04258519, 
    0.03878835, 0.03984511, 0.03683997, 0.03758177, 0.03687457, 0.03708814, 
    0.0368718, 0.03796354, 0.03749331, 0.03846309, 0.04238913, 0.04121059, 
    0.04478628, 0.04702424, 0.04854783, 0.0496466, 0.04949037, 0.04919332, 
    0.04768394, 0.04629076, 0.04524578, 0.04455484, 0.04388041, 0.04187685, 
    0.04084009, 0.03857674, 0.0389794, 0.03829893, 0.03765609, 0.036592, 
    0.03676584, 0.03630172, 0.03831689, 0.03696989, 0.03920989, 0.03858897, 
    0.04369752, 0.04574835, 0.04663689, 0.04742365, 0.04937043, 0.04802095, 
    0.04855023, 0.04729691, 0.0465107, 0.04689857, 0.04453604, 0.04544568, 
    0.04077915, 0.04275108, 0.03773071, 0.03889655, 0.03745461, 0.03818614, 
    0.0369381, 0.03806015, 0.03612998, 0.03571803, 0.03599921, 0.03492695, 
    0.03812296, 0.03687452, 0.04690944, 0.04684603, 0.0465514, 0.04785495, 
    0.04793543, 0.04915054, 0.0480685, 0.04761206, 0.04646542, 0.04579501, 
    0.04516324, 0.04379297, 0.04229302, 0.04024958, 0.03882029, 0.03788025, 
    0.03845499, 0.03794729, 0.0385151, 0.03878309, 0.035872, 0.03748891, 
    0.0350799, 0.03521057, 0.0362907, 0.03519583, 0.04680155, 0.04716691, 
    0.04844854, 0.04744379, 0.04928398, 0.04824866, 0.04765928, 0.04542642, 
    0.04494468, 0.04450059, 0.04363155, 0.04253156, 0.04064355, 0.03904405, 
    0.03761892, 0.03772222, 0.03768583, 0.0373716, 0.03815292, 0.03724431, 
    0.03709311, 0.03748917, 0.03522809, 0.03586497, 0.03521335, 0.0356271, 
    0.04704798, 0.04643517, 0.04676569, 0.0461453, 0.0465818, 0.0446598, 
    0.04409314, 0.04150055, 0.04255301, 0.04088583, 0.04238182, 0.04211428, 
    0.04083189, 0.04230017, 0.03913108, 0.04126265, 0.03735942, 0.03942751, 
    0.03723214, 0.03762501, 0.03697601, 0.03640075, 0.03568524, 0.03438852, 
    0.03468609, 0.03361932, 0.04553069, 0.04475244, 0.04482074, 0.04401438, 
    0.04342376, 0.04216056, 0.0401823, 0.04091933, 0.03957278, 0.03930579, 
    0.04135412, 0.04008869, 0.04423625, 0.04354894, 0.04395745, 0.04546893, 
    0.0407486, 0.04313128, 0.03879692, 0.04003903, 0.0364824, 0.03822507, 
    0.03485058, 0.03346789, 0.03219975, 0.03075721, 0.04433127, 0.04485614, 
    0.04391912, 0.04264243, 0.04147886, 0.03996255, 0.03980944, 0.03952992, 
    0.03881172, 0.03821419, 0.03944168, 0.03806532, 0.04339025, 0.04054578, 
    0.04505546, 0.04366651, 0.0427171, 0.04313211, 0.04100413, 0.04051222, 
    0.03855118, 0.0395574, 0.03380572, 0.03627982, 0.02968791, 0.03144431, 
    0.04504039, 0.04433313, 0.04192471, 0.04306034, 0.03986263, 0.03909888, 
    0.03848491, 0.03770876, 0.03762564, 0.03717111, 0.03791775, 0.03720047, 
    0.03995935, 0.03871116, 0.04219595, 0.04133049, 0.0417273, 0.04216517, 
    0.04082284, 0.03942214, 0.03939272, 0.03895021, 0.03771975, 0.03984999, 
    0.03349421, 0.03733642, 0.04356968, 0.04224072, 0.0420532, 0.04256355, 
    0.03917503, 0.04038263, 0.03718217, 0.03803084, 0.03664667, 0.03733043, 
    0.03743169, 0.03832317, 0.03888482, 0.04032672, 0.04152419, 0.04248932, 
    0.0422637, 0.04120776, 0.03933749, 0.03761804, 0.03799054, 0.03675073, 
    0.04008935, 0.0386671, 0.03921293, 0.03779977, 0.04093899, 0.03825534, 
    0.04164314, 0.04133898, 0.04040683, 0.03857167, 0.03817313, 0.03775014, 
    0.03801084, 0.03929075, 0.03950306, 0.04042937, 0.0406874, 0.0414051, 
    0.04200508, 0.04145664, 0.04088543, 0.03929028, 0.03788651, 0.03639257, 
    0.03603282, 0.03434571, 0.03571495, 0.03347352, 0.03537287, 0.03212753, 
    0.03810357, 0.03543009, 0.04036479, 0.03981371, 0.03882874, 0.03662823, 
    0.03780634, 0.03643096, 0.0395114, 0.04117153, 0.04160822, 0.04243022, 
    0.04158955, 0.04165754, 0.04086201, 0.04111663, 0.03923799, 0.04024032, 
    0.03743419, 0.03644174, 0.03373006, 0.03213359, 0.03055988, 0.02988136, 
    0.02967683, 0.02959159,
  0.001314405, 0.001238281, 0.001252822, 0.001193305, 0.00122606, 
    0.001187466, 0.001298705, 0.001235324, 0.001275519, 0.00130742, 
    0.001083766, 0.0011907, 0.0009804169, 0.001042971, 0.0008912049, 
    0.0009899591, 0.0008722227, 0.0008939523, 0.0008297676, 0.0008477895, 
    0.0007695429, 0.0008215479, 0.0007317304, 0.0007817327, 0.0007736571, 
    0.0008233066, 0.001168588, 0.001096674, 0.001172954, 0.001162464, 
    0.001167164, 0.001225375, 0.001255499, 0.001320365, 0.001308413, 
    0.001260859, 0.00115777, 0.001192046, 0.001107074, 0.001108942, 
    0.001019585, 0.001059186, 0.0009171605, 0.0009559871, 0.0008470315, 
    0.0008735065, 0.0008482604, 0.0008558577, 0.0008481618, 0.0008872399, 
    0.0008703347, 0.0009053209, 0.001051683, 0.001006964, 0.001144662, 
    0.001233859, 0.001295875, 0.001341239, 0.001334756, 0.001322461, 
    0.001260584, 0.001204374, 0.00116279, 0.001135569, 0.001109211, 
    0.001032163, 0.0009930431, 0.0009094519, 0.0009241388, 0.0008993655, 
    0.0008761741, 0.0008382439, 0.0008444012, 0.0008279966, 0.0009000166, 
    0.0008516483, 0.0009325822, 0.0009098966, 0.0011021, 0.001182728, 
    0.001218258, 0.001250016, 0.001329787, 0.001274312, 0.001295974, 
    0.001244881, 0.00121319, 0.00122879, 0.001134831, 0.001170706, 
    0.0009907595, 0.00106555, 0.0008788558, 0.0009211104, 0.0008689482, 
    0.0008952817, 0.0008505178, 0.0008907272, 0.0008219545, 0.0008075231, 
    0.0008173638, 0.0007800563, 0.0008929967, 0.0008482586, 0.001229228, 
    0.001226673, 0.001214824, 0.001267544, 0.001270824, 0.001320693, 
    0.001276253, 0.001257663, 0.001211373, 0.001184584, 0.001159527, 
    0.001105809, 0.001048011, 0.0009709927, 0.000918326, 0.0008842378, 
    0.000905027, 0.0008866541, 0.0009072106, 0.0009169683, 0.0008129066, 
    0.000870177, 0.0007853415, 0.0007898663, 0.0008276087, 0.0007893555, 
    0.001224882, 0.001239622, 0.001291802, 0.001250833, 0.001326209, 
    0.001283616, 0.001259582, 0.001169943, 0.0011509, 0.001133441, 
    0.001099538, 0.001057132, 0.0009856853, 0.0009265045, 0.0008748397, 
    0.0008785505, 0.0008772426, 0.0008659772, 0.0008940798, 0.0008614279, 
    0.000856035, 0.0008701864, 0.0007904737, 0.0008126606, 0.0007899627, 
    0.0008043495, 0.001234817, 0.00121016, 0.001223438, 0.001198556, 
    0.001216044, 0.00113969, 0.001117502, 0.001017905, 0.001057954, 
    0.000994758, 0.001051404, 0.001041195, 0.0009927355, 0.001048284, 
    0.0009296925, 0.001008925, 0.0008655416, 0.0009405781, 0.0008609935, 
    0.0008750584, 0.0008518661, 0.0008314876, 0.0008063781, 0.0007615492, 
    0.0007717586, 0.0007353757, 0.001174078, 0.001143331, 0.001146019, 
    0.00111443, 0.001091484, 0.001042958, 0.0009684911, 0.0009960147, 
    0.0009459286, 0.0009361032, 0.001012375, 0.0009650143, 0.001123091, 
    0.001096334, 0.001112211, 0.001171628, 0.0009896153, 0.001080182, 
    0.0009174731, 0.0009631713, 0.00083437, 0.0008966902, 0.000777422, 
    0.0007307801, 0.0006883058, 0.0006410813, 0.001126808, 0.001147412, 
    0.001110718, 0.00106138, 0.001017085, 0.0009603355, 0.0009546676, 
    0.0009443489, 0.000918013, 0.0008962965, 0.0009410997, 0.0008909139, 
    0.001090187, 0.0009820318, 0.00115527, 0.001100895, 0.001064245, 
    0.001080214, 0.0009991982, 0.0009807791, 0.0009085222, 0.0009453616, 
    0.0007416895, 0.0008272253, 0.0006068415, 0.0006634283, 0.001154675, 
    0.001126881, 0.001033982, 0.001077446, 0.0009566353, 0.0009285127, 
    0.0009061136, 0.0008780666, 0.0008750809, 0.0008588157, 0.0008855889, 
    0.000859863, 0.0009602173, 0.0009143461, 0.001044308, 0.001011483, 
    0.001026489, 0.001043134, 0.0009923966, 0.0009403806, 0.0009392985, 
    0.0009230716, 0.0008784614, 0.0009561675, 0.0007316711, 0.0008647192, 
    0.001097138, 0.001046015, 0.001038869, 0.001058358, 0.0009313037, 
    0.000975946, 0.0008592103, 0.0008896688, 0.0008401788, 0.0008645048, 
    0.0008681276, 0.000900244, 0.000920682, 0.0009738635, 0.001018798, 
    0.001055515, 0.001046892, 0.001006857, 0.0009372678, 0.000874808, 
    0.0008882141, 0.0008438656, 0.0009650385, 0.0009127407, 0.000932694, 
    0.0008813398, 0.0009967524, 0.0008977863, 0.0010233, 0.001011803, 
    0.0009768481, 0.0009092676, 0.0008948109, 0.0008795542, 0.0008889465, 
    0.0009355505, 0.0009433595, 0.0009776885, 0.0009873252, 0.001014299, 
    0.001037038, 0.001016245, 0.0009947432, 0.0009355332, 0.0008844633, 
    0.0008311993, 0.0008185429, 0.0007600842, 0.0008074152, 0.0007309707, 
    0.0007954988, 0.0006859135, 0.0008922957, 0.0007974879, 0.0009752814, 
    0.0009548253, 0.0009186342, 0.0008395259, 0.0008815763, 0.0008325538, 
    0.0009436668, 0.001005493, 0.001021978, 0.001053254, 0.001021271, 
    0.001023845, 0.0009938648, 0.001003427, 0.0009336137, 0.0009706481, 
    0.0008682171, 0.0008329343, 0.0007391244, 0.0006861141, 0.0006347131, 
    0.000612987, 0.0006064902, 0.0006037899,
  8.639937e-06, 7.87812e-06, 8.021895e-06, 7.438759e-06, 7.757933e-06, 
    7.382321e-06, 8.480997e-06, 7.848987e-06, 8.247979e-06, 8.569104e-06, 
    6.403892e-06, 7.413563e-06, 5.476304e-06, 6.031866e-06, 4.716954e-06, 
    5.559854e-06, 4.560644e-06, 4.739734e-06, 4.218054e-06, 4.362281e-06, 
    3.749385e-06, 4.152871e-06, 3.143563e-06, 3.842555e-06, 3.780733e-06, 
    4.166786e-06, 7.200818e-06, 6.523161e-06, 7.242659e-06, 7.14225e-06, 
    7.187181e-06, 7.751207e-06, 8.048453e-06, 8.700531e-06, 8.579162e-06, 
    8.10172e-06, 7.097467e-06, 7.426577e-06, 6.619782e-06, 6.637189e-06, 
    5.82202e-06, 6.17884e-06, 4.933733e-06, 5.264412e-06, 4.356179e-06, 
    4.571155e-06, 4.366074e-06, 4.427427e-06, 4.365279e-06, 4.684147e-06, 
    4.545201e-06, 4.834417e-06, 6.110681e-06, 5.709825e-06, 6.972911e-06, 
    7.834558e-06, 8.452444e-06, 8.913767e-06, 8.847368e-06, 8.721859e-06, 
    8.098988e-06, 7.546135e-06, 7.145363e-06, 6.886923e-06, 6.639694e-06, 
    5.93457e-06, 5.58695e-06, 4.868989e-06, 4.992606e-06, 4.784734e-06, 
    4.593025e-06, 4.285666e-06, 4.335029e-06, 4.203978e-06, 4.790157e-06, 
    4.393394e-06, 5.06417e-06, 4.872715e-06, 6.573509e-06, 7.336622e-06, 
    7.681513e-06, 7.994088e-06, 8.796578e-06, 8.235908e-06, 8.453441e-06, 
    7.943278e-06, 7.632003e-06, 7.784727e-06, 6.879964e-06, 7.221106e-06, 
    5.566882e-06, 6.236843e-06, 4.615047e-06, 4.967027e-06, 4.533873e-06, 
    4.750772e-06, 4.38427e-06, 4.712997e-06, 4.156087e-06, 4.042529e-06, 
    4.119835e-06, 3.82969e-06, 4.731806e-06, 4.366059e-06, 7.78903e-06, 
    7.763944e-06, 7.64795e-06, 8.168309e-06, 8.201046e-06, 8.703863e-06, 
    8.255324e-06, 8.069949e-06, 7.614281e-06, 7.354518e-06, 7.114218e-06, 
    6.608006e-06, 6.077419e-06, 5.394218e-06, 4.943548e-06, 4.659361e-06, 
    4.831961e-06, 4.679307e-06, 4.850221e-06, 4.932116e-06, 4.084753e-06, 
    4.543912e-06, 3.870305e-06, 3.905207e-06, 4.200897e-06, 3.901261e-06, 
    7.746372e-06, 7.891344e-06, 8.411406e-06, 8.002179e-06, 8.760063e-06, 
    8.329119e-06, 8.089021e-06, 7.213788e-06, 7.0321e-06, 6.866854e-06, 
    6.549723e-06, 6.160154e-06, 5.522379e-06, 5.012621e-06, 4.582081e-06, 
    4.612538e-06, 4.601795e-06, 4.509634e-06, 4.740793e-06, 4.472608e-06, 
    4.428862e-06, 4.543989e-06, 3.9099e-06, 4.082819e-06, 3.905951e-06, 
    4.017715e-06, 7.843992e-06, 7.602456e-06, 7.732221e-06, 7.489633e-06, 
    7.659875e-06, 6.925848e-06, 6.71714e-06, 5.807036e-06, 6.167625e-06, 
    5.602038e-06, 6.108149e-06, 6.015837e-06, 5.584246e-06, 6.079892e-06, 
    5.039637e-06, 5.727211e-06, 4.506083e-06, 5.132271e-06, 4.469079e-06, 
    4.583873e-06, 4.395153e-06, 4.231742e-06, 4.03357e-06, 3.688763e-06, 
    3.766255e-06, 3.492965e-06, 7.25345e-06, 6.960301e-06, 6.985767e-06, 
    6.68841e-06, 6.47512e-06, 6.031747e-06, 5.372502e-06, 5.613103e-06, 
    5.178021e-06, 5.094118e-06, 5.757831e-06, 5.34237e-06, 6.769515e-06, 
    6.520007e-06, 6.667684e-06, 7.229945e-06, 5.556837e-06, 6.370909e-06, 
    4.936365e-06, 5.326421e-06, 4.254716e-06, 4.762476e-06, 3.809507e-06, 
    3.138315e-06, 2.904989e-06, 2.648534e-06, 6.804419e-06, 6.998983e-06, 
    6.65375e-06, 6.198819e-06, 5.799735e-06, 5.301914e-06, 5.25305e-06, 
    5.164499e-06, 4.940912e-06, 4.759203e-06, 5.136725e-06, 4.714543e-06, 
    6.463133e-06, 5.490413e-06, 7.073654e-06, 6.562322e-06, 6.224935e-06, 
    6.371205e-06, 5.641166e-06, 5.479467e-06, 4.8612e-06, 5.173167e-06, 
    3.539816e-06, 4.197853e-06, 2.464689e-06, 2.769487e-06, 7.067995e-06, 
    6.805102e-06, 5.950903e-06, 6.345774e-06, 5.269997e-06, 5.029633e-06, 
    4.841045e-06, 4.608563e-06, 4.584058e-06, 4.451399e-06, 4.670511e-06, 
    4.459898e-06, 5.300893e-06, 4.910059e-06, 6.043933e-06, 5.749913e-06, 
    5.883701e-06, 6.033335e-06, 5.581267e-06, 5.130585e-06, 5.121352e-06, 
    4.983586e-06, 4.611806e-06, 5.265966e-06, 3.143235e-06, 4.499383e-06, 
    6.52746e-06, 6.059367e-06, 5.994871e-06, 6.171299e-06, 5.05331e-06, 
    5.437308e-06, 4.4546e-06, 4.704234e-06, 4.301155e-06, 4.497638e-06, 
    4.527174e-06, 4.792052e-06, 4.963412e-06, 5.419178e-06, 5.815004e-06, 
    6.14546e-06, 6.067294e-06, 5.708881e-06, 5.104039e-06, 4.58182e-06, 
    4.6922e-06, 4.330726e-06, 5.34258e-06, 4.896574e-06, 5.06512e-06, 
    4.635482e-06, 5.619602e-06, 4.77159e-06, 5.855183e-06, 5.752755e-06, 
    5.445168e-06, 4.867444e-06, 4.746862e-06, 4.62079e-06, 4.698257e-06, 
    5.089414e-06, 5.156036e-06, 5.452495e-06, 5.536748e-06, 5.774934e-06, 
    5.978386e-06, 5.792258e-06, 5.601908e-06, 5.089267e-06, 4.661221e-06, 
    4.229446e-06, 4.129136e-06, 3.677695e-06, 4.041685e-06, 3.139367e-06, 
    3.948817e-06, 2.891921e-06, 4.725993e-06, 3.964263e-06, 5.43152e-06, 
    5.254408e-06, 4.946145e-06, 4.295926e-06, 4.637428e-06, 4.240234e-06, 
    5.158665e-06, 5.696801e-06, 5.843371e-06, 6.124931e-06, 5.83706e-06, 
    5.860056e-06, 5.594179e-06, 5.678521e-06, 5.072937e-06, 5.391225e-06, 
    4.527904e-06, 4.243267e-06, 3.520752e-06, 2.893016e-06, 2.614204e-06, 
    2.49755e-06, 2.462813e-06, 2.448394e-06,
  7.925912e-09, 6.761332e-09, 6.978174e-09, 6.107835e-09, 6.581175e-09, 
    6.024933e-09, 7.679854e-09, 6.717568e-09, 7.321993e-09, 7.816062e-09, 
    4.62956e-09, 6.070795e-09, 3.392006e-09, 4.122109e-09, 2.457013e-09, 
    3.499521e-09, 2.275023e-09, 2.483859e-09, 1.890551e-09, 2.049894e-09, 
    1.400802e-09, 1.819798e-09, 1.122341e-09, 1.494503e-09, 1.432113e-09, 
    1.834834e-09, 5.760004e-09, 4.795123e-09, 5.820846e-09, 5.675076e-09, 
    5.740205e-09, 6.571121e-09, 7.018385e-09, 8.020127e-09, 7.83164e-09, 
    7.099178e-09, 5.610325e-09, 6.089919e-09, 4.930225e-09, 4.954655e-09, 
    3.842235e-09, 4.320914e-09, 2.715675e-09, 3.123232e-09, 2.043077e-09, 
    2.287137e-09, 2.054135e-09, 2.123087e-09, 2.053246e-09, 2.418493e-09, 
    2.257258e-09, 2.596295e-09, 4.22844e-09, 3.694597e-09, 5.431103e-09, 
    6.695915e-09, 7.635818e-09, 8.353427e-09, 8.249355e-09, 8.053343e-09, 
    7.09503e-09, 6.266231e-09, 5.679583e-09, 5.308137e-09, 4.958173e-09, 
    3.99175e-09, 3.53457e-09, 2.637685e-09, 2.787121e-09, 2.537127e-09, 
    2.3124e-09, 1.964778e-09, 2.019498e-09, 1.875204e-09, 2.543566e-09, 
    2.084757e-09, 2.874632e-09, 2.642157e-09, 4.865415e-09, 5.957986e-09, 
    6.467159e-09, 6.936124e-09, 8.169922e-09, 7.30355e-09, 7.637355e-09, 
    6.859427e-09, 6.393519e-09, 6.621249e-09, 5.298212e-09, 5.789489e-09, 
    3.508603e-09, 4.39998e-09, 2.337919e-09, 2.756018e-09, 2.244251e-09, 
    2.496896e-09, 2.074517e-09, 2.452359e-09, 1.823269e-09, 1.701894e-09, 
    1.784249e-09, 1.481451e-09, 2.474507e-09, 2.054118e-09, 6.627689e-09, 
    6.59016e-09, 6.41722e-09, 7.200446e-09, 7.250339e-09, 8.025316e-09, 
    7.33322e-09, 7.050966e-09, 6.367205e-09, 5.984182e-09, 5.634526e-09, 
    4.913712e-09, 4.183487e-09, 3.28721e-09, 2.727552e-09, 2.389505e-09, 
    2.593361e-09, 2.412824e-09, 2.615194e-09, 2.713719e-09, 1.74673e-09, 
    2.255777e-09, 1.522779e-09, 1.558577e-09, 1.87185e-09, 1.554517e-09, 
    6.563899e-09, 6.781216e-09, 7.572616e-09, 6.948354e-09, 8.112907e-09, 
    7.446209e-09, 7.079899e-09, 5.77885e-09, 5.516109e-09, 5.279527e-09, 
    4.832179e-09, 4.295515e-09, 3.451192e-09, 2.811523e-09, 2.299748e-09, 
    2.335008e-09, 2.322553e-09, 2.216492e-09, 2.485109e-09, 2.174281e-09, 
    2.124707e-09, 2.255865e-09, 1.563411e-09, 1.744669e-09, 1.559344e-09, 
    1.675712e-09, 6.71007e-09, 6.349658e-09, 6.542766e-09, 6.182773e-09, 
    6.434955e-09, 5.363722e-09, 5.067218e-09, 3.822436e-09, 4.305666e-09, 
    3.554125e-09, 4.225014e-09, 4.100564e-09, 3.531069e-09, 4.186826e-09, 
    2.844551e-09, 3.717382e-09, 2.212434e-09, 2.95857e-09, 2.170269e-09, 
    2.301819e-09, 2.086734e-09, 1.905509e-09, 1.692427e-09, 1.340884e-09, 
    1.417625e-09, 1.153304e-09, 5.836561e-09, 5.41303e-09, 5.44954e-09, 
    5.026703e-09, 4.728274e-09, 4.12195e-09, 3.259627e-09, 3.568482e-09, 
    3.015315e-09, 2.911466e-09, 3.757594e-09, 3.221454e-09, 5.141268e-09, 
    4.790729e-09, 4.997521e-09, 5.802344e-09, 3.495624e-09, 4.584015e-09, 
    2.718858e-09, 3.201296e-09, 1.930695e-09, 2.51074e-09, 1.461047e-09, 
    1.11589e-09, 8.457931e-10, 5.886177e-10, 5.190749e-09, 5.46851e-09, 
    4.977923e-09, 4.34811e-09, 3.812797e-09, 3.170384e-09, 3.108984e-09, 
    2.998514e-09, 2.72436e-09, 2.506866e-09, 2.964082e-09, 2.454177e-09, 
    4.711627e-09, 3.410102e-09, 5.575961e-09, 4.849776e-09, 4.38372e-09, 
    4.584423e-09, 3.604962e-09, 3.396061e-09, 2.628345e-09, 3.009281e-09, 
    1.197335e-09, 1.868538e-09, 4.315928e-10, 7.045379e-10, 5.567802e-09, 
    5.191719e-09, 4.013562e-09, 4.549377e-09, 3.130242e-09, 2.832308e-09, 
    2.604216e-09, 2.330397e-09, 2.302033e-09, 2.150205e-09, 2.402533e-09, 
    2.159844e-09, 3.169098e-09, 2.687087e-09, 4.138348e-09, 3.747186e-09, 
    3.924002e-09, 4.124085e-09, 3.527211e-09, 2.956484e-09, 2.945069e-09, 
    2.776142e-09, 2.334158e-09, 3.125182e-09, 1.121937e-09, 2.204782e-09, 
    4.801117e-09, 4.159137e-09, 4.072424e-09, 4.310659e-09, 2.861306e-09, 
    3.342117e-09, 2.153834e-09, 2.442059e-09, 1.981901e-09, 2.202791e-09, 
    2.236569e-09, 2.545818e-09, 2.75163e-09, 3.318987e-09, 3.832961e-09, 
    4.275567e-09, 4.169826e-09, 3.693362e-09, 2.923695e-09, 2.299447e-09, 
    2.427933e-09, 2.014711e-09, 3.221719e-09, 2.670838e-09, 2.875798e-09, 
    2.361667e-09, 3.576922e-09, 2.521535e-09, 3.886145e-09, 3.75092e-09, 
    3.352158e-09, 2.635832e-09, 2.492275e-09, 2.344586e-09, 2.435041e-09, 
    2.905671e-09, 2.988011e-09, 3.361524e-09, 3.469703e-09, 3.780101e-09, 
    4.050331e-09, 3.802932e-09, 3.553955e-09, 2.90549e-09, 2.391676e-09, 
    1.902998e-09, 1.794235e-09, 1.330035e-09, 1.701001e-09, 1.117182e-09, 
    1.603669e-09, 8.316579e-10, 2.467656e-09, 1.619735e-09, 3.334728e-09, 
    3.110685e-09, 2.730697e-09, 1.976115e-09, 2.363933e-09, 1.914808e-09, 
    2.991273e-09, 3.677552e-09, 3.870491e-09, 4.247734e-09, 3.862134e-09, 
    3.892607e-09, 3.543935e-09, 3.653662e-09, 2.885402e-09, 3.283405e-09, 
    2.237406e-09, 1.918131e-09, 1.179352e-09, 8.328389e-10, 5.575134e-10, 
    4.579189e-10, 4.301126e-10, 4.188245e-10,
  4.321133e-13, 4.275416e-13, 4.283935e-13, 4.249726e-13, 4.268336e-13, 
    4.246465e-13, 4.31148e-13, 4.273696e-13, 4.297435e-13, 4.316824e-13, 
    4.191504e-13, 4.248269e-13, 4.142626e-13, 4.171478e-13, 4.105605e-13, 
    4.146878e-13, 4.098387e-13, 4.10667e-13, 4.083124e-13, 4.089452e-13, 
    4.063649e-13, 4.080313e-13, 4.052611e-13, 4.067378e-13, 4.064895e-13, 
    4.08091e-13, 4.236041e-13, 4.198033e-13, 4.238435e-13, 4.232698e-13, 
    4.235262e-13, 4.267942e-13, 4.285514e-13, 4.324828e-13, 4.317435e-13, 
    4.288687e-13, 4.230149e-13, 4.249021e-13, 4.203359e-13, 4.204322e-13, 
    4.160424e-13, 4.179326e-13, 4.115857e-13, 4.131993e-13, 4.089182e-13, 
    4.098868e-13, 4.089621e-13, 4.092358e-13, 4.089586e-13, 4.104078e-13, 
    4.097682e-13, 4.111126e-13, 4.175676e-13, 4.15459e-13, 4.223093e-13, 
    4.272846e-13, 4.309752e-13, 4.337896e-13, 4.333816e-13, 4.32613e-13, 
    4.288524e-13, 4.255955e-13, 4.232875e-13, 4.21825e-13, 4.20446e-13, 
    4.166331e-13, 4.148264e-13, 4.112767e-13, 4.118687e-13, 4.108781e-13, 
    4.09987e-13, 4.086073e-13, 4.088246e-13, 4.082514e-13, 4.109037e-13, 
    4.090837e-13, 4.122153e-13, 4.112944e-13, 4.200804e-13, 4.243831e-13, 
    4.263855e-13, 4.282283e-13, 4.330702e-13, 4.296711e-13, 4.309813e-13, 
    4.27927e-13, 4.26096e-13, 4.269912e-13, 4.217859e-13, 4.237201e-13, 
    4.147238e-13, 4.182447e-13, 4.100882e-13, 4.117455e-13, 4.097166e-13, 
    4.107186e-13, 4.09043e-13, 4.105421e-13, 4.080451e-13, 4.075627e-13, 
    4.0789e-13, 4.066859e-13, 4.106299e-13, 4.08962e-13, 4.270165e-13, 
    4.26869e-13, 4.261892e-13, 4.292663e-13, 4.294622e-13, 4.325031e-13, 
    4.297876e-13, 4.286793e-13, 4.259926e-13, 4.244862e-13, 4.231102e-13, 
    4.202708e-13, 4.173902e-13, 4.138481e-13, 4.116327e-13, 4.102928e-13, 
    4.11101e-13, 4.103853e-13, 4.111875e-13, 4.115779e-13, 4.077409e-13, 
    4.097624e-13, 4.068503e-13, 4.069927e-13, 4.082381e-13, 4.069766e-13, 
    4.267657e-13, 4.276197e-13, 4.307272e-13, 4.282763e-13, 4.328466e-13, 
    4.302311e-13, 4.28793e-13, 4.236783e-13, 4.22644e-13, 4.217123e-13, 
    4.199494e-13, 4.178324e-13, 4.144967e-13, 4.119653e-13, 4.099368e-13, 
    4.100767e-13, 4.100273e-13, 4.096065e-13, 4.106719e-13, 4.09439e-13, 
    4.092422e-13, 4.097627e-13, 4.07012e-13, 4.077327e-13, 4.069958e-13, 
    4.074586e-13, 4.273402e-13, 4.259236e-13, 4.266827e-13, 4.252674e-13, 
    4.262589e-13, 4.220439e-13, 4.208758e-13, 4.159642e-13, 4.178725e-13, 
    4.149037e-13, 4.175541e-13, 4.170628e-13, 4.148126e-13, 4.174034e-13, 
    4.120961e-13, 4.155491e-13, 4.095904e-13, 4.125476e-13, 4.094231e-13, 
    4.09945e-13, 4.090915e-13, 4.083718e-13, 4.07525e-13, 4.061264e-13, 
    4.064319e-13, 4.053792e-13, 4.239054e-13, 4.222381e-13, 4.223819e-13, 
    4.207161e-13, 4.195397e-13, 4.171472e-13, 4.13739e-13, 4.149605e-13, 
    4.127722e-13, 4.123611e-13, 4.15708e-13, 4.135879e-13, 4.211676e-13, 
    4.19786e-13, 4.206011e-13, 4.237707e-13, 4.146724e-13, 4.189707e-13, 
    4.115983e-13, 4.135082e-13, 4.084719e-13, 4.107735e-13, 4.066047e-13, 
    4.052353e-13, 4.041568e-13, 4.031284e-13, 4.213625e-13, 4.224566e-13, 
    4.205239e-13, 4.1804e-13, 4.159261e-13, 4.133859e-13, 4.131429e-13, 
    4.127057e-13, 4.116201e-13, 4.107582e-13, 4.125694e-13, 4.105493e-13, 
    4.19474e-13, 4.143342e-13, 4.228796e-13, 4.200188e-13, 4.181805e-13, 
    4.189723e-13, 4.151047e-13, 4.142787e-13, 4.112396e-13, 4.127483e-13, 
    4.055546e-13, 4.082249e-13, 4.024998e-13, 4.035921e-13, 4.228475e-13, 
    4.213664e-13, 4.167192e-13, 4.188341e-13, 4.132271e-13, 4.120476e-13, 
    4.11144e-13, 4.100584e-13, 4.099459e-13, 4.093435e-13, 4.103445e-13, 
    4.093817e-13, 4.133808e-13, 4.114724e-13, 4.17212e-13, 4.156668e-13, 
    4.163655e-13, 4.171556e-13, 4.147973e-13, 4.125394e-13, 4.124941e-13, 
    4.118252e-13, 4.100733e-13, 4.13207e-13, 4.052594e-13, 4.0956e-13, 
    4.198269e-13, 4.17294e-13, 4.169517e-13, 4.178922e-13, 4.121625e-13, 
    4.140653e-13, 4.093579e-13, 4.105012e-13, 4.086753e-13, 4.095521e-13, 
    4.096862e-13, 4.109126e-13, 4.117281e-13, 4.139738e-13, 4.160058e-13, 
    4.177537e-13, 4.173363e-13, 4.154542e-13, 4.124095e-13, 4.099356e-13, 
    4.104452e-13, 4.088055e-13, 4.13589e-13, 4.11408e-13, 4.122199e-13, 
    4.101824e-13, 4.149939e-13, 4.108163e-13, 4.162159e-13, 4.156816e-13, 
    4.14105e-13, 4.112693e-13, 4.107003e-13, 4.101147e-13, 4.104734e-13, 
    4.123382e-13, 4.126642e-13, 4.141421e-13, 4.145699e-13, 4.157969e-13, 
    4.168644e-13, 4.158872e-13, 4.149031e-13, 4.123375e-13, 4.103014e-13, 
    4.083618e-13, 4.079297e-13, 4.060832e-13, 4.075591e-13, 4.052405e-13, 
    4.071721e-13, 4.041003e-13, 4.106027e-13, 4.07236e-13, 4.140361e-13, 
    4.131497e-13, 4.116452e-13, 4.086523e-13, 4.101914e-13, 4.084088e-13, 
    4.126771e-13, 4.153917e-13, 4.161541e-13, 4.176438e-13, 4.16121e-13, 
    4.162414e-13, 4.148635e-13, 4.152972e-13, 4.122579e-13, 4.138331e-13, 
    4.096895e-13, 4.08422e-13, 4.05483e-13, 4.041051e-13, 4.03004e-13, 
    4.026052e-13, 4.024938e-13, 4.024486e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC =
  9.300609e-07, 9.300608e-07, 9.300609e-07, 9.300608e-07, 9.300608e-07, 
    9.300608e-07, 9.300609e-07, 9.300608e-07, 9.300609e-07, 9.300609e-07, 
    9.300607e-07, 9.300608e-07, 9.300606e-07, 9.300607e-07, 9.300605e-07, 
    9.300607e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 
    9.300604e-07, 9.300605e-07, 9.300604e-07, 9.300604e-07, 9.300604e-07, 
    9.300605e-07, 9.300608e-07, 9.300607e-07, 9.300608e-07, 9.300608e-07, 
    9.300608e-07, 9.300608e-07, 9.300609e-07, 9.300609e-07, 9.300609e-07, 
    9.300609e-07, 9.300608e-07, 9.300608e-07, 9.300607e-07, 9.300608e-07, 
    9.300607e-07, 9.300607e-07, 9.300605e-07, 9.300606e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300607e-07, 9.300607e-07, 9.300608e-07, 
    9.300608e-07, 9.300609e-07, 9.300609e-07, 9.300609e-07, 9.300609e-07, 
    9.300609e-07, 9.300608e-07, 9.300608e-07, 9.300608e-07, 9.300608e-07, 
    9.300607e-07, 9.300607e-07, 9.300605e-07, 9.300606e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 
    9.300605e-07, 9.300606e-07, 9.300605e-07, 9.300607e-07, 9.300608e-07, 
    9.300608e-07, 9.300609e-07, 9.300609e-07, 9.300609e-07, 9.300609e-07, 
    9.300609e-07, 9.300608e-07, 9.300608e-07, 9.300608e-07, 9.300608e-07, 
    9.300607e-07, 9.300607e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300604e-07, 
    9.300605e-07, 9.300604e-07, 9.300605e-07, 9.300605e-07, 9.300608e-07, 
    9.300608e-07, 9.300608e-07, 9.300609e-07, 9.300609e-07, 9.300609e-07, 
    9.300609e-07, 9.300609e-07, 9.300608e-07, 9.300608e-07, 9.300608e-07, 
    9.300607e-07, 9.300607e-07, 9.300606e-07, 9.300605e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300604e-07, 
    9.300605e-07, 9.300604e-07, 9.300604e-07, 9.300605e-07, 9.300604e-07, 
    9.300608e-07, 9.300608e-07, 9.300609e-07, 9.300609e-07, 9.300609e-07, 
    9.300609e-07, 9.300609e-07, 9.300608e-07, 9.300608e-07, 9.300608e-07, 
    9.300607e-07, 9.300607e-07, 9.300607e-07, 9.300606e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300604e-07, 9.300604e-07, 9.300604e-07, 
    9.300604e-07, 9.300608e-07, 9.300608e-07, 9.300608e-07, 9.300608e-07, 
    9.300608e-07, 9.300608e-07, 9.300608e-07, 9.300607e-07, 9.300607e-07, 
    9.300607e-07, 9.300607e-07, 9.300607e-07, 9.300607e-07, 9.300607e-07, 
    9.300606e-07, 9.300607e-07, 9.300605e-07, 9.300606e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300604e-07, 9.300604e-07, 
    9.300604e-07, 9.300604e-07, 9.300608e-07, 9.300608e-07, 9.300608e-07, 
    9.300608e-07, 9.300607e-07, 9.300607e-07, 9.300606e-07, 9.300607e-07, 
    9.300606e-07, 9.300606e-07, 9.300607e-07, 9.300606e-07, 9.300608e-07, 
    9.300607e-07, 9.300608e-07, 9.300608e-07, 9.300607e-07, 9.300607e-07, 
    9.300605e-07, 9.300606e-07, 9.300605e-07, 9.300605e-07, 9.300604e-07, 
    9.300604e-07, 9.300603e-07, 9.300603e-07, 9.300608e-07, 9.300608e-07, 
    9.300608e-07, 9.300607e-07, 9.300607e-07, 9.300606e-07, 9.300606e-07, 
    9.300606e-07, 9.300605e-07, 9.300605e-07, 9.300606e-07, 9.300605e-07, 
    9.300607e-07, 9.300607e-07, 9.300608e-07, 9.300607e-07, 9.300607e-07, 
    9.300607e-07, 9.300607e-07, 9.300606e-07, 9.300605e-07, 9.300606e-07, 
    9.300604e-07, 9.300605e-07, 9.300602e-07, 9.300603e-07, 9.300608e-07, 
    9.300608e-07, 9.300607e-07, 9.300607e-07, 9.300606e-07, 9.300606e-07, 
    9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 
    9.300605e-07, 9.300606e-07, 9.300605e-07, 9.300607e-07, 9.300607e-07, 
    9.300607e-07, 9.300607e-07, 9.300607e-07, 9.300606e-07, 9.300606e-07, 
    9.300605e-07, 9.300605e-07, 9.300606e-07, 9.300604e-07, 9.300605e-07, 
    9.300607e-07, 9.300607e-07, 9.300607e-07, 9.300607e-07, 9.300606e-07, 
    9.300606e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300606e-07, 9.300607e-07, 
    9.300607e-07, 9.300607e-07, 9.300607e-07, 9.300606e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300606e-07, 9.300605e-07, 9.300606e-07, 
    9.300605e-07, 9.300607e-07, 9.300605e-07, 9.300607e-07, 9.300607e-07, 
    9.300606e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 
    9.300606e-07, 9.300606e-07, 9.300606e-07, 9.300607e-07, 9.300607e-07, 
    9.300607e-07, 9.300607e-07, 9.300607e-07, 9.300606e-07, 9.300605e-07, 
    9.300605e-07, 9.300605e-07, 9.300604e-07, 9.300604e-07, 9.300604e-07, 
    9.300604e-07, 9.300603e-07, 9.300605e-07, 9.300604e-07, 9.300606e-07, 
    9.300606e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 9.300605e-07, 
    9.300606e-07, 9.300607e-07, 9.300607e-07, 9.300607e-07, 9.300607e-07, 
    9.300607e-07, 9.300607e-07, 9.300607e-07, 9.300606e-07, 9.300606e-07, 
    9.300605e-07, 9.300605e-07, 9.300604e-07, 9.300603e-07, 9.300603e-07, 
    9.300602e-07, 9.300602e-07, 9.300602e-07 ;

 CWDC_HR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC_LOSS =
  6.323393e-16, 6.340528e-16, 6.337199e-16, 6.351007e-16, 6.343351e-16, 
    6.352389e-16, 6.32687e-16, 6.341205e-16, 6.332057e-16, 6.324939e-16, 
    6.377764e-16, 6.351623e-16, 6.404895e-16, 6.388253e-16, 6.43003e-16, 
    6.402303e-16, 6.435617e-16, 6.429236e-16, 6.448445e-16, 6.442945e-16, 
    6.467478e-16, 6.450983e-16, 6.480189e-16, 6.463543e-16, 6.466146e-16, 
    6.450438e-16, 6.356892e-16, 6.374509e-16, 6.355847e-16, 6.358361e-16, 
    6.357234e-16, 6.343507e-16, 6.336582e-16, 6.322086e-16, 6.324719e-16, 
    6.335368e-16, 6.359491e-16, 6.35131e-16, 6.371931e-16, 6.371466e-16, 
    6.39439e-16, 6.384058e-16, 6.422541e-16, 6.411616e-16, 6.443175e-16, 
    6.435242e-16, 6.442801e-16, 6.44051e-16, 6.442831e-16, 6.431196e-16, 
    6.436182e-16, 6.425941e-16, 6.385993e-16, 6.397743e-16, 6.36267e-16, 
    6.341536e-16, 6.327498e-16, 6.317525e-16, 6.318936e-16, 6.321623e-16, 
    6.33543e-16, 6.348407e-16, 6.358287e-16, 6.364892e-16, 6.371399e-16, 
    6.391064e-16, 6.401474e-16, 6.424746e-16, 6.420553e-16, 6.42766e-16, 
    6.434453e-16, 6.445846e-16, 6.443971e-16, 6.448988e-16, 6.427476e-16, 
    6.441774e-16, 6.418163e-16, 6.424624e-16, 6.373149e-16, 6.353518e-16, 
    6.345151e-16, 6.337838e-16, 6.320019e-16, 6.332326e-16, 6.327475e-16, 
    6.339017e-16, 6.346344e-16, 6.342721e-16, 6.365073e-16, 6.356386e-16, 
    6.40209e-16, 6.38242e-16, 6.433661e-16, 6.421414e-16, 6.436595e-16, 
    6.428851e-16, 6.442116e-16, 6.430179e-16, 6.450856e-16, 6.455352e-16, 
    6.452279e-16, 6.464087e-16, 6.429516e-16, 6.442799e-16, 6.342619e-16, 
    6.34321e-16, 6.345963e-16, 6.333853e-16, 6.333113e-16, 6.322013e-16, 
    6.331892e-16, 6.336095e-16, 6.34677e-16, 6.353077e-16, 6.359071e-16, 
    6.372244e-16, 6.38694e-16, 6.407473e-16, 6.422208e-16, 6.432079e-16, 
    6.426028e-16, 6.43137e-16, 6.425398e-16, 6.422598e-16, 6.453666e-16, 
    6.436227e-16, 6.46239e-16, 6.460943e-16, 6.449106e-16, 6.461106e-16, 
    6.343625e-16, 6.340224e-16, 6.328407e-16, 6.337656e-16, 6.320804e-16, 
    6.330236e-16, 6.335656e-16, 6.356564e-16, 6.361158e-16, 6.365412e-16, 
    6.373813e-16, 6.384587e-16, 6.403468e-16, 6.419878e-16, 6.434849e-16, 
    6.433753e-16, 6.434139e-16, 6.43748e-16, 6.4292e-16, 6.438838e-16, 
    6.440454e-16, 6.436227e-16, 6.46075e-16, 6.453748e-16, 6.460913e-16, 
    6.456355e-16, 6.34133e-16, 6.347052e-16, 6.34396e-16, 6.349772e-16, 
    6.345676e-16, 6.363878e-16, 6.369331e-16, 6.394829e-16, 6.384374e-16, 
    6.401015e-16, 6.386067e-16, 6.388715e-16, 6.401549e-16, 6.386876e-16, 
    6.41897e-16, 6.397212e-16, 6.437609e-16, 6.4159e-16, 6.438969e-16, 
    6.434784e-16, 6.441713e-16, 6.447914e-16, 6.455716e-16, 6.470095e-16, 
    6.466767e-16, 6.478788e-16, 6.35558e-16, 6.362993e-16, 6.362344e-16, 
    6.370101e-16, 6.375835e-16, 6.388259e-16, 6.408163e-16, 6.400682e-16, 
    6.414416e-16, 6.417168e-16, 6.396306e-16, 6.409117e-16, 6.367955e-16, 
    6.374609e-16, 6.37065e-16, 6.356163e-16, 6.402401e-16, 6.378686e-16, 
    6.422451e-16, 6.409628e-16, 6.44703e-16, 6.428435e-16, 6.464934e-16, 
    6.480502e-16, 6.495157e-16, 6.512244e-16, 6.367041e-16, 6.362005e-16, 
    6.371024e-16, 6.383488e-16, 6.395053e-16, 6.41041e-16, 6.411982e-16, 
    6.414856e-16, 6.4223e-16, 6.428556e-16, 6.415762e-16, 6.430125e-16, 
    6.376144e-16, 6.40446e-16, 6.360098e-16, 6.373464e-16, 6.382755e-16, 
    6.378684e-16, 6.399828e-16, 6.404806e-16, 6.425015e-16, 6.414575e-16, 
    6.476658e-16, 6.449219e-16, 6.525255e-16, 6.504041e-16, 6.360244e-16, 
    6.367025e-16, 6.390598e-16, 6.379387e-16, 6.411436e-16, 6.419311e-16, 
    6.425715e-16, 6.433892e-16, 6.434777e-16, 6.43962e-16, 6.431683e-16, 
    6.439308e-16, 6.410443e-16, 6.423347e-16, 6.38791e-16, 6.396541e-16, 
    6.392572e-16, 6.388214e-16, 6.401658e-16, 6.415962e-16, 6.416274e-16, 
    6.420853e-16, 6.43375e-16, 6.411566e-16, 6.480185e-16, 6.437831e-16, 
    6.374416e-16, 6.387455e-16, 6.389324e-16, 6.384274e-16, 6.418521e-16, 
    6.406122e-16, 6.439503e-16, 6.430488e-16, 6.445257e-16, 6.437919e-16, 
    6.436839e-16, 6.42741e-16, 6.421536e-16, 6.406689e-16, 6.394598e-16, 
    6.385007e-16, 6.387238e-16, 6.397772e-16, 6.416838e-16, 6.434854e-16, 
    6.430908e-16, 6.444135e-16, 6.409115e-16, 6.423804e-16, 6.418125e-16, 
    6.432929e-16, 6.400482e-16, 6.428099e-16, 6.393413e-16, 6.396458e-16, 
    6.405875e-16, 6.424796e-16, 6.428988e-16, 6.433453e-16, 6.4307e-16, 
    6.41732e-16, 6.415132e-16, 6.405648e-16, 6.403025e-16, 6.395795e-16, 
    6.389805e-16, 6.395277e-16, 6.401021e-16, 6.417328e-16, 6.432009e-16, 
    6.448002e-16, 6.451916e-16, 6.470563e-16, 6.455377e-16, 6.48042e-16, 
    6.459119e-16, 6.495979e-16, 6.429706e-16, 6.458504e-16, 6.406306e-16, 
    6.411939e-16, 6.422114e-16, 6.445446e-16, 6.43286e-16, 6.447581e-16, 
    6.415047e-16, 6.398133e-16, 6.393761e-16, 6.385589e-16, 6.393948e-16, 
    6.393268e-16, 6.401263e-16, 6.398694e-16, 6.417869e-16, 6.407574e-16, 
    6.43681e-16, 6.447466e-16, 6.477526e-16, 6.495922e-16, 6.514634e-16, 
    6.522884e-16, 6.525395e-16, 6.526444e-16 ;

 CWDC_TO_LITR2C =
  4.805778e-16, 4.818801e-16, 4.816271e-16, 4.826765e-16, 4.820947e-16, 
    4.827816e-16, 4.808421e-16, 4.819316e-16, 4.812363e-16, 4.806954e-16, 
    4.847101e-16, 4.827234e-16, 4.86772e-16, 4.855072e-16, 4.886823e-16, 
    4.86575e-16, 4.891068e-16, 4.886219e-16, 4.900819e-16, 4.896638e-16, 
    4.915283e-16, 4.902747e-16, 4.924943e-16, 4.912293e-16, 4.914271e-16, 
    4.902333e-16, 4.831238e-16, 4.844627e-16, 4.830444e-16, 4.832354e-16, 
    4.831498e-16, 4.821065e-16, 4.815802e-16, 4.804785e-16, 4.806787e-16, 
    4.81488e-16, 4.833213e-16, 4.826996e-16, 4.842668e-16, 4.842314e-16, 
    4.859737e-16, 4.851884e-16, 4.881131e-16, 4.872828e-16, 4.896813e-16, 
    4.890784e-16, 4.896529e-16, 4.894788e-16, 4.896552e-16, 4.887709e-16, 
    4.891498e-16, 4.883716e-16, 4.853354e-16, 4.862285e-16, 4.835629e-16, 
    4.819568e-16, 4.808899e-16, 4.801319e-16, 4.802391e-16, 4.804433e-16, 
    4.814927e-16, 4.824789e-16, 4.832299e-16, 4.837318e-16, 4.842263e-16, 
    4.857208e-16, 4.86512e-16, 4.882807e-16, 4.87962e-16, 4.885022e-16, 
    4.890184e-16, 4.898843e-16, 4.897419e-16, 4.901231e-16, 4.884881e-16, 
    4.895748e-16, 4.877804e-16, 4.882714e-16, 4.843593e-16, 4.828674e-16, 
    4.822315e-16, 4.816757e-16, 4.803215e-16, 4.812568e-16, 4.808881e-16, 
    4.817653e-16, 4.823221e-16, 4.820468e-16, 4.837455e-16, 4.830853e-16, 
    4.865589e-16, 4.85064e-16, 4.889582e-16, 4.880275e-16, 4.891813e-16, 
    4.885927e-16, 4.896009e-16, 4.886936e-16, 4.902651e-16, 4.906068e-16, 
    4.903732e-16, 4.912706e-16, 4.886432e-16, 4.896528e-16, 4.82039e-16, 
    4.820839e-16, 4.822933e-16, 4.813728e-16, 4.813166e-16, 4.80473e-16, 
    4.812238e-16, 4.815433e-16, 4.823545e-16, 4.828338e-16, 4.832894e-16, 
    4.842906e-16, 4.854075e-16, 4.86968e-16, 4.880878e-16, 4.88838e-16, 
    4.883781e-16, 4.887841e-16, 4.883302e-16, 4.881175e-16, 4.904787e-16, 
    4.891533e-16, 4.911416e-16, 4.910317e-16, 4.901321e-16, 4.910441e-16, 
    4.821155e-16, 4.81857e-16, 4.809589e-16, 4.816618e-16, 4.803811e-16, 
    4.81098e-16, 4.815099e-16, 4.830988e-16, 4.83448e-16, 4.837713e-16, 
    4.844098e-16, 4.852286e-16, 4.866636e-16, 4.879107e-16, 4.890485e-16, 
    4.889652e-16, 4.889946e-16, 4.892485e-16, 4.886192e-16, 4.893517e-16, 
    4.894745e-16, 4.891533e-16, 4.91017e-16, 4.904849e-16, 4.910294e-16, 
    4.90683e-16, 4.819411e-16, 4.823759e-16, 4.821409e-16, 4.825827e-16, 
    4.822714e-16, 4.836547e-16, 4.840692e-16, 4.86007e-16, 4.852124e-16, 
    4.864771e-16, 4.853411e-16, 4.855424e-16, 4.865178e-16, 4.854026e-16, 
    4.878417e-16, 4.861881e-16, 4.892583e-16, 4.876084e-16, 4.893616e-16, 
    4.890436e-16, 4.895702e-16, 4.900415e-16, 4.906344e-16, 4.917272e-16, 
    4.914743e-16, 4.923879e-16, 4.830241e-16, 4.835875e-16, 4.835381e-16, 
    4.841277e-16, 4.845634e-16, 4.855077e-16, 4.870204e-16, 4.864518e-16, 
    4.874957e-16, 4.877047e-16, 4.861193e-16, 4.870929e-16, 4.839646e-16, 
    4.844703e-16, 4.841694e-16, 4.830683e-16, 4.865825e-16, 4.847801e-16, 
    4.881063e-16, 4.871317e-16, 4.899743e-16, 4.88561e-16, 4.91335e-16, 
    4.925182e-16, 4.936319e-16, 4.949306e-16, 4.838952e-16, 4.835124e-16, 
    4.841978e-16, 4.851451e-16, 4.86024e-16, 4.871912e-16, 4.873107e-16, 
    4.875291e-16, 4.880947e-16, 4.885702e-16, 4.875979e-16, 4.886895e-16, 
    4.84587e-16, 4.86739e-16, 4.833674e-16, 4.843833e-16, 4.850894e-16, 
    4.847799e-16, 4.863869e-16, 4.867653e-16, 4.883012e-16, 4.875077e-16, 
    4.92226e-16, 4.901406e-16, 4.959194e-16, 4.943071e-16, 4.833786e-16, 
    4.838939e-16, 4.856855e-16, 4.848334e-16, 4.872692e-16, 4.878676e-16, 
    4.883543e-16, 4.889758e-16, 4.89043e-16, 4.894111e-16, 4.888079e-16, 
    4.893874e-16, 4.871937e-16, 4.881744e-16, 4.854811e-16, 4.861371e-16, 
    4.858354e-16, 4.855043e-16, 4.86526e-16, 4.876132e-16, 4.876368e-16, 
    4.879848e-16, 4.88965e-16, 4.87279e-16, 4.924941e-16, 4.892751e-16, 
    4.844556e-16, 4.854466e-16, 4.855886e-16, 4.852048e-16, 4.878076e-16, 
    4.868652e-16, 4.894022e-16, 4.887171e-16, 4.898395e-16, 4.892819e-16, 
    4.891998e-16, 4.884832e-16, 4.880367e-16, 4.869084e-16, 4.859894e-16, 
    4.852605e-16, 4.854301e-16, 4.862307e-16, 4.876797e-16, 4.890489e-16, 
    4.88749e-16, 4.897543e-16, 4.870927e-16, 4.882091e-16, 4.877775e-16, 
    4.889027e-16, 4.864366e-16, 4.885355e-16, 4.858993e-16, 4.861308e-16, 
    4.868465e-16, 4.882845e-16, 4.886031e-16, 4.889424e-16, 4.887331e-16, 
    4.877163e-16, 4.8755e-16, 4.868292e-16, 4.8663e-16, 4.860804e-16, 
    4.856252e-16, 4.860411e-16, 4.864775e-16, 4.877169e-16, 4.888327e-16, 
    4.900482e-16, 4.903456e-16, 4.917627e-16, 4.906086e-16, 4.925119e-16, 
    4.90893e-16, 4.936944e-16, 4.886577e-16, 4.908463e-16, 4.868792e-16, 
    4.873074e-16, 4.880807e-16, 4.898539e-16, 4.888974e-16, 4.900161e-16, 
    4.875436e-16, 4.862581e-16, 4.859258e-16, 4.853048e-16, 4.8594e-16, 
    4.858884e-16, 4.86496e-16, 4.863008e-16, 4.87758e-16, 4.869756e-16, 
    4.891976e-16, 4.900074e-16, 4.92292e-16, 4.9369e-16, 4.951121e-16, 
    4.957392e-16, 4.9593e-16, 4.960097e-16 ;

 CWDC_TO_LITR3C =
  1.517614e-16, 1.521727e-16, 1.520928e-16, 1.524242e-16, 1.522404e-16, 
    1.524573e-16, 1.518449e-16, 1.521889e-16, 1.519694e-16, 1.517985e-16, 
    1.530663e-16, 1.52439e-16, 1.537175e-16, 1.533181e-16, 1.543207e-16, 
    1.536553e-16, 1.544548e-16, 1.543017e-16, 1.547627e-16, 1.546307e-16, 
    1.552195e-16, 1.548236e-16, 1.555245e-16, 1.55125e-16, 1.551875e-16, 
    1.548105e-16, 1.525654e-16, 1.529882e-16, 1.525403e-16, 1.526007e-16, 
    1.525736e-16, 1.522442e-16, 1.52078e-16, 1.517301e-16, 1.517933e-16, 
    1.520488e-16, 1.526278e-16, 1.524314e-16, 1.529264e-16, 1.529152e-16, 
    1.534654e-16, 1.532174e-16, 1.54141e-16, 1.538788e-16, 1.546362e-16, 
    1.544458e-16, 1.546272e-16, 1.545722e-16, 1.546279e-16, 1.543487e-16, 
    1.544684e-16, 1.542226e-16, 1.532638e-16, 1.535458e-16, 1.527041e-16, 
    1.521969e-16, 1.5186e-16, 1.516206e-16, 1.516545e-16, 1.517189e-16, 
    1.520503e-16, 1.523618e-16, 1.525989e-16, 1.527574e-16, 1.529136e-16, 
    1.533855e-16, 1.536354e-16, 1.541939e-16, 1.540933e-16, 1.542638e-16, 
    1.544269e-16, 1.547003e-16, 1.546553e-16, 1.547757e-16, 1.542594e-16, 
    1.546026e-16, 1.540359e-16, 1.54191e-16, 1.529556e-16, 1.524844e-16, 
    1.522836e-16, 1.521081e-16, 1.516805e-16, 1.519758e-16, 1.518594e-16, 
    1.521364e-16, 1.523122e-16, 1.522253e-16, 1.527618e-16, 1.525533e-16, 
    1.536502e-16, 1.531781e-16, 1.544079e-16, 1.541139e-16, 1.544783e-16, 
    1.542924e-16, 1.546108e-16, 1.543243e-16, 1.548205e-16, 1.549285e-16, 
    1.548547e-16, 1.551381e-16, 1.543084e-16, 1.546272e-16, 1.522228e-16, 
    1.52237e-16, 1.523031e-16, 1.520125e-16, 1.519947e-16, 1.517283e-16, 
    1.519654e-16, 1.520663e-16, 1.523225e-16, 1.524738e-16, 1.526177e-16, 
    1.529339e-16, 1.532866e-16, 1.537794e-16, 1.54133e-16, 1.543699e-16, 
    1.542247e-16, 1.543529e-16, 1.542095e-16, 1.541424e-16, 1.54888e-16, 
    1.544694e-16, 1.550973e-16, 1.550626e-16, 1.547785e-16, 1.550666e-16, 
    1.52247e-16, 1.521654e-16, 1.518818e-16, 1.521037e-16, 1.516993e-16, 
    1.519257e-16, 1.520558e-16, 1.525575e-16, 1.526678e-16, 1.527699e-16, 
    1.529715e-16, 1.532301e-16, 1.536832e-16, 1.540771e-16, 1.544364e-16, 
    1.544101e-16, 1.544193e-16, 1.544995e-16, 1.543008e-16, 1.545321e-16, 
    1.545709e-16, 1.544695e-16, 1.55058e-16, 1.5489e-16, 1.550619e-16, 
    1.549525e-16, 1.521919e-16, 1.523292e-16, 1.52255e-16, 1.523945e-16, 
    1.522962e-16, 1.527331e-16, 1.528639e-16, 1.534759e-16, 1.53225e-16, 
    1.536244e-16, 1.532656e-16, 1.533292e-16, 1.536372e-16, 1.53285e-16, 
    1.540553e-16, 1.535331e-16, 1.545026e-16, 1.539816e-16, 1.545352e-16, 
    1.544348e-16, 1.546011e-16, 1.547499e-16, 1.549372e-16, 1.552823e-16, 
    1.552024e-16, 1.554909e-16, 1.525339e-16, 1.527118e-16, 1.526963e-16, 
    1.528824e-16, 1.5302e-16, 1.533182e-16, 1.537959e-16, 1.536164e-16, 
    1.53946e-16, 1.54012e-16, 1.535114e-16, 1.538188e-16, 1.528309e-16, 
    1.529906e-16, 1.528956e-16, 1.525479e-16, 1.536576e-16, 1.530885e-16, 
    1.541388e-16, 1.538311e-16, 1.547287e-16, 1.542824e-16, 1.551584e-16, 
    1.555321e-16, 1.558838e-16, 1.562939e-16, 1.52809e-16, 1.526881e-16, 
    1.529046e-16, 1.532037e-16, 1.534813e-16, 1.538498e-16, 1.538876e-16, 
    1.539565e-16, 1.541352e-16, 1.542853e-16, 1.539783e-16, 1.54323e-16, 
    1.530275e-16, 1.53707e-16, 1.526423e-16, 1.529631e-16, 1.531861e-16, 
    1.530884e-16, 1.535959e-16, 1.537153e-16, 1.542004e-16, 1.539498e-16, 
    1.554398e-16, 1.547813e-16, 1.566061e-16, 1.56097e-16, 1.526459e-16, 
    1.528086e-16, 1.533743e-16, 1.531053e-16, 1.538745e-16, 1.540635e-16, 
    1.542172e-16, 1.544134e-16, 1.544346e-16, 1.545509e-16, 1.543604e-16, 
    1.545434e-16, 1.538506e-16, 1.541603e-16, 1.533098e-16, 1.53517e-16, 
    1.534217e-16, 1.533171e-16, 1.536398e-16, 1.539831e-16, 1.539906e-16, 
    1.541005e-16, 1.5441e-16, 1.538776e-16, 1.555244e-16, 1.545079e-16, 
    1.52986e-16, 1.532989e-16, 1.533438e-16, 1.532226e-16, 1.540445e-16, 
    1.537469e-16, 1.545481e-16, 1.543317e-16, 1.546862e-16, 1.545101e-16, 
    1.544841e-16, 1.542579e-16, 1.541169e-16, 1.537605e-16, 1.534704e-16, 
    1.532402e-16, 1.532937e-16, 1.535465e-16, 1.540041e-16, 1.544365e-16, 
    1.543418e-16, 1.546592e-16, 1.538187e-16, 1.541713e-16, 1.54035e-16, 
    1.543903e-16, 1.536116e-16, 1.542744e-16, 1.534419e-16, 1.53515e-16, 
    1.53741e-16, 1.541951e-16, 1.542957e-16, 1.544029e-16, 1.543368e-16, 
    1.540157e-16, 1.539632e-16, 1.537356e-16, 1.536726e-16, 1.534991e-16, 
    1.533553e-16, 1.534866e-16, 1.536245e-16, 1.540159e-16, 1.543682e-16, 
    1.54752e-16, 1.54846e-16, 1.552935e-16, 1.54929e-16, 1.555301e-16, 
    1.550188e-16, 1.559035e-16, 1.54313e-16, 1.550041e-16, 1.537513e-16, 
    1.538865e-16, 1.541307e-16, 1.546907e-16, 1.543886e-16, 1.547419e-16, 
    1.539611e-16, 1.535552e-16, 1.534503e-16, 1.532541e-16, 1.534547e-16, 
    1.534384e-16, 1.536303e-16, 1.535687e-16, 1.540289e-16, 1.537818e-16, 
    1.544834e-16, 1.547392e-16, 1.554606e-16, 1.559021e-16, 1.563512e-16, 
    1.565492e-16, 1.566095e-16, 1.566347e-16 ;

 CWDC_vr =
  5.310744e-05, 5.310744e-05, 5.310744e-05, 5.310743e-05, 5.310744e-05, 
    5.310743e-05, 5.310744e-05, 5.310744e-05, 5.310744e-05, 5.310744e-05, 
    5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310743e-05, 5.310742e-05, 
    5.310742e-05, 5.310741e-05, 5.310742e-05, 5.310741e-05, 5.310741e-05, 
    5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310741e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310744e-05, 5.310744e-05, 5.310744e-05, 5.310744e-05, 
    5.310744e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310742e-05, 5.310741e-05, 
    5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310742e-05, 
    5.310741e-05, 5.310742e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310744e-05, 5.310744e-05, 5.310744e-05, 5.310744e-05, 5.310744e-05, 
    5.310744e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 
    5.310742e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310742e-05, 
    5.310741e-05, 5.310742e-05, 5.310742e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310744e-05, 5.310744e-05, 5.310744e-05, 5.310744e-05, 
    5.310744e-05, 5.310743e-05, 5.310744e-05, 5.310743e-05, 5.310743e-05, 
    5.310742e-05, 5.310743e-05, 5.310742e-05, 5.310742e-05, 5.310741e-05, 
    5.310742e-05, 5.310741e-05, 5.310742e-05, 5.310741e-05, 5.310741e-05, 
    5.310741e-05, 5.310741e-05, 5.310742e-05, 5.310741e-05, 5.310744e-05, 
    5.310744e-05, 5.310743e-05, 5.310744e-05, 5.310744e-05, 5.310744e-05, 
    5.310744e-05, 5.310744e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 
    5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310741e-05, 
    5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310744e-05, 5.310744e-05, 5.310744e-05, 5.310744e-05, 5.310744e-05, 
    5.310744e-05, 5.310744e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 
    5.310742e-05, 5.310742e-05, 5.310741e-05, 5.310742e-05, 5.310741e-05, 
    5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310741e-05, 5.310744e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310742e-05, 5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310743e-05, 
    5.310742e-05, 5.310743e-05, 5.310741e-05, 5.310742e-05, 5.310741e-05, 
    5.310742e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310741e-05, 5.310741e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310742e-05, 
    5.310742e-05, 5.310742e-05, 5.310743e-05, 5.310742e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310743e-05, 
    5.310742e-05, 5.310742e-05, 5.310741e-05, 5.310742e-05, 5.310741e-05, 
    5.310741e-05, 5.31074e-05, 5.31074e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310742e-05, 
    5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 
    5.310743e-05, 5.310742e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 
    5.310741e-05, 5.310741e-05, 5.31074e-05, 5.31074e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310742e-05, 
    5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310741e-05, 5.310742e-05, 
    5.310741e-05, 5.310742e-05, 5.310742e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 
    5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310741e-05, 5.310741e-05, 
    5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310742e-05, 
    5.310742e-05, 5.310741e-05, 5.310742e-05, 5.310741e-05, 5.310741e-05, 
    5.310741e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310742e-05, 
    5.310742e-05, 5.310741e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 
    5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310743e-05, 5.310743e-05, 
    5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 
    5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310743e-05, 
    5.310743e-05, 5.310743e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 
    5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 5.310741e-05, 
    5.310741e-05, 5.31074e-05, 5.310742e-05, 5.310741e-05, 5.310742e-05, 
    5.310742e-05, 5.310742e-05, 5.310741e-05, 5.310742e-05, 5.310741e-05, 
    5.310742e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 5.310743e-05, 
    5.310743e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 5.310742e-05, 
    5.310741e-05, 5.310741e-05, 5.310741e-05, 5.31074e-05, 5.31074e-05, 
    5.31074e-05, 5.31074e-05, 5.31074e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDN =
  1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860121e-09, 1.860122e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860122e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860122e-09, 
    1.860122e-09, 1.860122e-09, 1.860122e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860122e-09, 1.860122e-09, 
    1.860122e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860122e-09, 1.860122e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.86012e-09, 1.860121e-09, 1.860122e-09, 
    1.860122e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860122e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 1.860121e-09, 
    1.86012e-09, 1.86012e-09, 1.86012e-09 ;

 CWDN_TO_LITR2N =
  9.611556e-19, 9.637602e-19, 9.632543e-19, 9.653531e-19, 9.641893e-19, 
    9.655631e-19, 9.616843e-19, 9.638632e-19, 9.624726e-19, 9.613908e-19, 
    9.694201e-19, 9.654467e-19, 9.73544e-19, 9.710144e-19, 9.773646e-19, 
    9.731501e-19, 9.782137e-19, 9.772439e-19, 9.801637e-19, 9.793277e-19, 
    9.830566e-19, 9.805495e-19, 9.849887e-19, 9.824585e-19, 9.828542e-19, 
    9.804666e-19, 9.662477e-19, 9.689255e-19, 9.660887e-19, 9.664708e-19, 
    9.662996e-19, 9.642131e-19, 9.631604e-19, 9.60957e-19, 9.613574e-19, 
    9.62976e-19, 9.666426e-19, 9.653991e-19, 9.685336e-19, 9.684629e-19, 
    9.719474e-19, 9.703768e-19, 9.762262e-19, 9.745657e-19, 9.793626e-19, 
    9.781568e-19, 9.793057e-19, 9.789576e-19, 9.793103e-19, 9.775418e-19, 
    9.782996e-19, 9.76743e-19, 9.706709e-19, 9.724569e-19, 9.671258e-19, 
    9.639135e-19, 9.617798e-19, 9.602638e-19, 9.604783e-19, 9.608866e-19, 
    9.629854e-19, 9.649578e-19, 9.664596e-19, 9.674637e-19, 9.684526e-19, 
    9.714416e-19, 9.73024e-19, 9.765615e-19, 9.75924e-19, 9.770043e-19, 
    9.780368e-19, 9.797686e-19, 9.794837e-19, 9.802461e-19, 9.769763e-19, 
    9.791497e-19, 9.755607e-19, 9.765428e-19, 9.687187e-19, 9.657348e-19, 
    9.64463e-19, 9.633514e-19, 9.60643e-19, 9.625136e-19, 9.617762e-19, 
    9.635306e-19, 9.646443e-19, 9.640936e-19, 9.674911e-19, 9.661707e-19, 
    9.731177e-19, 9.701279e-19, 9.779165e-19, 9.760549e-19, 9.783626e-19, 
    9.771855e-19, 9.792017e-19, 9.773872e-19, 9.805301e-19, 9.812135e-19, 
    9.807465e-19, 9.825413e-19, 9.772865e-19, 9.793055e-19, 9.640781e-19, 
    9.641678e-19, 9.645865e-19, 9.627457e-19, 9.626332e-19, 9.60946e-19, 
    9.624476e-19, 9.630865e-19, 9.64709e-19, 9.656677e-19, 9.665788e-19, 
    9.685811e-19, 9.708149e-19, 9.739359e-19, 9.761756e-19, 9.77676e-19, 
    9.767563e-19, 9.775683e-19, 9.766604e-19, 9.762349e-19, 9.809573e-19, 
    9.783065e-19, 9.822832e-19, 9.820635e-19, 9.802641e-19, 9.820882e-19, 
    9.642309e-19, 9.63714e-19, 9.619178e-19, 9.633237e-19, 9.607621e-19, 
    9.621959e-19, 9.630198e-19, 9.661977e-19, 9.668961e-19, 9.675426e-19, 
    9.688197e-19, 9.704573e-19, 9.733271e-19, 9.758215e-19, 9.78097e-19, 
    9.779305e-19, 9.779891e-19, 9.784969e-19, 9.772384e-19, 9.787035e-19, 
    9.789489e-19, 9.783065e-19, 9.82034e-19, 9.809697e-19, 9.820587e-19, 
    9.813659e-19, 9.638821e-19, 9.647519e-19, 9.642819e-19, 9.651654e-19, 
    9.645427e-19, 9.673095e-19, 9.681383e-19, 9.72014e-19, 9.704248e-19, 
    9.729542e-19, 9.706822e-19, 9.710847e-19, 9.730355e-19, 9.708051e-19, 
    9.756834e-19, 9.723762e-19, 9.785166e-19, 9.752168e-19, 9.787232e-19, 
    9.780872e-19, 9.791404e-19, 9.80083e-19, 9.812687e-19, 9.834544e-19, 
    9.829485e-19, 9.847757e-19, 9.660481e-19, 9.671749e-19, 9.670763e-19, 
    9.682553e-19, 9.691269e-19, 9.710154e-19, 9.740407e-19, 9.729037e-19, 
    9.749913e-19, 9.754095e-19, 9.722385e-19, 9.741857e-19, 9.679291e-19, 
    9.689406e-19, 9.683388e-19, 9.661367e-19, 9.731651e-19, 9.695603e-19, 
    9.762125e-19, 9.742635e-19, 9.799486e-19, 9.771221e-19, 9.8267e-19, 
    9.850363e-19, 9.872637e-19, 9.898612e-19, 9.677903e-19, 9.670248e-19, 
    9.683956e-19, 9.702901e-19, 9.720481e-19, 9.743824e-19, 9.746213e-19, 
    9.750582e-19, 9.761895e-19, 9.771405e-19, 9.751958e-19, 9.773789e-19, 
    9.691739e-19, 9.734779e-19, 9.667349e-19, 9.687665e-19, 9.701787e-19, 
    9.695599e-19, 9.727738e-19, 9.735305e-19, 9.766023e-19, 9.750154e-19, 
    9.84452e-19, 9.802813e-19, 9.918388e-19, 9.886143e-19, 9.667572e-19, 
    9.677879e-19, 9.713709e-19, 9.696668e-19, 9.745384e-19, 9.757352e-19, 
    9.767086e-19, 9.779515e-19, 9.780861e-19, 9.788223e-19, 9.776157e-19, 
    9.787748e-19, 9.743872e-19, 9.763488e-19, 9.709623e-19, 9.722742e-19, 
    9.716709e-19, 9.710086e-19, 9.730521e-19, 9.752263e-19, 9.752735e-19, 
    9.759696e-19, 9.7793e-19, 9.74558e-19, 9.849882e-19, 9.785503e-19, 
    9.689113e-19, 9.708932e-19, 9.711772e-19, 9.704096e-19, 9.756152e-19, 
    9.737304e-19, 9.788044e-19, 9.774341e-19, 9.796791e-19, 9.785638e-19, 
    9.783996e-19, 9.769664e-19, 9.760735e-19, 9.738168e-19, 9.719789e-19, 
    9.70521e-19, 9.708601e-19, 9.724614e-19, 9.753594e-19, 9.780979e-19, 
    9.77498e-19, 9.795086e-19, 9.741854e-19, 9.764182e-19, 9.75555e-19, 
    9.778052e-19, 9.728733e-19, 9.770711e-19, 9.717987e-19, 9.722616e-19, 
    9.73693e-19, 9.76569e-19, 9.772062e-19, 9.778849e-19, 9.774663e-19, 
    9.754326e-19, 9.751002e-19, 9.736585e-19, 9.732599e-19, 9.721609e-19, 
    9.712503e-19, 9.720821e-19, 9.729552e-19, 9.754338e-19, 9.776653e-19, 
    9.800963e-19, 9.806912e-19, 9.835255e-19, 9.812173e-19, 9.850238e-19, 
    9.81786e-19, 9.873889e-19, 9.773153e-19, 9.816926e-19, 9.737585e-19, 
    9.746147e-19, 9.761613e-19, 9.797078e-19, 9.777947e-19, 9.800323e-19, 
    9.750871e-19, 9.725162e-19, 9.718516e-19, 9.706095e-19, 9.7188e-19, 
    9.717767e-19, 9.729919e-19, 9.726015e-19, 9.75516e-19, 9.739512e-19, 
    9.783952e-19, 9.800148e-19, 9.84584e-19, 9.873801e-19, 9.902243e-19, 
    9.914783e-19, 9.9186e-19, 9.920195e-19 ;

 CWDN_TO_LITR3N =
  3.035228e-19, 3.043453e-19, 3.041856e-19, 3.048483e-19, 3.044808e-19, 
    3.049147e-19, 3.036898e-19, 3.043779e-19, 3.039387e-19, 3.035971e-19, 
    3.061327e-19, 3.048779e-19, 3.07435e-19, 3.066361e-19, 3.086414e-19, 
    3.073105e-19, 3.089096e-19, 3.086033e-19, 3.095254e-19, 3.092614e-19, 
    3.104389e-19, 3.096472e-19, 3.110491e-19, 3.102501e-19, 3.10375e-19, 
    3.09621e-19, 3.051308e-19, 3.059765e-19, 3.050807e-19, 3.052013e-19, 
    3.051472e-19, 3.044883e-19, 3.041559e-19, 3.034601e-19, 3.035865e-19, 
    3.040977e-19, 3.052556e-19, 3.048629e-19, 3.058527e-19, 3.058304e-19, 
    3.069307e-19, 3.064348e-19, 3.082819e-19, 3.077576e-19, 3.092724e-19, 
    3.088916e-19, 3.092544e-19, 3.091445e-19, 3.092559e-19, 3.086974e-19, 
    3.089367e-19, 3.084452e-19, 3.065276e-19, 3.070917e-19, 3.054081e-19, 
    3.043937e-19, 3.037199e-19, 3.032412e-19, 3.033089e-19, 3.034379e-19, 
    3.041006e-19, 3.047235e-19, 3.051978e-19, 3.055148e-19, 3.058272e-19, 
    3.06771e-19, 3.072707e-19, 3.083878e-19, 3.081865e-19, 3.085277e-19, 
    3.088538e-19, 3.094006e-19, 3.093106e-19, 3.095514e-19, 3.085188e-19, 
    3.092052e-19, 3.080718e-19, 3.083819e-19, 3.059111e-19, 3.049689e-19, 
    3.045673e-19, 3.042162e-19, 3.033609e-19, 3.039517e-19, 3.037188e-19, 
    3.042728e-19, 3.046245e-19, 3.044506e-19, 3.055235e-19, 3.051065e-19, 
    3.073003e-19, 3.063562e-19, 3.088157e-19, 3.082279e-19, 3.089566e-19, 
    3.085849e-19, 3.092216e-19, 3.086486e-19, 3.096411e-19, 3.098569e-19, 
    3.097094e-19, 3.102762e-19, 3.086168e-19, 3.092544e-19, 3.044457e-19, 
    3.04474e-19, 3.046063e-19, 3.04025e-19, 3.039894e-19, 3.034566e-19, 
    3.039308e-19, 3.041326e-19, 3.04645e-19, 3.049477e-19, 3.052354e-19, 
    3.058677e-19, 3.065731e-19, 3.075587e-19, 3.08266e-19, 3.087398e-19, 
    3.084493e-19, 3.087058e-19, 3.084191e-19, 3.082847e-19, 3.09776e-19, 
    3.089389e-19, 3.101947e-19, 3.101253e-19, 3.095571e-19, 3.101331e-19, 
    3.04494e-19, 3.043308e-19, 3.037635e-19, 3.042075e-19, 3.033986e-19, 
    3.038514e-19, 3.041115e-19, 3.051151e-19, 3.053356e-19, 3.055398e-19, 
    3.05943e-19, 3.064602e-19, 3.073665e-19, 3.081541e-19, 3.088728e-19, 
    3.088202e-19, 3.088387e-19, 3.08999e-19, 3.086016e-19, 3.090642e-19, 
    3.091418e-19, 3.089389e-19, 3.10116e-19, 3.097799e-19, 3.101238e-19, 
    3.09905e-19, 3.043838e-19, 3.046585e-19, 3.045101e-19, 3.047891e-19, 
    3.045925e-19, 3.054661e-19, 3.057279e-19, 3.069518e-19, 3.064499e-19, 
    3.072487e-19, 3.065312e-19, 3.066583e-19, 3.072744e-19, 3.065701e-19, 
    3.081105e-19, 3.070662e-19, 3.090053e-19, 3.079632e-19, 3.090705e-19, 
    3.088697e-19, 3.092022e-19, 3.094999e-19, 3.098743e-19, 3.105645e-19, 
    3.104048e-19, 3.109818e-19, 3.050678e-19, 3.054237e-19, 3.053925e-19, 
    3.057648e-19, 3.060401e-19, 3.066364e-19, 3.075918e-19, 3.072327e-19, 
    3.07892e-19, 3.08024e-19, 3.070227e-19, 3.076376e-19, 3.056618e-19, 
    3.059812e-19, 3.057912e-19, 3.050958e-19, 3.073153e-19, 3.061769e-19, 
    3.082777e-19, 3.076622e-19, 3.094574e-19, 3.085649e-19, 3.103168e-19, 
    3.110641e-19, 3.117675e-19, 3.125877e-19, 3.05618e-19, 3.053763e-19, 
    3.058092e-19, 3.064074e-19, 3.069625e-19, 3.076997e-19, 3.077752e-19, 
    3.079131e-19, 3.082704e-19, 3.085707e-19, 3.079566e-19, 3.08646e-19, 
    3.060549e-19, 3.074141e-19, 3.052847e-19, 3.059263e-19, 3.063722e-19, 
    3.061768e-19, 3.071917e-19, 3.074307e-19, 3.084007e-19, 3.078996e-19, 
    3.108796e-19, 3.095625e-19, 3.132122e-19, 3.12194e-19, 3.052917e-19, 
    3.056172e-19, 3.067487e-19, 3.062106e-19, 3.07749e-19, 3.081269e-19, 
    3.084343e-19, 3.088268e-19, 3.088693e-19, 3.091018e-19, 3.087208e-19, 
    3.090868e-19, 3.077012e-19, 3.083206e-19, 3.066197e-19, 3.07034e-19, 
    3.068434e-19, 3.066343e-19, 3.072796e-19, 3.079662e-19, 3.079811e-19, 
    3.082009e-19, 3.0882e-19, 3.077552e-19, 3.110489e-19, 3.090159e-19, 
    3.05972e-19, 3.065979e-19, 3.066876e-19, 3.064451e-19, 3.08089e-19, 
    3.074938e-19, 3.090961e-19, 3.086634e-19, 3.093723e-19, 3.090201e-19, 
    3.089683e-19, 3.085157e-19, 3.082337e-19, 3.075211e-19, 3.069407e-19, 
    3.064803e-19, 3.065874e-19, 3.070931e-19, 3.080082e-19, 3.08873e-19, 
    3.086836e-19, 3.093185e-19, 3.076375e-19, 3.083426e-19, 3.0807e-19, 
    3.087806e-19, 3.072231e-19, 3.085488e-19, 3.068838e-19, 3.0703e-19, 
    3.07482e-19, 3.083902e-19, 3.085914e-19, 3.088057e-19, 3.086736e-19, 
    3.080313e-19, 3.079264e-19, 3.074711e-19, 3.073452e-19, 3.069982e-19, 
    3.067106e-19, 3.069733e-19, 3.07249e-19, 3.080317e-19, 3.087364e-19, 
    3.095041e-19, 3.096919e-19, 3.10587e-19, 3.098581e-19, 3.110602e-19, 
    3.100377e-19, 3.11807e-19, 3.086259e-19, 3.100082e-19, 3.075027e-19, 
    3.077731e-19, 3.082614e-19, 3.093814e-19, 3.087773e-19, 3.094839e-19, 
    3.079222e-19, 3.071104e-19, 3.069005e-19, 3.065083e-19, 3.069095e-19, 
    3.068769e-19, 3.072606e-19, 3.071373e-19, 3.080577e-19, 3.075635e-19, 
    3.089669e-19, 3.094784e-19, 3.109212e-19, 3.118042e-19, 3.127024e-19, 
    3.130984e-19, 3.132189e-19, 3.132693e-19 ;

 CWDN_vr =
  1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062148e-07, 1.062149e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062149e-07, 1.062148e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062148e-07, 1.062149e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062148e-07, 1.062149e-07, 
    1.062148e-07, 1.062149e-07, 1.062148e-07, 1.062148e-07, 1.062149e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062149e-07, 1.062148e-07, 1.062149e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062149e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062149e-07, 1.062148e-07, 1.062149e-07, 1.062149e-07, 1.062149e-07, 
    1.062149e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062149e-07, 
    1.062149e-07, 1.062148e-07, 1.062149e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062149e-07, 1.062148e-07, 1.062148e-07, 1.062149e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062149e-07, 1.062149e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062149e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 1.062148e-07, 
    1.062148e-07, 1.062148e-07, 1.062148e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADSTEMC =
  0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504 ;

 DEADSTEMN =
  6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 6.149009e-05, 
    6.149009e-05, 6.149009e-05, 6.149009e-05 ;

 DENIT =
  1.095188e-14, 1.099342e-14, 1.09853e-14, 1.101883e-14, 1.10002e-14, 
    1.102213e-14, 1.09602e-14, 1.099496e-14, 1.097274e-14, 1.095546e-14, 
    1.108377e-14, 1.102018e-14, 1.114976e-14, 1.110917e-14, 1.121104e-14, 
    1.114341e-14, 1.122466e-14, 1.120902e-14, 1.125594e-14, 1.124247e-14, 
    1.130251e-14, 1.12621e-14, 1.133359e-14, 1.129282e-14, 1.129918e-14, 
    1.126068e-14, 1.103308e-14, 1.107599e-14, 1.103051e-14, 1.103663e-14, 
    1.103386e-14, 1.100052e-14, 1.098373e-14, 1.094853e-14, 1.095489e-14, 
    1.098072e-14, 1.103925e-14, 1.101933e-14, 1.10694e-14, 1.106828e-14, 
    1.112404e-14, 1.109888e-14, 1.119266e-14, 1.116596e-14, 1.124301e-14, 
    1.12236e-14, 1.124207e-14, 1.123643e-14, 1.124209e-14, 1.121367e-14, 
    1.12258e-14, 1.12008e-14, 1.110381e-14, 1.11324e-14, 1.104706e-14, 
    1.099576e-14, 1.096165e-14, 1.093749e-14, 1.094087e-14, 1.094739e-14, 
    1.098084e-14, 1.101227e-14, 1.103625e-14, 1.105227e-14, 1.106806e-14, 
    1.111598e-14, 1.114129e-14, 1.119802e-14, 1.118775e-14, 1.120509e-14, 
    1.122165e-14, 1.124947e-14, 1.124487e-14, 1.125712e-14, 1.120452e-14, 
    1.123947e-14, 1.118175e-14, 1.119753e-14, 1.10726e-14, 1.102478e-14, 
    1.10045e-14, 1.09867e-14, 1.094348e-14, 1.097332e-14, 1.096153e-14, 
    1.098947e-14, 1.100724e-14, 1.099842e-14, 1.105269e-14, 1.103156e-14, 
    1.114276e-14, 1.109485e-14, 1.121974e-14, 1.118981e-14, 1.122686e-14, 
    1.120794e-14, 1.124032e-14, 1.121115e-14, 1.126164e-14, 1.127266e-14, 
    1.12651e-14, 1.129398e-14, 1.120942e-14, 1.124189e-14, 1.099828e-14, 
    1.099972e-14, 1.100638e-14, 1.097699e-14, 1.097519e-14, 1.094825e-14, 
    1.097216e-14, 1.098237e-14, 1.100822e-14, 1.102351e-14, 1.103805e-14, 
    1.107007e-14, 1.110582e-14, 1.115581e-14, 1.119173e-14, 1.121579e-14, 
    1.120101e-14, 1.121403e-14, 1.119944e-14, 1.119257e-14, 1.126848e-14, 
    1.122585e-14, 1.128978e-14, 1.128624e-14, 1.125727e-14, 1.128658e-14, 
    1.100069e-14, 1.099241e-14, 1.096376e-14, 1.098615e-14, 1.094528e-14, 
    1.096815e-14, 1.098128e-14, 1.103199e-14, 1.10431e-14, 1.105345e-14, 
    1.107384e-14, 1.110003e-14, 1.114602e-14, 1.118601e-14, 1.122254e-14, 
    1.121983e-14, 1.122077e-14, 1.122891e-14, 1.120868e-14, 1.123219e-14, 
    1.123612e-14, 1.122579e-14, 1.128571e-14, 1.126858e-14, 1.128609e-14, 
    1.12749e-14, 1.099507e-14, 1.100893e-14, 1.10014e-14, 1.101552e-14, 
    1.100554e-14, 1.104976e-14, 1.1063e-14, 1.112502e-14, 1.109951e-14, 
    1.114006e-14, 1.110359e-14, 1.111005e-14, 1.114134e-14, 1.110551e-14, 
    1.118376e-14, 1.113069e-14, 1.12292e-14, 1.117622e-14, 1.123249e-14, 
    1.122223e-14, 1.123914e-14, 1.125431e-14, 1.127334e-14, 1.130856e-14, 
    1.130037e-14, 1.132981e-14, 1.102961e-14, 1.104761e-14, 1.1046e-14, 
    1.106483e-14, 1.107876e-14, 1.110899e-14, 1.115746e-14, 1.113919e-14, 
    1.117265e-14, 1.117938e-14, 1.112847e-14, 1.115971e-14, 1.105948e-14, 
    1.107565e-14, 1.106599e-14, 1.103076e-14, 1.114326e-14, 1.108549e-14, 
    1.119211e-14, 1.116079e-14, 1.125209e-14, 1.120668e-14, 1.129586e-14, 
    1.133405e-14, 1.136991e-14, 1.141187e-14, 1.105741e-14, 1.104514e-14, 
    1.106704e-14, 1.109739e-14, 1.112549e-14, 1.116292e-14, 1.116672e-14, 
    1.11737e-14, 1.119184e-14, 1.120712e-14, 1.117589e-14, 1.12109e-14, 
    1.10794e-14, 1.114826e-14, 1.104028e-14, 1.10728e-14, 1.109534e-14, 
    1.108543e-14, 1.113687e-14, 1.114897e-14, 1.119827e-14, 1.117277e-14, 
    1.132458e-14, 1.125739e-14, 1.144378e-14, 1.139168e-14, 1.104084e-14, 
    1.105729e-14, 1.111464e-14, 1.108734e-14, 1.116536e-14, 1.118458e-14, 
    1.120016e-14, 1.122015e-14, 1.122226e-14, 1.123411e-14, 1.121466e-14, 
    1.12333e-14, 1.11628e-14, 1.119429e-14, 1.110786e-14, 1.112887e-14, 
    1.111918e-14, 1.110854e-14, 1.114126e-14, 1.117618e-14, 1.117688e-14, 
    1.118805e-14, 1.121963e-14, 1.116533e-14, 1.133321e-14, 1.122952e-14, 
    1.107524e-14, 1.110698e-14, 1.111147e-14, 1.109917e-14, 1.11826e-14, 
    1.115236e-14, 1.123381e-14, 1.121176e-14, 1.124782e-14, 1.122989e-14, 
    1.122722e-14, 1.120419e-14, 1.118981e-14, 1.115361e-14, 1.11241e-14, 
    1.110074e-14, 1.110613e-14, 1.11318e-14, 1.117825e-14, 1.122224e-14, 
    1.121258e-14, 1.124485e-14, 1.115932e-14, 1.119518e-14, 1.118129e-14, 
    1.121741e-14, 1.113864e-14, 1.12061e-14, 1.112138e-14, 1.112877e-14, 
    1.115171e-14, 1.119791e-14, 1.120806e-14, 1.121898e-14, 1.12122e-14, 
    1.117957e-14, 1.117419e-14, 1.115102e-14, 1.114462e-14, 1.112699e-14, 
    1.111236e-14, 1.11257e-14, 1.113967e-14, 1.117943e-14, 1.121525e-14, 
    1.12543e-14, 1.126385e-14, 1.130953e-14, 1.127234e-14, 1.13337e-14, 
    1.128153e-14, 1.137178e-14, 1.120993e-14, 1.128034e-14, 1.115275e-14, 
    1.116646e-14, 1.119131e-14, 1.124829e-14, 1.121747e-14, 1.125348e-14, 
    1.117397e-14, 1.113273e-14, 1.112202e-14, 1.110213e-14, 1.112244e-14, 
    1.112079e-14, 1.114024e-14, 1.113395e-14, 1.11807e-14, 1.115558e-14, 
    1.122691e-14, 1.125297e-14, 1.132652e-14, 1.137161e-14, 1.141751e-14, 
    1.143776e-14, 1.144392e-14, 1.144648e-14 ;

 DISPVEGC =
  0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 0.1735638, 
    0.1735638, 0.1735638 ;

 DISPVEGN =
  0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959, 0.003631959, 0.003631959, 
    0.003631959, 0.003631959, 0.003631959 ;

 DSTDEP =
  2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 2.347785e-12, 
    2.347785e-12, 2.347785e-12, 2.347785e-12 ;

 DSTFLXT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_NFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_GRND_LAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 EFLX_LH_TOT =
  6.257064, 6.273336, 6.270175, 6.28331, 6.276031, 6.284628, 6.260372, 
    6.273972, 6.265294, 6.258544, 6.308742, 6.283899, 6.334722, 6.318814, 
    6.360476, 6.332225, 6.365878, 6.359734, 6.378316, 6.372989, 6.396751, 
    6.380776, 6.409156, 6.392949, 6.395471, 6.380245, 6.288925, 6.305635, 
    6.28793, 6.290312, 6.28925, 6.276171, 6.269567, 6.255841, 6.258336, 
    6.268428, 6.291384, 6.283615, 6.303249, 6.302806, 6.324682, 6.314816, 
    6.353277, 6.341199, 6.373212, 6.365537, 6.372846, 6.370632, 6.372875, 
    6.361624, 6.36644, 6.356558, 6.316658, 6.327885, 6.294414, 6.274263, 
    6.260962, 6.25152, 6.252854, 6.255393, 6.268486, 6.280848, 6.290258, 
    6.296541, 6.302742, 6.321459, 6.331442, 6.35539, 6.351368, 6.358202, 
    6.364775, 6.375791, 6.37398, 6.378832, 6.35804, 6.371841, 6.349073, 
    6.355289, 6.304333, 6.285721, 6.27771, 6.270779, 6.253878, 6.26554, 
    6.260938, 6.271912, 6.278882, 6.275437, 6.296713, 6.288447, 6.332035, 
    6.31324, 6.364008, 6.352196, 6.366847, 6.359371, 6.372177, 6.360651, 
    6.380647, 6.384997, 6.382021, 6.393495, 6.36001, 6.372836, 6.275336, 
    6.275898, 6.278523, 6.266988, 6.266289, 6.255768, 6.265137, 6.269124, 
    6.279294, 6.285299, 6.290998, 6.30354, 6.317551, 6.337207, 6.35296, 
    6.362486, 6.356649, 6.361801, 6.356038, 6.353343, 6.38336, 6.366478, 
    6.391843, 6.39044, 6.378942, 6.390599, 6.276293, 6.273062, 6.261827, 
    6.270618, 6.254625, 6.26356, 6.268696, 6.2886, 6.292987, 6.297029, 
    6.30504, 6.31532, 6.333368, 6.350708, 6.365162, 6.364104, 6.364475, 
    6.367698, 6.359704, 6.369013, 6.370566, 6.366489, 6.390252, 6.383455, 
    6.39041, 6.385986, 6.274115, 6.279557, 6.276614, 6.282145, 6.27824, 
    6.295551, 6.300739, 6.325082, 6.315112, 6.331014, 6.316733, 6.319256, 
    6.331492, 6.317511, 6.349818, 6.327353, 6.367824, 6.345267, 6.369139, 
    6.365099, 6.371799, 6.377794, 6.385363, 6.399323, 6.396091, 6.407802, 
    6.287682, 6.294719, 6.294116, 6.301501, 6.306962, 6.31883, 6.337878, 
    6.330713, 6.343891, 6.348107, 6.326526, 6.338786, 6.299446, 6.305773, 
    6.302018, 6.288226, 6.332338, 6.309666, 6.353191, 6.339287, 6.376936, 
    6.358944, 6.394309, 6.409437, 6.4238, 6.440518, 6.298582, 6.293795, 
    6.302384, 6.314251, 6.325317, 6.340034, 6.341552, 6.344307, 6.353055, 
    6.359085, 6.345161, 6.3606, 6.307205, 6.334319, 6.291969, 6.304678, 
    6.31356, 6.309682, 6.329899, 6.334667, 6.355653, 6.344043, 6.405683, 
    6.379033, 6.453344, 6.432476, 6.292119, 6.298573, 6.321049, 6.310356, 
    6.341028, 6.350169, 6.356347, 6.364224, 6.365089, 6.369764, 6.362103, 
    6.369469, 6.340065, 6.354059, 6.318501, 6.326742, 6.322955, 6.318791, 
    6.33165, 6.345351, 6.345673, 6.351646, 6.364004, 6.341152, 6.409071, 
    6.367958, 6.305617, 6.318035, 6.319843, 6.315027, 6.349408, 6.335922, 
    6.369655, 6.36095, 6.375227, 6.368125, 6.36708, 6.35798, 6.352314, 
    6.336462, 6.324881, 6.315729, 6.317858, 6.327917, 6.346196, 6.365154, 
    6.361337, 6.374142, 6.338798, 6.354488, 6.349015, 6.363302, 6.330516, 
    6.358564, 6.323759, 6.326671, 6.335686, 6.355427, 6.359501, 6.363801, 
    6.361154, 6.348241, 6.34457, 6.335474, 6.33295, 6.326039, 6.320311, 
    6.325537, 6.331025, 6.348259, 6.362404, 6.377875, 6.381678, 6.399734, 
    6.384988, 6.409294, 6.388557, 6.42453, 6.360147, 6.388014, 6.336106, 
    6.341512, 6.352848, 6.375375, 6.363235, 6.37745, 6.34449, 6.328249, 
    6.32409, 6.316279, 6.324269, 6.32362, 6.331274, 6.328815, 6.348781, 
    6.337322, 6.367045, 6.377345, 6.406561, 6.424519, 6.442905, 6.45102, 
    6.453496, 6.454528 ;

 EFLX_LH_TOT_R =
  6.257064, 6.273336, 6.270175, 6.28331, 6.276031, 6.284628, 6.260372, 
    6.273972, 6.265294, 6.258544, 6.308742, 6.283899, 6.334722, 6.318814, 
    6.360476, 6.332225, 6.365878, 6.359734, 6.378316, 6.372989, 6.396751, 
    6.380776, 6.409156, 6.392949, 6.395471, 6.380245, 6.288925, 6.305635, 
    6.28793, 6.290312, 6.28925, 6.276171, 6.269567, 6.255841, 6.258336, 
    6.268428, 6.291384, 6.283615, 6.303249, 6.302806, 6.324682, 6.314816, 
    6.353277, 6.341199, 6.373212, 6.365537, 6.372846, 6.370632, 6.372875, 
    6.361624, 6.36644, 6.356558, 6.316658, 6.327885, 6.294414, 6.274263, 
    6.260962, 6.25152, 6.252854, 6.255393, 6.268486, 6.280848, 6.290258, 
    6.296541, 6.302742, 6.321459, 6.331442, 6.35539, 6.351368, 6.358202, 
    6.364775, 6.375791, 6.37398, 6.378832, 6.35804, 6.371841, 6.349073, 
    6.355289, 6.304333, 6.285721, 6.27771, 6.270779, 6.253878, 6.26554, 
    6.260938, 6.271912, 6.278882, 6.275437, 6.296713, 6.288447, 6.332035, 
    6.31324, 6.364008, 6.352196, 6.366847, 6.359371, 6.372177, 6.360651, 
    6.380647, 6.384997, 6.382021, 6.393495, 6.36001, 6.372836, 6.275336, 
    6.275898, 6.278523, 6.266988, 6.266289, 6.255768, 6.265137, 6.269124, 
    6.279294, 6.285299, 6.290998, 6.30354, 6.317551, 6.337207, 6.35296, 
    6.362486, 6.356649, 6.361801, 6.356038, 6.353343, 6.38336, 6.366478, 
    6.391843, 6.39044, 6.378942, 6.390599, 6.276293, 6.273062, 6.261827, 
    6.270618, 6.254625, 6.26356, 6.268696, 6.2886, 6.292987, 6.297029, 
    6.30504, 6.31532, 6.333368, 6.350708, 6.365162, 6.364104, 6.364475, 
    6.367698, 6.359704, 6.369013, 6.370566, 6.366489, 6.390252, 6.383455, 
    6.39041, 6.385986, 6.274115, 6.279557, 6.276614, 6.282145, 6.27824, 
    6.295551, 6.300739, 6.325082, 6.315112, 6.331014, 6.316733, 6.319256, 
    6.331492, 6.317511, 6.349818, 6.327353, 6.367824, 6.345267, 6.369139, 
    6.365099, 6.371799, 6.377794, 6.385363, 6.399323, 6.396091, 6.407802, 
    6.287682, 6.294719, 6.294116, 6.301501, 6.306962, 6.31883, 6.337878, 
    6.330713, 6.343891, 6.348107, 6.326526, 6.338786, 6.299446, 6.305773, 
    6.302018, 6.288226, 6.332338, 6.309666, 6.353191, 6.339287, 6.376936, 
    6.358944, 6.394309, 6.409437, 6.4238, 6.440518, 6.298582, 6.293795, 
    6.302384, 6.314251, 6.325317, 6.340034, 6.341552, 6.344307, 6.353055, 
    6.359085, 6.345161, 6.3606, 6.307205, 6.334319, 6.291969, 6.304678, 
    6.31356, 6.309682, 6.329899, 6.334667, 6.355653, 6.344043, 6.405683, 
    6.379033, 6.453344, 6.432476, 6.292119, 6.298573, 6.321049, 6.310356, 
    6.341028, 6.350169, 6.356347, 6.364224, 6.365089, 6.369764, 6.362103, 
    6.369469, 6.340065, 6.354059, 6.318501, 6.326742, 6.322955, 6.318791, 
    6.33165, 6.345351, 6.345673, 6.351646, 6.364004, 6.341152, 6.409071, 
    6.367958, 6.305617, 6.318035, 6.319843, 6.315027, 6.349408, 6.335922, 
    6.369655, 6.36095, 6.375227, 6.368125, 6.36708, 6.35798, 6.352314, 
    6.336462, 6.324881, 6.315729, 6.317858, 6.327917, 6.346196, 6.365154, 
    6.361337, 6.374142, 6.338798, 6.354488, 6.349015, 6.363302, 6.330516, 
    6.358564, 6.323759, 6.326671, 6.335686, 6.355427, 6.359501, 6.363801, 
    6.361154, 6.348241, 6.34457, 6.335474, 6.33295, 6.326039, 6.320311, 
    6.325537, 6.331025, 6.348259, 6.362404, 6.377875, 6.381678, 6.399734, 
    6.384988, 6.409294, 6.388557, 6.42453, 6.360147, 6.388014, 6.336106, 
    6.341512, 6.352848, 6.375375, 6.363235, 6.37745, 6.34449, 6.328249, 
    6.32409, 6.316279, 6.324269, 6.32362, 6.331274, 6.328815, 6.348781, 
    6.337322, 6.367045, 6.377345, 6.406561, 6.424519, 6.442905, 6.45102, 
    6.453496, 6.454528 ;

 EFLX_LH_TOT_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 ELAI =
  0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122 ;

 ER =
  6.358388e-08, 6.386347e-08, 6.380911e-08, 6.403462e-08, 6.390952e-08, 
    6.405718e-08, 6.364056e-08, 6.387457e-08, 6.372518e-08, 6.360905e-08, 
    6.447225e-08, 6.404468e-08, 6.491634e-08, 6.464366e-08, 6.532863e-08, 
    6.487392e-08, 6.542031e-08, 6.53155e-08, 6.563094e-08, 6.554057e-08, 
    6.594404e-08, 6.567264e-08, 6.615318e-08, 6.587923e-08, 6.592209e-08, 
    6.566369e-08, 6.413072e-08, 6.441902e-08, 6.411364e-08, 6.415475e-08, 
    6.41363e-08, 6.391211e-08, 6.379913e-08, 6.356251e-08, 6.360547e-08, 
    6.377926e-08, 6.417324e-08, 6.403949e-08, 6.437654e-08, 6.436893e-08, 
    6.474416e-08, 6.457498e-08, 6.520563e-08, 6.502638e-08, 6.554434e-08, 
    6.541408e-08, 6.553822e-08, 6.550058e-08, 6.553871e-08, 6.534768e-08, 
    6.542952e-08, 6.526142e-08, 6.460666e-08, 6.47991e-08, 6.422516e-08, 
    6.388007e-08, 6.365083e-08, 6.348817e-08, 6.351116e-08, 6.3555e-08, 
    6.378028e-08, 6.399208e-08, 6.415348e-08, 6.426145e-08, 6.436783e-08, 
    6.468986e-08, 6.486028e-08, 6.524188e-08, 6.5173e-08, 6.528968e-08, 
    6.540112e-08, 6.558825e-08, 6.555744e-08, 6.563989e-08, 6.528659e-08, 
    6.55214e-08, 6.513378e-08, 6.52398e-08, 6.439678e-08, 6.407557e-08, 
    6.393907e-08, 6.381956e-08, 6.352884e-08, 6.372961e-08, 6.365047e-08, 
    6.383875e-08, 6.395839e-08, 6.389921e-08, 6.426441e-08, 6.412242e-08, 
    6.487038e-08, 6.454822e-08, 6.538812e-08, 6.518714e-08, 6.54363e-08, 
    6.530916e-08, 6.5527e-08, 6.533094e-08, 6.567057e-08, 6.574452e-08, 
    6.569399e-08, 6.588811e-08, 6.532007e-08, 6.553822e-08, 6.389756e-08, 
    6.390721e-08, 6.395216e-08, 6.375454e-08, 6.374245e-08, 6.356133e-08, 
    6.372249e-08, 6.379111e-08, 6.396532e-08, 6.406837e-08, 6.416632e-08, 
    6.438169e-08, 6.462222e-08, 6.495855e-08, 6.520017e-08, 6.536213e-08, 
    6.526282e-08, 6.53505e-08, 6.525248e-08, 6.520654e-08, 6.571682e-08, 
    6.543029e-08, 6.586019e-08, 6.58364e-08, 6.564185e-08, 6.583908e-08, 
    6.391399e-08, 6.385844e-08, 6.366564e-08, 6.381653e-08, 6.354161e-08, 
    6.36955e-08, 6.378399e-08, 6.41254e-08, 6.420041e-08, 6.426996e-08, 
    6.440733e-08, 6.458363e-08, 6.489289e-08, 6.516198e-08, 6.54076e-08, 
    6.538961e-08, 6.539594e-08, 6.545082e-08, 6.531489e-08, 6.547314e-08, 
    6.54997e-08, 6.543026e-08, 6.583321e-08, 6.571809e-08, 6.58359e-08, 
    6.576094e-08, 6.38765e-08, 6.396994e-08, 6.391945e-08, 6.40144e-08, 
    6.394751e-08, 6.424496e-08, 6.433414e-08, 6.475143e-08, 6.458016e-08, 
    6.485271e-08, 6.460785e-08, 6.465124e-08, 6.486162e-08, 6.462108e-08, 
    6.514714e-08, 6.47905e-08, 6.545295e-08, 6.509682e-08, 6.547527e-08, 
    6.540655e-08, 6.552033e-08, 6.562224e-08, 6.575045e-08, 6.598701e-08, 
    6.593223e-08, 6.613006e-08, 6.410925e-08, 6.423046e-08, 6.421978e-08, 
    6.434662e-08, 6.444042e-08, 6.464373e-08, 6.496981e-08, 6.484719e-08, 
    6.507229e-08, 6.511748e-08, 6.477549e-08, 6.498548e-08, 6.431157e-08, 
    6.442045e-08, 6.435562e-08, 6.411882e-08, 6.487545e-08, 6.448715e-08, 
    6.520416e-08, 6.499381e-08, 6.560771e-08, 6.530242e-08, 6.590207e-08, 
    6.615844e-08, 6.639969e-08, 6.668164e-08, 6.42966e-08, 6.421424e-08, 
    6.43617e-08, 6.456572e-08, 6.4755e-08, 6.500665e-08, 6.503239e-08, 
    6.507953e-08, 6.520164e-08, 6.530431e-08, 6.509445e-08, 6.533005e-08, 
    6.444572e-08, 6.490915e-08, 6.418311e-08, 6.440175e-08, 6.455369e-08, 
    6.448703e-08, 6.483317e-08, 6.491475e-08, 6.524627e-08, 6.507489e-08, 
    6.609517e-08, 6.564377e-08, 6.689631e-08, 6.654629e-08, 6.418547e-08, 
    6.429631e-08, 6.468208e-08, 6.449854e-08, 6.502344e-08, 6.515264e-08, 
    6.525767e-08, 6.539194e-08, 6.540643e-08, 6.548598e-08, 6.535562e-08, 
    6.548083e-08, 6.500718e-08, 6.521884e-08, 6.463799e-08, 6.477936e-08, 
    6.471433e-08, 6.464298e-08, 6.486317e-08, 6.509775e-08, 6.510275e-08, 
    6.517797e-08, 6.538995e-08, 6.502557e-08, 6.615345e-08, 6.545692e-08, 
    6.441718e-08, 6.463069e-08, 6.466117e-08, 6.457847e-08, 6.513969e-08, 
    6.493634e-08, 6.548404e-08, 6.533602e-08, 6.557855e-08, 6.545803e-08, 
    6.54403e-08, 6.528551e-08, 6.518914e-08, 6.494567e-08, 6.474756e-08, 
    6.459047e-08, 6.4627e-08, 6.479956e-08, 6.51121e-08, 6.540775e-08, 
    6.534299e-08, 6.556012e-08, 6.498538e-08, 6.522639e-08, 6.513324e-08, 
    6.537611e-08, 6.484393e-08, 6.529714e-08, 6.472809e-08, 6.477798e-08, 
    6.493231e-08, 6.524274e-08, 6.53114e-08, 6.538474e-08, 6.533948e-08, 
    6.512003e-08, 6.508407e-08, 6.492856e-08, 6.488562e-08, 6.476711e-08, 
    6.466901e-08, 6.475865e-08, 6.485278e-08, 6.512012e-08, 6.536104e-08, 
    6.562369e-08, 6.568797e-08, 6.599488e-08, 6.574506e-08, 6.615733e-08, 
    6.580684e-08, 6.641355e-08, 6.532339e-08, 6.579651e-08, 6.493933e-08, 
    6.503167e-08, 6.519871e-08, 6.558179e-08, 6.537497e-08, 6.561685e-08, 
    6.508266e-08, 6.480552e-08, 6.47338e-08, 6.460002e-08, 6.473686e-08, 
    6.472573e-08, 6.485668e-08, 6.48146e-08, 6.512899e-08, 6.496011e-08, 
    6.543986e-08, 6.561493e-08, 6.610933e-08, 6.641241e-08, 6.672092e-08, 
    6.685712e-08, 6.689857e-08, 6.69159e-08 ;

 ERRH2O =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 ERRH2OSNO =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 ERRSEB =
  -1.053313e-14, -8.699309e-16, -1.602822e-14, -7.371716e-15, -5.029286e-15, 
    -1.340398e-14, -1.336219e-14, -1.143902e-14, -1.319324e-14, 1.808731e-15, 
    -6.351236e-15, -1.016574e-14, -1.314459e-14, -8.039349e-15, 
    -1.241416e-14, -6.043374e-15, -2.259766e-14, -7.866874e-15, 
    -1.109628e-14, -1.07206e-14, -5.427586e-15, -1.768885e-14, -1.224179e-14, 
    -1.441249e-14, -1.501101e-14, -2.450391e-14, -1.868933e-14, 
    -2.077158e-15, -1.094377e-14, -1.513513e-14, -6.698661e-15, 
    -7.815619e-15, -1.311137e-14, -1.012186e-14, -5.959289e-15, -1.26745e-15, 
    -6.280636e-15, -2.438427e-15, -1.171454e-14, -1.277582e-14, 
    -1.131977e-14, -4.364106e-15, -4.501632e-15, -8.902969e-15, 2.162014e-15, 
    -6.814942e-15, -1.243615e-14, -1.130549e-14, -7.54729e-15, -6.266311e-15, 
    -7.37178e-15, 1.087319e-15, -1.395234e-14, -1.546415e-14, -1.249528e-14, 
    -1.695866e-14, -9.369465e-15, -5.651065e-15, -1.78993e-15, -1.673835e-14, 
    -1.556529e-14, -1.091806e-14, -1.572832e-14, -2.237173e-15, 
    -1.661143e-14, -1.204155e-14, -4.751109e-15, -2.049015e-14, 
    -1.660581e-14, -1.208397e-14, -1.552576e-14, -7.93124e-15, -9.432355e-15, 
    -1.023809e-14, -1.290397e-14, -8.177498e-15, -8.84312e-15, -1.316013e-14, 
    -4.728607e-15, -1.179538e-14, -8.429735e-15, -8.490905e-15, 
    -9.899004e-15, -1.405593e-14, -1.106075e-14, -1.793059e-14, 
    -8.755658e-15, -2.364313e-15, -2.833433e-15, -7.886077e-15, 
    -7.385713e-15, -1.661434e-14, -5.032269e-15, -9.886239e-15, 
    -9.693221e-15, -1.40377e-14, -9.041399e-15, -1.139155e-14, -9.973731e-15, 
    -6.272298e-15, -7.127709e-15, -1.076657e-14, -7.187108e-15, 
    -1.121365e-14, -1.122835e-14, -1.64806e-14, -8.507869e-15, -7.660613e-15, 
    -1.626585e-14, -2.26274e-15, -1.155358e-14, -6.733264e-15, -4.762765e-15, 
    1.25352e-15, -3.260113e-17, -4.795735e-15, -1.064453e-14, -3.968613e-15, 
    -8.108688e-15, -9.037883e-15, -1.000065e-14, -1.562457e-14, 
    -1.622849e-14, -1.648379e-14, -1.027772e-14, -1.517898e-14, 
    -1.477495e-14, -9.628307e-15, -3.248537e-15, -1.785506e-14, 
    -1.400419e-14, -6.207885e-15, -1.726228e-14, -1.448213e-14, 
    -1.629336e-14, -6.785617e-15, -7.109593e-15, -5.825849e-15, 
    -1.424195e-14, -1.456014e-14, -1.405533e-14, -6.591279e-15, 
    -1.618264e-14, 1.820294e-16, -1.112845e-14, -6.725151e-15, -1.64705e-14, 
    -9.681121e-15, -6.42374e-15, -5.19824e-15, -1.042711e-14, -1.519215e-14, 
    -1.270663e-14, -1.323337e-14, -1.803796e-15, -1.096906e-14, 
    -5.731919e-15, 3.990911e-17, -4.985185e-15, -8.035304e-15, -9.691286e-15, 
    -7.432891e-15, -7.702077e-15, -3.310563e-15, -1.177629e-14, 
    -1.142949e-14, -1.287394e-14, -4.145745e-15, -1.894322e-14, 
    -4.083134e-15, -1.580036e-14, -1.321846e-14, -1.481669e-14, 
    -1.510152e-14, -9.213716e-15, -1.248358e-14, -1.697648e-14, 
    -1.230256e-14, -1.250956e-14, -1.855058e-14, -4.99417e-15, -2.743905e-15, 
    1.031351e-15, -1.29076e-14, -1.478074e-14, -1.364245e-14, -1.140283e-14, 
    -4.389402e-15, -1.739589e-15, -3.165486e-15, -1.268234e-14, 
    -2.305677e-14, -6.695962e-15, -1.84876e-14, -6.102727e-15, -1.127535e-14, 
    -1.451179e-14, -1.26007e-14, -1.11392e-14, -1.27976e-14, -1.404705e-14, 
    -1.558802e-14, -1.392889e-14, -8.90018e-15, -8.789849e-15, -1.276235e-14, 
    -1.911267e-14, -1.426556e-14, -1.087911e-14, -4.463036e-15, 
    -5.485711e-15, -1.329055e-14, 5.12898e-16, -6.375071e-15, -3.225053e-15, 
    -1.654468e-14, -9.92638e-15, -1.330885e-14, -2.490386e-15, -9.045378e-15, 
    -1.566735e-14, -2.910854e-15, -1.290031e-14, -1.038301e-14, 
    -4.001604e-15, -5.768823e-15, -2.140405e-15, -1.654102e-14, 
    -1.001677e-14, -9.673664e-15, -2.557437e-15, -1.29631e-14, -1.295457e-14, 
    -8.445686e-15, -8.216403e-15, -1.203967e-14, 1.853344e-15, -8.70483e-15, 
    -1.001491e-15, -5.124247e-16, -1.42726e-14, -5.181331e-15, -1.116796e-14, 
    -2.274718e-15, -7.418719e-15, -1.404445e-14, -8.276093e-15, 
    -5.036296e-15, -1.316149e-14, -1.039251e-14, -1.439116e-14, 
    -1.065918e-14, -1.738716e-14, -7.439621e-15, -1.549085e-14, 
    -1.514036e-14, -2.001386e-14, -1.010933e-14, -1.226672e-14, 
    -2.177959e-14, -1.234264e-14, 8.048573e-16, -1.740949e-14, -8.400019e-15, 
    -1.202079e-14, -7.794442e-15, -1.483278e-14, -5.114677e-15, 
    -1.071163e-14, -7.945765e-15, -7.197081e-15, -1.01325e-14, -9.410236e-15, 
    -6.966376e-15, -8.130203e-15, -1.375013e-14, -1.044085e-14, 
    -8.750309e-15, -1.172131e-14, -7.239302e-15, -3.964436e-15, 
    -1.007552e-14, -1.315425e-14, -1.642577e-14, -5.263744e-15, 
    -1.097125e-14, -1.431619e-15, -2.170512e-14, -3.724356e-15, 
    -1.072958e-14, -9.461915e-15, -1.03674e-14, -4.876308e-15, -1.029846e-14, 
    -7.709762e-15, -1.105344e-14, -3.07541e-15, -1.028082e-14, -2.079139e-15, 
    -1.303432e-14, -2.080964e-14, -6.110069e-15, -1.217172e-14, 
    -9.884825e-15, -1.25409e-14, -8.231585e-15, -8.104746e-15, -7.047064e-15, 
    -1.006634e-14, -1.793697e-14, -9.275433e-15, -1.337089e-14, 
    -2.178819e-14, -8.972363e-15, -1.5938e-14, -8.875955e-15, -1.145503e-14, 
    -6.90242e-15, -8.15315e-15, -7.933089e-15, -7.936789e-15, -1.074087e-14, 
    -8.427038e-15, -1.689644e-14, 5.622376e-17, -1.194212e-14, -9.096164e-15, 
    -1.192986e-14, -1.563313e-14, -1.189722e-14, -3.510844e-15, 
    -1.759615e-14, -1.973349e-14, -1.179447e-14, -1.665455e-14, 
    -1.221551e-14, -5.956403e-15, -1.241767e-14 ;

 ERRSOI =
  -71.24087, -71.33397, -71.31628, -71.3905, -71.35, -71.39811, -71.26054, 
    -71.33696, -71.28863, -71.25035, -71.53255, -71.39401, -71.68469, 
    -71.59469, -71.82368, -71.66957, -71.85513, -71.82108, -71.92818, 
    -71.89758, -72.03098, -71.94232, -72.10334, -72.01078, -72.02454, 
    -71.9391, -71.42362, -71.51469, -71.41781, -71.43089, -71.42544, 
    -71.3502, -71.31114, -71.23501, -71.24916, -71.30576, -71.43681, 
    -71.39349, -71.50633, -71.50382, -71.62858, -71.57224, -71.78399, 
    -71.72404, -71.8989, -71.85459, -71.89649, -71.88402, -71.89666, 
    -71.83181, -71.85948, -71.80305, -71.58244, -71.64655, -71.45469, 
    -71.337, -71.26357, -71.21014, -71.21768, -71.2317, -71.30606, -71.37767, 
    -71.43178, -71.46773, -71.50343, -71.60693, -71.66586, -71.79521, 
    -71.77341, -71.81155, -71.85027, -71.91322, -71.90308, -71.93047, 
    -71.81168, -71.89002, -71.76064, -71.79578, -71.5069, -71.40545, 
    -71.35706, -71.31945, -71.22336, -71.28936, -71.26318, -71.32681, 
    -71.36637, -71.34705, -71.46872, -71.42113, -71.66936, -71.56229, 
    -71.84576, -71.77802, -71.86224, -71.81955, -71.89221, -71.82683, 
    -71.94117, -71.96539, -71.9487, -72.01498, -71.82304, -71.8959, 
    -71.34621, -71.34933, -71.36456, -71.29752, -71.29379, -71.23431, 
    -71.28779, -71.31007, -71.36916, -71.40298, -71.43558, -71.50743, 
    -71.58677, -71.69984, -71.78233, -71.83739, -71.80403, -71.83344, 
    -71.80033, -71.7851, -71.9559, -71.85936, -72.00542, -71.99754, 
    -71.93087, -71.99845, -71.35162, -71.33351, -71.2687, -71.31943, 
    -71.22793, -71.27834, -71.30688, -71.42077, -71.44733, -71.47002, 
    -71.51633, -71.57509, -71.67798, -71.76885, -71.85279, -71.84676, 
    -71.84882, -71.86694, -71.82119, -71.87452, -71.88287, -71.86009, 
    -71.99646, -71.95753, -71.99738, -71.97218, -71.33955, -71.37032, 
    -71.35359, -71.38471, -71.36228, -71.4603, -71.48969, -71.62943, 
    -71.57358, -71.66422, -71.58327, -71.59724, -71.66454, -71.58805, 
    -71.76264, -71.64179, -71.86767, -71.74413, -71.87526, -71.85241, 
    -71.89087, -71.92465, -71.96836, -72.04733, -72.02928, -72.09644, 
    -71.4168, -71.45623, -71.45392, -71.49605, -71.52695, -71.59553, 
    -71.70437, -71.66377, -71.73962, -71.75455, -71.63995, -71.70908, 
    -71.48352, -71.51865, -71.4986, -71.41922, -71.67151, -71.5411, 
    -71.78348, -71.71272, -71.91968, -71.81544, -72.01907, -72.10339, 
    -72.18842, -72.2816, -71.47904, -71.4521, -71.50139, -71.56753, 
    -71.63233, -71.71681, -71.72611, -71.74161, -71.78336, -71.81782, 
    -71.74537, -71.82659, -71.52444, -71.6834, -71.44083, -71.51214, 
    -71.56414, -71.54251, -71.65944, -71.68663, -71.79702, -71.74054, 
    -72.08152, -71.93013, -72.35668, -72.23619, -71.44241, -71.4795, 
    -71.60713, -71.54653, -71.72309, -71.76624, -71.80231, -71.84653, 
    -71.85217, -71.87856, -71.8352, -71.8773, -71.71699, -71.78878, 
    -71.59393, -71.64054, -71.6195, -71.59554, -71.66935, -71.74622, 
    -71.74976, -71.77421, -71.83955, -71.72383, -72.0976, -71.86306, 
    -71.51985, -71.58887, -71.60104, -71.57388, -71.76186, -71.69333, 
    -71.87819, -71.82857, -71.91041, -71.86954, -71.86345, -71.81149, 
    -71.77868, -71.6961, -71.62968, -71.57805, -71.59019, -71.64698, 
    -71.75136, -71.85184, -71.82956, -71.90421, -71.71017, -71.79048, 
    -71.75883, -71.84176, -71.66227, -71.80934, -71.62415, -71.64073, 
    -71.69199, -71.79466, -71.82021, -71.8441, -71.82976, -71.75447, 
    -71.7429, -71.69121, -71.67601, -71.63726, -71.60432, -71.63394, 
    -71.66468, -71.75529, -71.83598, -71.92486, -71.94736, -72.04677, 
    -71.9632, -72.09853, -71.97948, -72.18777, -71.82066, -71.97987, 
    -71.69496, -71.726, -71.78025, -71.9089, -71.84138, -71.92127, -71.74261, 
    -71.64799, -71.62591, -71.58083, -71.62694, -71.62326, -71.6673, 
    -71.65326, -71.75833, -71.70187, -71.86279, -71.92111, -72.0887, 
    -72.19061, -72.29771, -72.34407, -72.35837, -72.36423 ;

 ERRSOL =
  4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 4.625929e-18, 
    4.625929e-18, 4.625929e-18, 4.625929e-18 ;

 ESAI =
  0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173 ;

 FAREA_BURNED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCEV =
  -1.94949, -1.948384, -1.948594, -1.947711, -1.948193, -1.947621, -1.949256, 
    -1.948349, -1.948922, -1.949376, -1.946018, -1.947669, -1.944212, 
    -1.945276, -1.94257, -1.944392, -1.942195, -1.942599, -1.941323, 
    -1.941688, -1.940096, -1.941154, -1.939227, -1.940337, -1.940172, 
    -1.941193, -1.947316, -1.946232, -1.947385, -1.94723, -1.947294, 
    -1.948191, -1.948656, -1.949558, -1.949391, -1.948719, -1.947159, 
    -1.947675, -1.946328, -1.946358, -1.944876, -1.945542, -1.94304, 
    -1.943744, -1.941672, -1.9422, -1.941701, -1.94185, -1.941699, -1.942472, 
    -1.942142, -1.942813, -1.945421, -1.944663, -1.946946, -1.948349, 
    -1.94922, -1.949853, -1.949764, -1.949598, -1.948716, -1.947863, 
    -1.947218, -1.946789, -1.946363, -1.945134, -1.944435, -1.942907, 
    -1.943165, -1.942713, -1.942252, -1.941502, -1.941623, -1.941296, 
    -1.942711, -1.941779, -1.943317, -1.9429, -1.946325, -1.947532, -1.94811, 
    -1.948556, -1.949697, -1.948914, -1.949225, -1.948468, -1.947998, 
    -1.948228, -1.946777, -1.947345, -1.944394, -1.94566, -1.942306, 
    -1.943111, -1.942109, -1.942617, -1.941753, -1.942531, -1.941168, 
    -1.940879, -1.941079, -1.940286, -1.942576, -1.941709, -1.948238, 
    -1.948201, -1.948019, -1.948817, -1.948861, -1.949567, -1.948932, 
    -1.948668, -1.947964, -1.947562, -1.947173, -1.946315, -1.945371, 
    -1.944032, -1.94306, -1.942405, -1.942801, -1.942452, -1.942846, 
    -1.943026, -1.940993, -1.942144, -1.9404, -1.940494, -1.941292, 
    -1.940483, -1.948173, -1.948389, -1.949159, -1.948556, -1.949642, 
    -1.949045, -1.948706, -1.94735, -1.947033, -1.946762, -1.946209, 
    -1.945508, -1.944291, -1.94322, -1.942222, -1.942294, -1.942269, 
    -1.942053, -1.942598, -1.941963, -1.941864, -1.942135, -1.940507, 
    -1.940973, -1.940496, -1.940798, -1.948317, -1.947951, -1.94815, 
    -1.94778, -1.948047, -1.946879, -1.946528, -1.944867, -1.945526, 
    -1.944454, -1.945411, -1.945246, -1.944452, -1.945354, -1.943295, 
    -1.944721, -1.942045, -1.943508, -1.941954, -1.942226, -1.941768, 
    -1.941366, -1.940843, -1.939899, -1.940115, -1.93931, -1.947397, 
    -1.946927, -1.946954, -1.946451, -1.946082, -1.945266, -1.943978, 
    -1.944458, -1.94356, -1.943389, -1.944741, -1.943922, -1.946601, 
    -1.946182, -1.946421, -1.947368, -1.944368, -1.945913, -1.943046, 
    -1.943879, -1.941425, -1.942667, -1.940237, -1.939228, -1.938203, 
    -1.937081, -1.946655, -1.946976, -1.946387, -1.945599, -1.944831, 
    -1.94383, -1.94372, -1.943536, -1.943047, -1.942638, -1.943493, 
    -1.942533, -1.946115, -1.944227, -1.947111, -1.94626, -1.945639, 
    -1.945896, -1.94451, -1.944188, -1.942886, -1.943549, -1.939491, 
    -1.941301, -1.936172, -1.937629, -1.947091, -1.946649, -1.94513, 
    -1.945848, -1.943756, -1.943251, -1.942822, -1.942297, -1.942229, 
    -1.941915, -1.942431, -1.94193, -1.943828, -1.942983, -1.945285, 
    -1.944734, -1.944982, -1.945266, -1.944392, -1.943483, -1.943439, 
    -1.943156, -1.942384, -1.943747, -1.9393, -1.942103, -1.946166, 
    -1.945346, -1.945201, -1.945522, -1.943303, -1.944109, -1.941919, 
    -1.94251, -1.941535, -1.942022, -1.942095, -1.942713, -1.943103, 
    -1.944076, -1.944863, -1.945473, -1.945329, -1.944658, -1.943421, 
    -1.942234, -1.942499, -1.941609, -1.943909, -1.942963, -1.943339, 
    -1.942353, -1.944477, -1.942742, -1.944927, -1.944731, -1.944124, 
    -1.942914, -1.942609, -1.942326, -1.942496, -1.943391, -1.943521, 
    -1.944133, -1.944314, -1.944772, -1.945162, -1.944812, -1.944448, 
    -1.94338, -1.942422, -1.941363, -1.941094, -1.939908, -1.940907, 
    -1.939289, -1.940715, -1.938215, -1.942606, -1.940709, -1.944089, 
    -1.943721, -1.943085, -1.941555, -1.942358, -1.941407, -1.943525, 
    -1.944647, -1.944907, -1.94544, -1.944895, -1.944938, -1.944417, 
    -1.944583, -1.943344, -1.944007, -1.942103, -1.941409, -1.939403, 
    -1.938178, -1.936885, -1.936324, -1.936151, -1.93608 ;

 FCH4 =
  1.671817e-13, 1.656402e-13, 1.659412e-13, 1.646884e-13, 1.653847e-13, 
    1.645624e-13, 1.668705e-13, 1.655787e-13, 1.664047e-13, 1.670436e-13, 
    1.622262e-13, 1.646322e-13, 1.587796e-13, 1.601956e-13, 1.565869e-13, 
    1.590017e-13, 1.56091e-13, 1.566576e-13, 1.549404e-13, 1.55436e-13, 
    1.532019e-13, 1.547108e-13, 1.52022e-13, 1.535645e-13, 1.533249e-13, 
    1.547601e-13, 1.641511e-13, 1.625279e-13, 1.642467e-13, 1.640165e-13, 
    1.641198e-13, 1.653703e-13, 1.659965e-13, 1.672988e-13, 1.670632e-13, 
    1.661063e-13, 1.639128e-13, 1.646611e-13, 1.62768e-13, 1.62811e-13, 
    1.596769e-13, 1.60548e-13, 1.572474e-13, 1.582002e-13, 1.554153e-13, 
    1.561247e-13, 1.554488e-13, 1.556543e-13, 1.554461e-13, 1.564841e-13, 
    1.560409e-13, 1.569484e-13, 1.603857e-13, 1.593918e-13, 1.636212e-13, 
    1.655483e-13, 1.668141e-13, 1.677054e-13, 1.675798e-13, 1.673399e-13, 
    1.661007e-13, 1.649255e-13, 1.640235e-13, 1.634171e-13, 1.628172e-13, 
    1.599578e-13, 1.590729e-13, 1.570533e-13, 1.574217e-13, 1.567967e-13, 
    1.56195e-13, 1.551749e-13, 1.553436e-13, 1.548912e-13, 1.568132e-13, 
    1.555408e-13, 1.576307e-13, 1.570645e-13, 1.626537e-13, 1.644596e-13, 
    1.652206e-13, 1.658834e-13, 1.674831e-13, 1.663804e-13, 1.668161e-13, 
    1.657772e-13, 1.651131e-13, 1.654419e-13, 1.634005e-13, 1.641975e-13, 
    1.590202e-13, 1.606848e-13, 1.562654e-13, 1.573462e-13, 1.560042e-13, 
    1.566917e-13, 1.555101e-13, 1.565743e-13, 1.547222e-13, 1.543136e-13, 
    1.545931e-13, 1.535148e-13, 1.566329e-13, 1.554488e-13, 1.654511e-13, 
    1.653975e-13, 1.651477e-13, 1.662428e-13, 1.663095e-13, 1.673052e-13, 
    1.664196e-13, 1.660408e-13, 1.650745e-13, 1.644999e-13, 1.639516e-13, 
    1.627389e-13, 1.603058e-13, 1.585579e-13, 1.572766e-13, 1.564059e-13, 
    1.569409e-13, 1.564688e-13, 1.569964e-13, 1.572425e-13, 1.54467e-13, 
    1.560368e-13, 1.536707e-13, 1.538033e-13, 1.548804e-13, 1.537883e-13, 
    1.653599e-13, 1.65668e-13, 1.667327e-13, 1.659002e-13, 1.674132e-13, 
    1.665683e-13, 1.660802e-13, 1.641809e-13, 1.637603e-13, 1.633692e-13, 
    1.625938e-13, 1.605037e-13, 1.589023e-13, 1.574806e-13, 1.561598e-13, 
    1.562573e-13, 1.56223e-13, 1.559253e-13, 1.566609e-13, 1.558039e-13, 
    1.556592e-13, 1.56037e-13, 1.53821e-13, 1.544598e-13, 1.538061e-13, 
    1.542226e-13, 1.655679e-13, 1.650487e-13, 1.653295e-13, 1.648011e-13, 
    1.651736e-13, 1.6351e-13, 1.630075e-13, 1.596393e-13, 1.605214e-13, 
    1.591124e-13, 1.603795e-13, 1.601566e-13, 1.59066e-13, 1.603116e-13, 
    1.575597e-13, 1.594365e-13, 1.559137e-13, 1.578274e-13, 1.557922e-13, 
    1.561656e-13, 1.555465e-13, 1.549883e-13, 1.542808e-13, 1.529606e-13, 
    1.53268e-13, 1.521532e-13, 1.642713e-13, 1.635915e-13, 1.636514e-13, 
    1.62937e-13, 1.624065e-13, 1.601952e-13, 1.584986e-13, 1.591412e-13, 
    1.579573e-13, 1.577174e-13, 1.595143e-13, 1.584161e-13, 1.631348e-13, 
    1.625196e-13, 1.628862e-13, 1.642178e-13, 1.589936e-13, 1.621416e-13, 
    1.572552e-13, 1.583722e-13, 1.550681e-13, 1.567281e-13, 1.534368e-13, 
    1.519923e-13, 1.506132e-13, 1.489787e-13, 1.632192e-13, 1.636825e-13, 
    1.628518e-13, 1.605954e-13, 1.596207e-13, 1.583045e-13, 1.581685e-13, 
    1.57919e-13, 1.572687e-13, 1.567178e-13, 1.578399e-13, 1.565791e-13, 
    1.623766e-13, 1.588172e-13, 1.638574e-13, 1.626255e-13, 1.606569e-13, 
    1.621422e-13, 1.592143e-13, 1.587878e-13, 1.570298e-13, 1.579435e-13, 
    1.523509e-13, 1.548699e-13, 1.477183e-13, 1.497664e-13, 1.638441e-13, 
    1.632208e-13, 1.599977e-13, 1.620769e-13, 1.582158e-13, 1.575303e-13, 
    1.569685e-13, 1.562447e-13, 1.561662e-13, 1.557339e-13, 1.564411e-13, 
    1.557619e-13, 1.583017e-13, 1.571767e-13, 1.602248e-13, 1.594942e-13, 
    1.598312e-13, 1.601991e-13, 1.590578e-13, 1.578224e-13, 1.577957e-13, 
    1.573952e-13, 1.562558e-13, 1.582046e-13, 1.520208e-13, 1.558924e-13, 
    1.625381e-13, 1.602624e-13, 1.601054e-13, 1.605301e-13, 1.575993e-13, 
    1.586745e-13, 1.557445e-13, 1.565469e-13, 1.55228e-13, 1.55886e-13, 
    1.559824e-13, 1.56819e-13, 1.573355e-13, 1.586256e-13, 1.596592e-13, 
    1.604686e-13, 1.602812e-13, 1.593893e-13, 1.577461e-13, 1.561591e-13, 
    1.565094e-13, 1.55329e-13, 1.584166e-13, 1.571363e-13, 1.576337e-13, 
    1.563304e-13, 1.591582e-13, 1.567567e-13, 1.5976e-13, 1.595014e-13, 
    1.586957e-13, 1.570488e-13, 1.566796e-13, 1.562837e-13, 1.565282e-13, 
    1.577039e-13, 1.578949e-13, 1.587154e-13, 1.589404e-13, 1.595578e-13, 
    1.600651e-13, 1.596017e-13, 1.59112e-13, 1.577034e-13, 1.564119e-13, 
    1.549803e-13, 1.546262e-13, 1.529165e-13, 1.543108e-13, 1.519988e-13, 
    1.539682e-13, 1.505337e-13, 1.566152e-13, 1.540254e-13, 1.586588e-13, 
    1.581723e-13, 1.572845e-13, 1.552104e-13, 1.563366e-13, 1.55018e-13, 
    1.579024e-13, 1.593584e-13, 1.597305e-13, 1.604197e-13, 1.597146e-13, 
    1.597722e-13, 1.590916e-13, 1.59311e-13, 1.576562e-13, 1.585496e-13, 
    1.559848e-13, 1.550285e-13, 1.522706e-13, 1.5054e-13, 1.48749e-13, 
    1.479494e-13, 1.477049e-13, 1.476026e-13 ;

 FCH4TOCO2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4_DFSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCOV =
  0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584 ;

 FCTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FGEV =
  8.206553, 8.22172, 8.218769, 8.231021, 8.224223, 8.232248, 8.209627, 
    8.222321, 8.214216, 8.20792, 8.25476, 8.231567, 8.278934, 8.264091, 
    8.303046, 8.276617, 8.308073, 8.302333, 8.319639, 8.314677, 8.336847, 
    8.321931, 8.348383, 8.333286, 8.335643, 8.321438, 8.236241, 8.251867, 
    8.235315, 8.237541, 8.236544, 8.224361, 8.218223, 8.2054, 8.207726, 
    8.217148, 8.238543, 8.23129, 8.249578, 8.249164, 8.269558, 8.260358, 
    8.296317, 8.284944, 8.314884, 8.307737, 8.314548, 8.312482, 8.314574, 
    8.304095, 8.308583, 8.299372, 8.262079, 8.272549, 8.24136, 8.222613, 
    8.210183, 8.201373, 8.202619, 8.20499, 8.217202, 8.228711, 8.237476, 
    8.24333, 8.249104, 8.266593, 8.275877, 8.298298, 8.294534, 8.300916, 
    8.307027, 8.317293, 8.315602, 8.320128, 8.300751, 8.313621, 8.29239, 
    8.298188, 8.250659, 8.233253, 8.225821, 8.219336, 8.203575, 8.214454, 
    8.210162, 8.220381, 8.226879, 8.223665, 8.24349, 8.235793, 8.276428, 
    8.258901, 8.306314, 8.295306, 8.308956, 8.301988, 8.31393, 8.303182, 
    8.321815, 8.325876, 8.3231, 8.33378, 8.302586, 8.314545, 8.223574, 
    8.224098, 8.226542, 8.215806, 8.215151, 8.205335, 8.214069, 8.217792, 
    8.227258, 8.232861, 8.238171, 8.249855, 8.262922, 8.281239, 8.296019, 
    8.304891, 8.29945, 8.304254, 8.298883, 8.29637, 8.324353, 8.308622, 
    8.332243, 8.330935, 8.320234, 8.331082, 8.224466, 8.221451, 8.210986, 
    8.219174, 8.204267, 8.212605, 8.217402, 8.23595, 8.24002, 8.243791, 
    8.251248, 8.260828, 8.277658, 8.293928, 8.307384, 8.306397, 8.306744, 
    8.309752, 8.302301, 8.310976, 8.31243, 8.308624, 8.330759, 8.324428, 
    8.330907, 8.326784, 8.222431, 8.227509, 8.224764, 8.229924, 8.226287, 
    8.242431, 8.247268, 8.269949, 8.260638, 8.275469, 8.262145, 8.264503, 
    8.275945, 8.262865, 8.293112, 8.272074, 8.309869, 8.288775, 8.311093, 
    8.307325, 8.313567, 8.31916, 8.326206, 8.339222, 8.336206, 8.347111, 
    8.235079, 8.241646, 8.241071, 8.247952, 8.253044, 8.264096, 8.281856, 
    8.275171, 8.28745, 8.291496, 8.271267, 8.282708, 8.246047, 8.251955, 
    8.248439, 8.235595, 8.276707, 8.255579, 8.296237, 8.283165, 8.318361, 
    8.301611, 8.334546, 8.348664, 8.362003, 8.377599, 8.245236, 8.24077, 
    8.248772, 8.259851, 8.270148, 8.283865, 8.285272, 8.287844, 8.296102, 
    8.301723, 8.288653, 8.303133, 8.253319, 8.278545, 8.239079, 8.250938, 
    8.259198, 8.255577, 8.274409, 8.278855, 8.298539, 8.287592, 8.345173, 
    8.320334, 8.389516, 8.370105, 8.23921, 8.245222, 8.266179, 8.256203, 
    8.284783, 8.293419, 8.299169, 8.306521, 8.307319, 8.31168, 8.304534, 
    8.311399, 8.283894, 8.297042, 8.263785, 8.271476, 8.267938, 8.264057, 
    8.276043, 8.288834, 8.289113, 8.294803, 8.306388, 8.284899, 8.348371, 
    8.310061, 8.251783, 8.263381, 8.265044, 8.26055, 8.29271, 8.28003, 
    8.311574, 8.303459, 8.316763, 8.310148, 8.309175, 8.300693, 8.295417, 
    8.280538, 8.269743, 8.261201, 8.263187, 8.272574, 8.289618, 8.307387, 
    8.303836, 8.315751, 8.282706, 8.297451, 8.292354, 8.305655, 8.274992, 
    8.301307, 8.268686, 8.271402, 8.27981, 8.298342, 8.302111, 8.306127, 
    8.30365, 8.291632, 8.288091, 8.279607, 8.277264, 8.270811, 8.265472, 
    8.270349, 8.275474, 8.29164, 8.304826, 8.319239, 8.322772, 8.339642, 
    8.325895, 8.348583, 8.329273, 8.362744, 8.302753, 8.328723, 8.280195, 
    8.285233, 8.295933, 8.31693, 8.305593, 8.318857, 8.288014, 8.272896, 
    8.268997, 8.26172, 8.269163, 8.268558, 8.27569, 8.273397, 8.292126, 
    8.281328, 8.309149, 8.318753, 8.345964, 8.362698, 8.379789, 8.387344, 
    8.389647, 8.390608 ;

 FGR =
  -324.7462, -325.5064, -325.359, -325.9713, -325.6324, -326.0328, -324.9012, 
    -325.5359, -325.1311, -324.8158, -327.1569, -325.9988, -328.3655, 
    -327.6271, -329.4947, -328.2495, -329.744, -329.4608, -330.3177, 
    -330.0723, -331.1647, -330.431, -331.734, -330.9904, -331.1061, 
    -330.4065, -326.2337, -327.0121, -326.1871, -326.2982, -326.2488, 
    -325.6387, -325.3301, -324.6894, -324.806, -325.2773, -326.3482, 
    -325.986, -326.9025, -326.8818, -327.8999, -327.4412, -329.1626, 
    -328.6664, -330.0826, -329.7287, -330.0657, -329.9637, -330.067, 
    -329.548, -329.7703, -329.3142, -327.5268, -328.0486, -326.4899, 
    -325.549, -324.9286, -324.4871, -324.5495, -324.6682, -325.28, -325.857, 
    -326.2961, -326.5895, -326.8788, -327.7492, -328.2134, -329.2599, 
    -329.0744, -329.3899, -329.6935, -330.2013, -330.118, -330.3413, 
    -329.3827, -330.0192, -328.9684, -329.2556, -326.9513, -326.084, 
    -325.7099, -325.3871, -324.5974, -325.1424, -324.9274, -325.4403, 
    -325.7653, -325.6048, -326.5975, -326.2114, -328.2409, -327.3676, 
    -329.6581, -329.1126, -329.7891, -329.4442, -330.0347, -329.5033, 
    -330.4249, -330.6249, -330.4881, -331.0157, -329.4737, -330.0651, -325.6, 
    -325.6262, -325.7487, -325.2101, -325.1775, -324.6859, -325.1239, 
    -325.3099, -325.7847, -326.0644, -326.3305, -326.9159, -327.5682, 
    -328.481, -329.1479, -329.588, -329.3185, -329.5564, -329.2903, 
    -329.1658, -330.5496, -329.772, -330.9398, -330.8754, -330.3463, 
    -330.8827, -325.6446, -325.494, -324.9691, -325.3799, -324.6324, -325.05, 
    -325.2897, -326.2181, -326.4235, -326.6121, -326.9859, -327.4647, 
    -328.303, -329.0436, -329.7115, -329.6627, -329.6798, -329.8284, 
    -329.4595, -329.889, -329.9605, -329.7726, -330.8668, -330.5542, 
    -330.874, -330.6707, -325.5431, -325.7968, -325.6596, -325.9173, 
    -325.7353, -326.5427, -326.7847, -327.9181, -327.4549, -328.1938, 
    -327.5305, -327.6477, -328.2152, -327.5667, -329.0022, -328.0234, 
    -329.8342, -328.854, -329.8948, -329.7086, -330.0175, -330.2935, 
    -330.6419, -331.2831, -331.1349, -331.6721, -326.1757, -326.5041, 
    -326.4763, -326.8209, -327.0754, -327.6281, -328.5123, -328.1801, 
    -328.7911, -328.9236, -327.9858, -328.5543, -326.7248, -327.0195, 
    -326.8449, -326.2009, -328.2551, -327.201, -329.1585, -328.5777, 
    -330.254, -329.4241, -331.053, -331.7466, -332.4048, -333.1678, 
    -326.6846, -326.4613, -326.8622, -327.4145, -327.9295, -328.6123, 
    -328.6828, -328.8103, -329.1524, -329.431, -328.8495, -329.5009, 
    -327.0855, -328.3471, -326.3758, -326.9684, -327.3825, -327.2021, 
    -328.1425, -328.3636, -329.2722, -328.7982, -331.5744, -330.3502, 
    -333.7527, -332.8008, -326.383, -326.6844, -327.7309, -327.2336, 
    -328.6585, -329.0189, -329.3046, -329.668, -329.7081, -329.9236, 
    -329.5703, -329.9101, -328.6137, -329.1988, -327.6128, -327.9956, 
    -327.8199, -327.6263, -328.2237, -328.8582, -328.8737, -329.087, 
    -329.6564, -328.6643, -331.729, -329.839, -327.0129, -327.5905, 
    -327.6751, -327.4512, -328.9837, -328.4217, -329.9186, -329.5171, 
    -330.1754, -329.8481, -329.7999, -329.3799, -329.118, -328.4466, 
    -327.9091, -327.4839, -327.5829, -328.0501, -328.8975, -329.7109, 
    -329.5347, -330.1254, -328.5551, -329.2184, -328.9653, -329.6256, 
    -328.1709, -329.4055, -327.8573, -327.9925, -328.4107, -329.2615, 
    -329.4502, -329.6484, -329.5265, -328.9295, -328.8224, -328.401, 
    -328.2838, -327.9632, -327.697, -327.9398, -328.1944, -328.9306, 
    -329.584, -330.2972, -330.4724, -331.3013, -330.624, -331.7391, 
    -330.7872, -332.4371, -329.4792, -330.763, -328.4304, -328.6809, 
    -329.1424, -330.1817, -329.6225, -330.2773, -328.8188, -328.0653, 
    -327.8727, -327.5094, -327.881, -327.8508, -328.2062, -328.0921, 
    -328.9547, -328.4868, -329.7982, -330.2726, -331.6152, -332.4372, 
    -333.2771, -333.6469, -333.7597, -333.8067 ;

 FGR12 =
  -224.3387, -224.3013, -224.3084, -224.2788, -224.2949, -224.2757, 
    -224.3307, -224.3001, -224.3194, -224.3348, -224.2226, -224.2774, 
    -224.1649, -224.1989, -224.1143, -224.1707, -224.1029, -224.1153, 
    -224.0764, -224.0875, -224.0399, -224.0714, -224.0145, -224.047, 
    -224.0421, -224.0726, -224.2655, -224.2295, -224.2679, -224.2626, 
    -224.2648, -224.2948, -224.3104, -224.341, -224.3353, -224.3125, 
    -224.2602, -224.2776, -224.2328, -224.2337, -224.1861, -224.2075, 
    -224.1289, -224.1503, -224.087, -224.1031, -224.0879, -224.0924, 
    -224.0878, -224.1114, -224.1013, -224.1219, -224.2036, -224.1792, 
    -224.2531, -224.3001, -224.3295, -224.3511, -224.3481, -224.3424, 
    -224.3124, -224.284, -224.2623, -224.2479, -224.2339, -224.1942, 
    -224.172, -224.1248, -224.1328, -224.1188, -224.1046, -224.0818, 
    -224.0855, -224.0756, -224.1187, -224.0902, -224.1375, -224.1246, 
    -224.2325, -224.2728, -224.2921, -224.3071, -224.3458, -224.3191, 
    -224.3297, -224.3041, -224.2884, -224.2961, -224.2475, -224.2665, 
    -224.1707, -224.2113, -224.1062, -224.1311, -224.1003, -224.1159, 
    -224.0894, -224.1132, -224.0718, -224.0632, -224.0691, -224.0455, 
    -224.1146, -224.0881, -224.2964, -224.2952, -224.2891, -224.3159, 
    -224.3173, -224.3413, -224.3198, -224.3108, -224.2873, -224.2738, 
    -224.2608, -224.2323, -224.2019, -224.1593, -224.1295, -224.1093, 
    -224.1215, -224.1108, -224.1229, -224.1285, -224.0665, -224.1014, 
    -224.0489, -224.0517, -224.0755, -224.0513, -224.2943, -224.3015, 
    -224.3274, -224.3071, -224.3439, -224.3235, -224.3121, -224.2666, 
    -224.2561, -224.247, -224.2289, -224.2064, -224.1675, -224.1344, 
    -224.1037, -224.1059, -224.1052, -224.0986, -224.1153, -224.0958, 
    -224.0928, -224.1011, -224.052, -224.0659, -224.0517, -224.0607, 
    -224.2991, -224.2869, -224.2935, -224.2812, -224.2901, -224.2508, 
    -224.2392, -224.1857, -224.207, -224.1726, -224.2032, -224.1979, 
    -224.1725, -224.2014, -224.1367, -224.1811, -224.0983, -224.1429, 
    -224.0956, -224.1039, -224.0899, -224.0777, -224.0621, -224.0341, 
    -224.0405, -224.0169, -224.2683, -224.2525, -224.2534, -224.2367, 
    -224.2248, -224.1986, -224.1576, -224.1728, -224.1445, -224.1397, 
    -224.1818, -224.1558, -224.2417, -224.228, -224.2357, -224.2673, 
    -224.1699, -224.2194, -224.1291, -224.1545, -224.0795, -224.1174, 
    -224.0441, -224.0145, -223.985, -223.9533, -224.2434, -224.2542, 
    -224.2347, -224.2092, -224.1846, -224.1529, -224.1495, -224.1437, 
    -224.1291, -224.1165, -224.1424, -224.1132, -224.2258, -224.1654, 
    -224.2587, -224.2305, -224.2105, -224.2188, -224.1744, -224.1642, 
    -224.1241, -224.1441, -224.0222, -224.0758, -223.928, -223.9687, 
    -224.258, -224.2433, -224.1942, -224.2173, -224.1506, -224.1354, 
    -224.1221, -224.106, -224.1039, -224.0944, -224.1101, -224.0948, 
    -224.1529, -224.1271, -224.1992, -224.1815, -224.1895, -224.1986, 
    -224.1707, -224.142, -224.1407, -224.1325, -224.1086, -224.1504, 
    -224.0166, -224.1001, -224.2276, -224.2011, -224.1965, -224.2068, 
    -224.137, -224.1617, -224.0945, -224.1125, -224.0828, -224.0976, 
    -224.0998, -224.1188, -224.1308, -224.1607, -224.1856, -224.2052, 
    -224.2006, -224.1791, -224.1402, -224.104, -224.1122, -224.0851, 
    -224.1555, -224.1265, -224.1382, -224.1077, -224.1734, -224.1196, 
    -224.1877, -224.1815, -224.1622, -224.125, -224.1156, -224.1069, 
    -224.1121, -224.1398, -224.1433, -224.1625, -224.1682, -224.1828, 
    -224.1953, -224.184, -224.1725, -224.1395, -224.1099, -224.0776, 
    -224.0696, -224.0344, -224.064, -224.0163, -224.0584, -223.9854, 
    -224.1155, -224.058, -224.1611, -224.1495, -224.1303, -224.0834, 
    -224.1079, -224.0789, -224.1434, -224.1788, -224.1871, -224.2042, 
    -224.1867, -224.1881, -224.1715, -224.1767, -224.1384, -224.1585, 
    -224.1001, -224.079, -224.0196, -223.9843, -223.9478, -223.9322, 
    -223.9274, -223.9255 ;

 FGR_R =
  -324.7462, -325.5064, -325.359, -325.9713, -325.6324, -326.0328, -324.9012, 
    -325.5359, -325.1311, -324.8158, -327.1569, -325.9988, -328.3655, 
    -327.6271, -329.4947, -328.2495, -329.744, -329.4608, -330.3177, 
    -330.0723, -331.1647, -330.431, -331.734, -330.9904, -331.1061, 
    -330.4065, -326.2337, -327.0121, -326.1871, -326.2982, -326.2488, 
    -325.6387, -325.3301, -324.6894, -324.806, -325.2773, -326.3482, 
    -325.986, -326.9025, -326.8818, -327.8999, -327.4412, -329.1626, 
    -328.6664, -330.0826, -329.7287, -330.0657, -329.9637, -330.067, 
    -329.548, -329.7703, -329.3142, -327.5268, -328.0486, -326.4899, 
    -325.549, -324.9286, -324.4871, -324.5495, -324.6682, -325.28, -325.857, 
    -326.2961, -326.5895, -326.8788, -327.7492, -328.2134, -329.2599, 
    -329.0744, -329.3899, -329.6935, -330.2013, -330.118, -330.3413, 
    -329.3827, -330.0192, -328.9684, -329.2556, -326.9513, -326.084, 
    -325.7099, -325.3871, -324.5974, -325.1424, -324.9274, -325.4403, 
    -325.7653, -325.6048, -326.5975, -326.2114, -328.2409, -327.3676, 
    -329.6581, -329.1126, -329.7891, -329.4442, -330.0347, -329.5033, 
    -330.4249, -330.6249, -330.4881, -331.0157, -329.4737, -330.0651, -325.6, 
    -325.6262, -325.7487, -325.2101, -325.1775, -324.6859, -325.1239, 
    -325.3099, -325.7847, -326.0644, -326.3305, -326.9159, -327.5682, 
    -328.481, -329.1479, -329.588, -329.3185, -329.5564, -329.2903, 
    -329.1658, -330.5496, -329.772, -330.9398, -330.8754, -330.3463, 
    -330.8827, -325.6446, -325.494, -324.9691, -325.3799, -324.6324, -325.05, 
    -325.2897, -326.2181, -326.4235, -326.6121, -326.9859, -327.4647, 
    -328.303, -329.0436, -329.7115, -329.6627, -329.6798, -329.8284, 
    -329.4595, -329.889, -329.9605, -329.7726, -330.8668, -330.5542, 
    -330.874, -330.6707, -325.5431, -325.7968, -325.6596, -325.9173, 
    -325.7353, -326.5427, -326.7847, -327.9181, -327.4549, -328.1938, 
    -327.5305, -327.6477, -328.2152, -327.5667, -329.0022, -328.0234, 
    -329.8342, -328.854, -329.8948, -329.7086, -330.0175, -330.2935, 
    -330.6419, -331.2831, -331.1349, -331.6721, -326.1757, -326.5041, 
    -326.4763, -326.8209, -327.0754, -327.6281, -328.5123, -328.1801, 
    -328.7911, -328.9236, -327.9858, -328.5543, -326.7248, -327.0195, 
    -326.8449, -326.2009, -328.2551, -327.201, -329.1585, -328.5777, 
    -330.254, -329.4241, -331.053, -331.7466, -332.4048, -333.1678, 
    -326.6846, -326.4613, -326.8622, -327.4145, -327.9295, -328.6123, 
    -328.6828, -328.8103, -329.1524, -329.431, -328.8495, -329.5009, 
    -327.0855, -328.3471, -326.3758, -326.9684, -327.3825, -327.2021, 
    -328.1425, -328.3636, -329.2722, -328.7982, -331.5744, -330.3502, 
    -333.7527, -332.8008, -326.383, -326.6844, -327.7309, -327.2336, 
    -328.6585, -329.0189, -329.3046, -329.668, -329.7081, -329.9236, 
    -329.5703, -329.9101, -328.6137, -329.1988, -327.6128, -327.9956, 
    -327.8199, -327.6263, -328.2237, -328.8582, -328.8737, -329.087, 
    -329.6564, -328.6643, -331.729, -329.839, -327.0129, -327.5905, 
    -327.6751, -327.4512, -328.9837, -328.4217, -329.9186, -329.5171, 
    -330.1754, -329.8481, -329.7999, -329.3799, -329.118, -328.4466, 
    -327.9091, -327.4839, -327.5829, -328.0501, -328.8975, -329.7109, 
    -329.5347, -330.1254, -328.5551, -329.2184, -328.9653, -329.6256, 
    -328.1709, -329.4055, -327.8573, -327.9925, -328.4107, -329.2615, 
    -329.4502, -329.6484, -329.5265, -328.9295, -328.8224, -328.401, 
    -328.2838, -327.9632, -327.697, -327.9398, -328.1944, -328.9306, 
    -329.584, -330.2972, -330.4724, -331.3013, -330.624, -331.7391, 
    -330.7872, -332.4371, -329.4792, -330.763, -328.4304, -328.6809, 
    -329.1424, -330.1817, -329.6225, -330.2773, -328.8188, -328.0653, 
    -327.8727, -327.5094, -327.881, -327.8508, -328.2062, -328.0921, 
    -328.9547, -328.4868, -329.7982, -330.2726, -331.6152, -332.4372, 
    -333.2771, -333.6469, -333.7597, -333.8067 ;

 FGR_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FIRA =
  74.69257, 74.7455, 74.73524, 74.77787, 74.75427, 74.78214, 74.70335, 
    74.74755, 74.71938, 74.69741, 74.86048, 74.77979, 74.94505, 74.89335, 
    75.02299, 74.93693, 75.04046, 75.02063, 75.08063, 75.06345, 75.13989, 
    75.08855, 75.17974, 75.12771, 75.1358, 75.08684, 74.79614, 74.8504, 
    74.7929, 74.80064, 74.7972, 74.75471, 74.73322, 74.68861, 74.69673, 
    74.72955, 74.80413, 74.77888, 74.84276, 74.84132, 74.91246, 74.88035, 
    74.99975, 74.96613, 75.06416, 75.03938, 75.06298, 75.05584, 75.06307, 
    75.02673, 75.0423, 75.01037, 74.88633, 74.92286, 74.814, 74.74847, 
    74.70527, 74.67452, 74.67886, 74.68713, 74.72974, 74.76991, 74.8005, 
    74.82095, 74.84111, 74.90189, 74.9344, 75.00656, 74.99358, 75.01566, 
    75.03693, 75.07247, 75.06664, 75.08227, 75.01516, 75.05972, 74.98615, 
    75.00626, 74.84615, 74.78571, 74.75967, 74.7372, 74.6822, 74.72015, 
    74.70518, 74.7409, 74.76353, 74.75235, 74.8215, 74.79459, 74.93633, 
    74.87519, 75.03445, 74.99625, 75.04362, 75.01947, 75.06081, 75.02361, 
    75.08813, 75.10212, 75.09254, 75.12948, 75.02153, 75.06293, 74.75202, 
    74.75384, 74.76237, 74.72487, 74.7226, 74.68836, 74.71886, 74.73182, 
    74.76487, 74.78434, 74.80289, 74.84369, 74.88922, 74.95314, 74.99872, 
    75.02953, 75.01067, 75.02732, 75.00869, 74.99998, 75.09685, 75.04241, 
    75.12417, 75.11966, 75.08263, 75.12017, 74.75513, 74.74464, 74.70809, 
    74.73669, 74.68464, 74.71372, 74.73041, 74.79506, 74.80938, 74.82252, 
    74.84858, 74.88199, 74.94068, 74.99142, 75.03819, 75.03477, 75.03596, 
    75.04636, 75.02054, 75.05061, 75.05561, 75.04247, 75.11906, 75.09718, 
    75.11956, 75.10533, 74.74805, 74.76572, 74.75617, 74.77411, 74.76144, 
    74.81768, 74.83455, 74.91373, 74.8813, 74.93303, 74.88659, 74.89479, 
    74.93452, 74.88913, 74.98851, 74.9211, 75.04677, 74.97926, 75.05102, 
    75.03798, 75.05961, 75.07893, 75.10332, 75.14819, 75.13782, 75.17542, 
    74.7921, 74.81499, 74.81306, 74.83707, 74.85481, 74.89342, 74.95534, 
    74.93208, 74.97488, 74.98301, 74.91847, 74.95827, 74.83038, 74.85091, 
    74.83875, 74.79385, 74.93732, 74.86356, 74.99947, 74.95992, 75.07616, 
    75.01805, 75.13209, 75.18061, 75.22667, 75.28004, 74.82758, 74.81201, 
    74.83995, 74.87847, 74.91453, 74.96234, 74.96728, 74.97622, 74.99904, 
    75.01854, 74.97896, 75.02344, 74.85551, 74.94376, 74.80605, 74.84735, 
    74.87624, 74.86364, 74.92944, 74.94493, 75.00742, 74.97537, 75.16856, 
    75.08289, 75.32095, 75.25437, 74.80655, 74.82756, 74.90062, 74.86583, 
    74.96558, 74.98968, 75.00969, 75.03513, 75.03794, 75.05303, 75.0283, 
    75.05209, 74.96244, 75.00228, 74.89235, 74.91916, 74.90686, 74.8933, 
    74.93513, 74.97957, 74.98065, 74.99445, 75.0343, 74.96599, 75.17937, 
    75.04709, 74.85046, 74.89078, 74.89671, 74.88104, 74.98722, 74.94899, 
    75.05268, 75.02457, 75.07066, 75.04774, 75.04437, 75.01497, 74.99663, 
    74.95074, 74.9131, 74.88333, 74.89026, 74.92297, 74.98232, 75.03814, 
    75.02579, 75.06716, 74.95834, 75.00365, 74.98593, 75.03217, 74.93143, 
    75.01674, 74.90948, 74.91895, 74.94823, 75.00667, 75.01989, 75.03377, 
    75.02523, 74.98342, 74.97706, 74.94755, 74.93933, 74.91689, 74.89825, 
    74.91525, 74.93307, 74.9835, 75.02925, 75.07919, 75.09145, 75.14945, 
    75.10205, 75.18008, 75.11346, 75.22892, 75.0219, 75.11178, 74.9496, 
    74.96716, 74.99833, 75.07109, 75.03195, 75.07779, 74.97681, 74.92403, 
    74.91055, 74.88512, 74.91113, 74.90902, 74.93391, 74.92592, 74.98519, 
    74.95354, 75.04425, 75.07746, 75.17142, 75.22894, 75.28769, 75.31355, 
    75.32144, 75.32473 ;

 FIRA_R =
  74.69257, 74.7455, 74.73524, 74.77787, 74.75427, 74.78214, 74.70335, 
    74.74755, 74.71938, 74.69741, 74.86048, 74.77979, 74.94505, 74.89335, 
    75.02299, 74.93693, 75.04046, 75.02063, 75.08063, 75.06345, 75.13989, 
    75.08855, 75.17974, 75.12771, 75.1358, 75.08684, 74.79614, 74.8504, 
    74.7929, 74.80064, 74.7972, 74.75471, 74.73322, 74.68861, 74.69673, 
    74.72955, 74.80413, 74.77888, 74.84276, 74.84132, 74.91246, 74.88035, 
    74.99975, 74.96613, 75.06416, 75.03938, 75.06298, 75.05584, 75.06307, 
    75.02673, 75.0423, 75.01037, 74.88633, 74.92286, 74.814, 74.74847, 
    74.70527, 74.67452, 74.67886, 74.68713, 74.72974, 74.76991, 74.8005, 
    74.82095, 74.84111, 74.90189, 74.9344, 75.00656, 74.99358, 75.01566, 
    75.03693, 75.07247, 75.06664, 75.08227, 75.01516, 75.05972, 74.98615, 
    75.00626, 74.84615, 74.78571, 74.75967, 74.7372, 74.6822, 74.72015, 
    74.70518, 74.7409, 74.76353, 74.75235, 74.8215, 74.79459, 74.93633, 
    74.87519, 75.03445, 74.99625, 75.04362, 75.01947, 75.06081, 75.02361, 
    75.08813, 75.10212, 75.09254, 75.12948, 75.02153, 75.06293, 74.75202, 
    74.75384, 74.76237, 74.72487, 74.7226, 74.68836, 74.71886, 74.73182, 
    74.76487, 74.78434, 74.80289, 74.84369, 74.88922, 74.95314, 74.99872, 
    75.02953, 75.01067, 75.02732, 75.00869, 74.99998, 75.09685, 75.04241, 
    75.12417, 75.11966, 75.08263, 75.12017, 74.75513, 74.74464, 74.70809, 
    74.73669, 74.68464, 74.71372, 74.73041, 74.79506, 74.80938, 74.82252, 
    74.84858, 74.88199, 74.94068, 74.99142, 75.03819, 75.03477, 75.03596, 
    75.04636, 75.02054, 75.05061, 75.05561, 75.04247, 75.11906, 75.09718, 
    75.11956, 75.10533, 74.74805, 74.76572, 74.75617, 74.77411, 74.76144, 
    74.81768, 74.83455, 74.91373, 74.8813, 74.93303, 74.88659, 74.89479, 
    74.93452, 74.88913, 74.98851, 74.9211, 75.04677, 74.97926, 75.05102, 
    75.03798, 75.05961, 75.07893, 75.10332, 75.14819, 75.13782, 75.17542, 
    74.7921, 74.81499, 74.81306, 74.83707, 74.85481, 74.89342, 74.95534, 
    74.93208, 74.97488, 74.98301, 74.91847, 74.95827, 74.83038, 74.85091, 
    74.83875, 74.79385, 74.93732, 74.86356, 74.99947, 74.95992, 75.07616, 
    75.01805, 75.13209, 75.18061, 75.22667, 75.28004, 74.82758, 74.81201, 
    74.83995, 74.87847, 74.91453, 74.96234, 74.96728, 74.97622, 74.99904, 
    75.01854, 74.97896, 75.02344, 74.85551, 74.94376, 74.80605, 74.84735, 
    74.87624, 74.86364, 74.92944, 74.94493, 75.00742, 74.97537, 75.16856, 
    75.08289, 75.32095, 75.25437, 74.80655, 74.82756, 74.90062, 74.86583, 
    74.96558, 74.98968, 75.00969, 75.03513, 75.03794, 75.05303, 75.0283, 
    75.05209, 74.96244, 75.00228, 74.89235, 74.91916, 74.90686, 74.8933, 
    74.93513, 74.97957, 74.98065, 74.99445, 75.0343, 74.96599, 75.17937, 
    75.04709, 74.85046, 74.89078, 74.89671, 74.88104, 74.98722, 74.94899, 
    75.05268, 75.02457, 75.07066, 75.04774, 75.04437, 75.01497, 74.99663, 
    74.95074, 74.9131, 74.88333, 74.89026, 74.92297, 74.98232, 75.03814, 
    75.02579, 75.06716, 74.95834, 75.00365, 74.98593, 75.03217, 74.93143, 
    75.01674, 74.90948, 74.91895, 74.94823, 75.00667, 75.01989, 75.03377, 
    75.02523, 74.98342, 74.97706, 74.94755, 74.93933, 74.91689, 74.89825, 
    74.91525, 74.93307, 74.9835, 75.02925, 75.07919, 75.09145, 75.14945, 
    75.10205, 75.18008, 75.11346, 75.22892, 75.0219, 75.11178, 74.9496, 
    74.96716, 74.99833, 75.07109, 75.03195, 75.07779, 74.97681, 74.92403, 
    74.91055, 74.88512, 74.91113, 74.90902, 74.93391, 74.92592, 74.98519, 
    74.95354, 75.04425, 75.07746, 75.17142, 75.22894, 75.28769, 75.31355, 
    75.32144, 75.32473 ;

 FIRA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FIRE =
  263.6535, 263.7065, 263.6962, 263.7388, 263.7152, 263.7431, 263.6643, 
    263.7085, 263.6803, 263.6584, 263.8214, 263.7407, 263.906, 263.8543, 
    263.9839, 263.8979, 264.0014, 263.9816, 264.0416, 264.0244, 264.1008, 
    264.0495, 264.1407, 264.0887, 264.0967, 264.0478, 263.7571, 263.8113, 
    263.7538, 263.7616, 263.7581, 263.7156, 263.6942, 263.6495, 263.6577, 
    263.6905, 263.7651, 263.7398, 263.8037, 263.8022, 263.8734, 263.8413, 
    263.9607, 263.9271, 264.0251, 264.0003, 264.0239, 264.0168, 264.024, 
    263.9877, 264.0032, 263.9713, 263.8473, 263.8838, 263.7749, 263.7094, 
    263.6662, 263.6355, 263.6398, 263.6481, 263.6907, 263.7308, 263.7614, 
    263.7819, 263.8021, 263.8628, 263.8953, 263.9675, 263.9545, 263.9766, 
    263.9979, 264.0334, 264.0276, 264.0432, 263.9761, 264.0207, 263.9471, 
    263.9672, 263.8071, 263.7466, 263.7206, 263.6982, 263.6431, 263.6811, 
    263.6661, 263.7018, 263.7245, 263.7133, 263.7824, 263.7555, 263.8973, 
    263.8361, 263.9954, 263.9572, 264.0045, 263.9804, 264.0218, 263.9846, 
    264.0491, 264.063, 264.0535, 264.0904, 263.9825, 264.0239, 263.713, 
    263.7148, 263.7233, 263.6858, 263.6835, 263.6493, 263.6798, 263.6927, 
    263.7258, 263.7453, 263.7638, 263.8046, 263.8502, 263.9141, 263.9597, 
    263.9905, 263.9716, 263.9883, 263.9696, 263.9609, 264.0578, 264.0034, 
    264.0851, 264.0806, 264.0435, 264.0811, 263.7161, 263.7056, 263.669, 
    263.6976, 263.6456, 263.6747, 263.6913, 263.756, 263.7703, 263.7834, 
    263.8095, 263.8429, 263.9016, 263.9524, 263.9991, 263.9957, 263.9969, 
    264.0073, 263.9815, 264.0115, 264.0165, 264.0034, 264.08, 264.0581, 
    264.0805, 264.0663, 263.709, 263.7267, 263.7171, 263.735, 263.7224, 
    263.7786, 263.7955, 263.8747, 263.8423, 263.894, 263.8475, 263.8557, 
    263.8955, 263.8501, 263.9494, 263.882, 264.0077, 263.9402, 264.012, 
    263.9989, 264.0205, 264.0399, 264.0643, 264.1091, 264.0988, 264.1364, 
    263.7531, 263.7759, 263.774, 263.798, 263.8158, 263.8544, 263.9163, 
    263.893, 263.9358, 263.9439, 263.8794, 263.9192, 263.7913, 263.8119, 
    263.7997, 263.7548, 263.8983, 263.8245, 263.9604, 263.9209, 264.0371, 
    263.979, 264.093, 264.1415, 264.1876, 264.241, 263.7885, 263.7729, 
    263.8009, 263.8394, 263.8755, 263.9233, 263.9282, 263.9372, 263.96, 
    263.9795, 263.9399, 263.9844, 263.8164, 263.9047, 263.767, 263.8083, 
    263.8372, 263.8246, 263.8904, 263.9059, 263.9684, 263.9363, 264.1295, 
    264.0438, 264.2819, 264.2153, 263.7675, 263.7885, 263.8615, 263.8268, 
    263.9265, 263.9506, 263.9706, 263.9961, 263.9989, 264.014, 263.9892, 
    264.013, 263.9234, 263.9632, 263.8533, 263.8801, 263.8678, 263.8542, 
    263.8961, 263.9405, 263.9416, 263.9554, 263.9952, 263.9269, 264.1403, 
    264.008, 263.8114, 263.8517, 263.8576, 263.842, 263.9482, 263.9099, 
    264.0136, 263.9855, 264.0316, 264.0087, 264.0053, 263.9759, 263.9576, 
    263.9117, 263.8741, 263.8443, 263.8512, 263.8839, 263.9433, 263.9991, 
    263.9867, 264.0281, 263.9193, 263.9646, 263.9469, 263.9931, 263.8924, 
    263.9777, 263.8704, 263.8799, 263.9091, 263.9676, 263.9808, 263.9947, 
    263.9862, 263.9444, 263.938, 263.9085, 263.9003, 263.8778, 263.8592, 
    263.8762, 263.894, 263.9444, 263.9902, 264.0401, 264.0524, 264.1104, 
    264.063, 264.141, 264.0744, 264.1898, 263.9828, 264.0727, 263.9106, 
    263.9281, 263.9593, 264.032, 263.9929, 264.0387, 263.9377, 263.885, 
    263.8715, 263.8461, 263.8721, 263.87, 263.8948, 263.8868, 263.9461, 
    263.9145, 264.0052, 264.0384, 264.1324, 264.1899, 264.2486, 264.2745, 
    264.2824, 264.2857 ;

 FIRE_R =
  263.6535, 263.7065, 263.6962, 263.7388, 263.7152, 263.7431, 263.6643, 
    263.7085, 263.6803, 263.6584, 263.8214, 263.7407, 263.906, 263.8543, 
    263.9839, 263.8979, 264.0014, 263.9816, 264.0416, 264.0244, 264.1008, 
    264.0495, 264.1407, 264.0887, 264.0967, 264.0478, 263.7571, 263.8113, 
    263.7538, 263.7616, 263.7581, 263.7156, 263.6942, 263.6495, 263.6577, 
    263.6905, 263.7651, 263.7398, 263.8037, 263.8022, 263.8734, 263.8413, 
    263.9607, 263.9271, 264.0251, 264.0003, 264.0239, 264.0168, 264.024, 
    263.9877, 264.0032, 263.9713, 263.8473, 263.8838, 263.7749, 263.7094, 
    263.6662, 263.6355, 263.6398, 263.6481, 263.6907, 263.7308, 263.7614, 
    263.7819, 263.8021, 263.8628, 263.8953, 263.9675, 263.9545, 263.9766, 
    263.9979, 264.0334, 264.0276, 264.0432, 263.9761, 264.0207, 263.9471, 
    263.9672, 263.8071, 263.7466, 263.7206, 263.6982, 263.6431, 263.6811, 
    263.6661, 263.7018, 263.7245, 263.7133, 263.7824, 263.7555, 263.8973, 
    263.8361, 263.9954, 263.9572, 264.0045, 263.9804, 264.0218, 263.9846, 
    264.0491, 264.063, 264.0535, 264.0904, 263.9825, 264.0239, 263.713, 
    263.7148, 263.7233, 263.6858, 263.6835, 263.6493, 263.6798, 263.6927, 
    263.7258, 263.7453, 263.7638, 263.8046, 263.8502, 263.9141, 263.9597, 
    263.9905, 263.9716, 263.9883, 263.9696, 263.9609, 264.0578, 264.0034, 
    264.0851, 264.0806, 264.0435, 264.0811, 263.7161, 263.7056, 263.669, 
    263.6976, 263.6456, 263.6747, 263.6913, 263.756, 263.7703, 263.7834, 
    263.8095, 263.8429, 263.9016, 263.9524, 263.9991, 263.9957, 263.9969, 
    264.0073, 263.9815, 264.0115, 264.0165, 264.0034, 264.08, 264.0581, 
    264.0805, 264.0663, 263.709, 263.7267, 263.7171, 263.735, 263.7224, 
    263.7786, 263.7955, 263.8747, 263.8423, 263.894, 263.8475, 263.8557, 
    263.8955, 263.8501, 263.9494, 263.882, 264.0077, 263.9402, 264.012, 
    263.9989, 264.0205, 264.0399, 264.0643, 264.1091, 264.0988, 264.1364, 
    263.7531, 263.7759, 263.774, 263.798, 263.8158, 263.8544, 263.9163, 
    263.893, 263.9358, 263.9439, 263.8794, 263.9192, 263.7913, 263.8119, 
    263.7997, 263.7548, 263.8983, 263.8245, 263.9604, 263.9209, 264.0371, 
    263.979, 264.093, 264.1415, 264.1876, 264.241, 263.7885, 263.7729, 
    263.8009, 263.8394, 263.8755, 263.9233, 263.9282, 263.9372, 263.96, 
    263.9795, 263.9399, 263.9844, 263.8164, 263.9047, 263.767, 263.8083, 
    263.8372, 263.8246, 263.8904, 263.9059, 263.9684, 263.9363, 264.1295, 
    264.0438, 264.2819, 264.2153, 263.7675, 263.7885, 263.8615, 263.8268, 
    263.9265, 263.9506, 263.9706, 263.9961, 263.9989, 264.014, 263.9892, 
    264.013, 263.9234, 263.9632, 263.8533, 263.8801, 263.8678, 263.8542, 
    263.8961, 263.9405, 263.9416, 263.9554, 263.9952, 263.9269, 264.1403, 
    264.008, 263.8114, 263.8517, 263.8576, 263.842, 263.9482, 263.9099, 
    264.0136, 263.9855, 264.0316, 264.0087, 264.0053, 263.9759, 263.9576, 
    263.9117, 263.8741, 263.8443, 263.8512, 263.8839, 263.9433, 263.9991, 
    263.9867, 264.0281, 263.9193, 263.9646, 263.9469, 263.9931, 263.8924, 
    263.9777, 263.8704, 263.8799, 263.9091, 263.9676, 263.9808, 263.9947, 
    263.9862, 263.9444, 263.938, 263.9085, 263.9003, 263.8778, 263.8592, 
    263.8762, 263.894, 263.9444, 263.9902, 264.0401, 264.0524, 264.1104, 
    264.063, 264.141, 264.0744, 264.1898, 263.9828, 264.0727, 263.9106, 
    263.9281, 263.9593, 264.032, 263.9929, 264.0387, 263.9377, 263.885, 
    263.8715, 263.8461, 263.8721, 263.87, 263.8948, 263.8868, 263.9461, 
    263.9145, 264.0052, 264.0384, 264.1324, 264.1899, 264.2486, 264.2745, 
    264.2824, 264.2857 ;

 FIRE_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FLDS =
  188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 188.9609, 
    188.9609, 188.9609 ;

 FPG =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI_vr =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WJ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROST_TABLE =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 FSA =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSAT =
  0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584 ;

 FSA_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSDS =
  1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658 ;

 FSDSND =
  0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004 ;

 FSDSNDLN =
  0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372 ;

 FSDSNI =
  0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284 ;

 FSDSVD =
  0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081 ;

 FSDSVDLN =
  0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678 ;

 FSDSVI =
  0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228 ;

 FSDSVILN =
  0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 0.7125012, 
    0.7125012, 0.7125012 ;

 FSH =
  243.7966, 244.4876, 244.3536, 244.9102, 244.6021, 244.966, 243.9374, 
    244.5144, 244.1465, 243.8598, 245.9876, 244.9352, 247.0857, 246.4149, 
    248.1112, 246.9804, 248.3377, 248.0805, 248.8588, 248.6359, 249.6281, 
    248.9617, 250.1451, 249.4698, 249.5748, 248.9394, 245.1486, 245.8561, 
    245.1063, 245.2073, 245.1624, 244.6078, 244.3273, 243.7449, 243.851, 
    244.2793, 245.2527, 244.9235, 245.7565, 245.7377, 246.6628, 246.2461, 
    247.8095, 247.3591, 248.6452, 248.3238, 248.6298, 248.5372, 248.6311, 
    248.1597, 248.3615, 247.9473, 246.3238, 246.7978, 245.3815, 244.5263, 
    243.9624, 243.5611, 243.6178, 243.7256, 244.2818, 244.8062, 245.2054, 
    245.472, 245.735, 246.5259, 246.9475, 247.898, 247.7295, 248.0161, 
    248.2919, 248.753, 248.6773, 248.8802, 248.0095, 248.5876, 247.6331, 
    247.894, 245.8008, 245.0126, 244.6725, 244.3792, 243.6613, 244.1567, 
    243.9613, 244.4275, 244.7229, 244.577, 245.4793, 245.1284, 246.9725, 
    246.1792, 248.2597, 247.7642, 248.3787, 248.0654, 248.6017, 248.119, 
    248.9561, 249.1378, 249.0135, 249.4928, 248.0921, 248.6293, 244.5727, 
    244.5964, 244.7078, 244.2182, 244.1886, 243.7417, 244.1399, 244.309, 
    244.7405, 244.9947, 245.2366, 245.7686, 246.3614, 247.1906, 247.7962, 
    248.196, 247.9512, 248.1673, 247.9255, 247.8125, 249.0694, 248.3631, 
    249.4238, 249.3653, 248.8848, 249.3719, 244.6132, 244.4763, 243.9992, 
    244.3726, 243.6932, 244.0727, 244.2906, 245.1345, 245.3212, 245.4925, 
    245.8323, 246.2674, 247.029, 247.7015, 248.3081, 248.2638, 248.2793, 
    248.4143, 248.0793, 248.4694, 248.5343, 248.3637, 249.3574, 249.0736, 
    249.3641, 249.1794, 244.521, 244.7516, 244.6269, 244.8611, 244.6956, 
    245.4295, 245.6494, 246.6793, 246.2585, 246.9297, 246.3271, 246.4336, 
    246.9492, 246.3601, 247.6639, 246.7749, 248.4196, 247.5294, 248.4746, 
    248.3055, 248.5861, 248.8368, 249.1533, 249.7356, 249.601, 250.0889, 
    245.0959, 245.3944, 245.3691, 245.6823, 245.9136, 246.4158, 247.2191, 
    246.9173, 247.4724, 247.5925, 246.7408, 247.2572, 245.5949, 245.8628, 
    245.7041, 245.1188, 246.9854, 246.0277, 247.8059, 247.2785, 248.8009, 
    248.0471, 249.5266, 250.1565, 250.7543, 251.4472, 245.5584, 245.3555, 
    245.7198, 246.2218, 246.6896, 247.3099, 247.3739, 247.4898, 247.8003, 
    248.0533, 247.5254, 248.1169, 245.9228, 247.069, 245.2778, 245.8163, 
    246.1927, 246.0288, 246.8831, 247.084, 247.9091, 247.4788, 250.0001, 
    248.8883, 251.9784, 251.114, 245.2843, 245.5582, 246.5092, 246.0574, 
    247.3519, 247.679, 247.9385, 248.2686, 248.305, 248.5008, 248.1799, 
    248.4885, 247.3112, 247.8424, 246.402, 246.7497, 246.5901, 246.4142, 
    246.9569, 247.5333, 247.5473, 247.7409, 248.2581, 247.3571, 250.1405, 
    248.424, 245.8568, 246.3816, 246.4585, 246.2551, 247.647, 247.1368, 
    248.4962, 248.1316, 248.7295, 248.4322, 248.3884, 248.007, 247.7691, 
    247.1594, 246.6712, 246.2848, 246.3748, 246.7992, 247.569, 248.3076, 
    248.1475, 248.6841, 247.258, 247.8603, 247.6304, 248.2301, 246.9089, 
    248.0302, 246.6241, 246.7469, 247.1268, 247.8994, 248.0708, 248.2509, 
    248.1401, 247.5979, 247.5008, 247.118, 247.0115, 246.7203, 246.4784, 
    246.699, 246.9303, 247.5988, 248.1923, 248.8401, 248.9993, 249.7521, 
    249.137, 250.1497, 249.2852, 250.7836, 248.0971, 249.2632, 247.1447, 
    247.3723, 247.7912, 248.7352, 248.2273, 248.8221, 247.4975, 246.813, 
    246.638, 246.308, 246.6456, 246.6182, 246.941, 246.8374, 247.6207, 
    247.1959, 248.3869, 248.8178, 250.0372, 250.7838, 251.5465, 251.8824, 
    251.9848, 252.0275 ;

 FSH_G =
  257.0626, 257.7545, 257.6204, 258.1776, 257.8691, 258.2336, 257.2036, 
    257.7813, 257.4129, 257.1259, 259.2565, 258.2027, 260.3561, 259.6845, 
    261.3829, 260.2506, 261.6097, 261.3522, 262.1315, 261.9084, 262.9018, 
    262.2346, 263.4196, 262.7433, 262.8485, 262.2122, 258.4164, 259.1248, 
    258.3741, 258.4752, 258.4302, 257.8749, 257.594, 257.0109, 257.117, 
    257.546, 258.5207, 258.191, 259.0251, 259.0063, 259.9326, 259.5154, 
    261.0809, 260.6299, 261.9177, 261.5958, 261.9023, 261.8096, 261.9035, 
    261.4315, 261.6336, 261.2188, 259.5932, 260.0678, 258.6496, 257.7932, 
    257.2286, 256.8268, 256.8836, 256.9915, 257.5484, 258.0736, 258.4732, 
    258.7402, 259.0036, 259.7955, 260.2177, 261.1695, 261.0007, 261.2877, 
    261.5638, 262.0256, 261.9498, 262.153, 261.2811, 261.86, 260.9043, 
    261.1655, 259.0695, 258.2802, 257.9397, 257.6459, 256.9271, 257.4232, 
    257.2275, 257.6943, 257.9901, 257.8441, 258.7476, 258.3962, 260.2428, 
    259.4484, 261.5316, 261.0355, 261.6508, 261.3371, 261.8741, 261.3908, 
    262.229, 262.4109, 262.2865, 262.7664, 261.3638, 261.9017, 257.8397, 
    257.8635, 257.975, 257.4848, 257.4551, 257.0077, 257.4063, 257.5756, 
    258.0078, 258.2623, 258.5045, 259.0373, 259.6308, 260.4612, 261.0676, 
    261.4678, 261.2227, 261.4391, 261.1971, 261.0839, 262.3424, 261.6352, 
    262.6973, 262.6387, 262.1576, 262.6454, 257.8803, 257.7432, 257.2655, 
    257.6394, 256.959, 257.3391, 257.5572, 258.4023, 258.5892, 258.7608, 
    259.101, 259.5367, 260.2993, 260.9727, 261.5801, 261.5357, 261.5513, 
    261.6865, 261.351, 261.7416, 261.8066, 261.6357, 262.6309, 262.3466, 
    262.6375, 262.4525, 257.7879, 258.0189, 257.894, 258.1285, 257.9628, 
    258.6977, 258.9179, 259.9492, 259.5278, 260.1999, 259.5966, 259.7032, 
    260.2194, 259.6295, 260.935, 260.0449, 261.6917, 260.8004, 261.7469, 
    261.5775, 261.8585, 262.1095, 262.4264, 263.0095, 262.8747, 263.3633, 
    258.3636, 258.6625, 258.6373, 258.9508, 259.1825, 259.6854, 260.4897, 
    260.1875, 260.7433, 260.8635, 260.0108, 260.5278, 258.8633, 259.1316, 
    258.9727, 258.3866, 260.2557, 259.2967, 261.0772, 260.5492, 262.0736, 
    261.3188, 262.8003, 263.431, 264.0296, 264.7234, 258.8268, 258.6236, 
    258.9884, 259.491, 259.9595, 260.5806, 260.6447, 260.7607, 261.0717, 
    261.325, 260.7964, 261.3886, 259.1916, 260.3394, 258.5458, 259.0851, 
    259.4619, 259.2978, 260.1533, 260.3545, 261.1806, 260.7498, 263.2744, 
    262.161, 265.2553, 264.3897, 258.5523, 258.8266, 259.7789, 259.3264, 
    260.6226, 260.9502, 261.2101, 261.5406, 261.5771, 261.773, 261.4518, 
    261.7608, 260.5819, 261.1138, 259.6715, 260.0197, 259.8599, 259.6838, 
    260.2272, 260.8043, 260.8184, 261.0122, 261.5299, 260.6279, 263.4149, 
    261.6961, 259.1256, 259.6511, 259.7281, 259.5244, 260.9182, 260.4073, 
    261.7685, 261.4034, 262.0021, 261.7044, 261.6606, 261.2786, 261.0404, 
    260.4299, 259.941, 259.5542, 259.6443, 260.0692, 260.84, 261.5796, 
    261.4193, 261.9566, 260.5286, 261.1317, 260.9015, 261.502, 260.1791, 
    261.3018, 259.8939, 260.0169, 260.3973, 261.1708, 261.3425, 261.5228, 
    261.4119, 260.8689, 260.7717, 260.3885, 260.2818, 259.9902, 259.748, 
    259.9689, 260.2005, 260.8699, 261.4642, 262.1129, 262.2722, 263.026, 
    262.4101, 263.4242, 262.5584, 264.0589, 261.3688, 262.5364, 260.4152, 
    260.6431, 261.0625, 262.0078, 261.4992, 262.0948, 260.7684, 260.083, 
    259.9078, 259.5774, 259.9154, 259.888, 260.2113, 260.1075, 260.8918, 
    260.4664, 261.659, 262.0905, 263.3115, 264.0591, 264.8229, 265.1592, 
    265.2617, 265.3045 ;

 FSH_NODYNLNDUSE =
  243.7966, 244.4876, 244.3536, 244.9102, 244.6021, 244.966, 243.9374, 
    244.5144, 244.1465, 243.8598, 245.9876, 244.9352, 247.0857, 246.4149, 
    248.1112, 246.9804, 248.3377, 248.0805, 248.8588, 248.6359, 249.6281, 
    248.9617, 250.1451, 249.4698, 249.5748, 248.9394, 245.1486, 245.8561, 
    245.1063, 245.2073, 245.1624, 244.6078, 244.3273, 243.7449, 243.851, 
    244.2793, 245.2527, 244.9235, 245.7565, 245.7377, 246.6628, 246.2461, 
    247.8095, 247.3591, 248.6452, 248.3238, 248.6298, 248.5372, 248.6311, 
    248.1597, 248.3615, 247.9473, 246.3238, 246.7978, 245.3815, 244.5263, 
    243.9624, 243.5611, 243.6178, 243.7256, 244.2818, 244.8062, 245.2054, 
    245.472, 245.735, 246.5259, 246.9475, 247.898, 247.7295, 248.0161, 
    248.2919, 248.753, 248.6773, 248.8802, 248.0095, 248.5876, 247.6331, 
    247.894, 245.8008, 245.0126, 244.6725, 244.3792, 243.6613, 244.1567, 
    243.9613, 244.4275, 244.7229, 244.577, 245.4793, 245.1284, 246.9725, 
    246.1792, 248.2597, 247.7642, 248.3787, 248.0654, 248.6017, 248.119, 
    248.9561, 249.1378, 249.0135, 249.4928, 248.0921, 248.6293, 244.5727, 
    244.5964, 244.7078, 244.2182, 244.1886, 243.7417, 244.1399, 244.309, 
    244.7405, 244.9947, 245.2366, 245.7686, 246.3614, 247.1906, 247.7962, 
    248.196, 247.9512, 248.1673, 247.9255, 247.8125, 249.0694, 248.3631, 
    249.4238, 249.3653, 248.8848, 249.3719, 244.6132, 244.4763, 243.9992, 
    244.3726, 243.6932, 244.0727, 244.2906, 245.1345, 245.3212, 245.4925, 
    245.8323, 246.2674, 247.029, 247.7015, 248.3081, 248.2638, 248.2793, 
    248.4143, 248.0793, 248.4694, 248.5343, 248.3637, 249.3574, 249.0736, 
    249.3641, 249.1794, 244.521, 244.7516, 244.6269, 244.8611, 244.6956, 
    245.4295, 245.6494, 246.6793, 246.2585, 246.9297, 246.3271, 246.4336, 
    246.9492, 246.3601, 247.6639, 246.7749, 248.4196, 247.5294, 248.4746, 
    248.3055, 248.5861, 248.8368, 249.1533, 249.7356, 249.601, 250.0889, 
    245.0959, 245.3944, 245.3691, 245.6823, 245.9136, 246.4158, 247.2191, 
    246.9173, 247.4724, 247.5925, 246.7408, 247.2572, 245.5949, 245.8628, 
    245.7041, 245.1188, 246.9854, 246.0277, 247.8059, 247.2785, 248.8009, 
    248.0471, 249.5266, 250.1565, 250.7543, 251.4472, 245.5584, 245.3555, 
    245.7198, 246.2218, 246.6896, 247.3099, 247.3739, 247.4898, 247.8003, 
    248.0533, 247.5254, 248.1169, 245.9228, 247.069, 245.2778, 245.8163, 
    246.1927, 246.0288, 246.8831, 247.084, 247.9091, 247.4788, 250.0001, 
    248.8883, 251.9784, 251.114, 245.2843, 245.5582, 246.5092, 246.0574, 
    247.3519, 247.679, 247.9385, 248.2686, 248.305, 248.5008, 248.1799, 
    248.4885, 247.3112, 247.8424, 246.402, 246.7497, 246.5901, 246.4142, 
    246.9569, 247.5333, 247.5473, 247.7409, 248.2581, 247.3571, 250.1405, 
    248.424, 245.8568, 246.3816, 246.4585, 246.2551, 247.647, 247.1368, 
    248.4962, 248.1316, 248.7295, 248.4322, 248.3884, 248.007, 247.7691, 
    247.1594, 246.6712, 246.2848, 246.3748, 246.7992, 247.569, 248.3076, 
    248.1475, 248.6841, 247.258, 247.8603, 247.6304, 248.2301, 246.9089, 
    248.0302, 246.6241, 246.7469, 247.1268, 247.8994, 248.0708, 248.2509, 
    248.1401, 247.5979, 247.5008, 247.118, 247.0115, 246.7203, 246.4784, 
    246.699, 246.9303, 247.5988, 248.1923, 248.8401, 248.9993, 249.7521, 
    249.137, 250.1497, 249.2852, 250.7836, 248.0971, 249.2632, 247.1447, 
    247.3723, 247.7912, 248.7352, 248.2273, 248.8221, 247.4975, 246.813, 
    246.638, 246.308, 246.6456, 246.6182, 246.941, 246.8374, 247.6207, 
    247.1959, 248.3869, 248.8178, 250.0372, 250.7838, 251.5465, 251.8824, 
    251.9848, 252.0275 ;

 FSH_R =
  243.7966, 244.4876, 244.3536, 244.9102, 244.6021, 244.966, 243.9374, 
    244.5144, 244.1465, 243.8598, 245.9876, 244.9352, 247.0857, 246.4149, 
    248.1112, 246.9804, 248.3377, 248.0805, 248.8588, 248.6359, 249.6281, 
    248.9617, 250.1451, 249.4698, 249.5748, 248.9394, 245.1486, 245.8561, 
    245.1063, 245.2073, 245.1624, 244.6078, 244.3273, 243.7449, 243.851, 
    244.2793, 245.2527, 244.9235, 245.7565, 245.7377, 246.6628, 246.2461, 
    247.8095, 247.3591, 248.6452, 248.3238, 248.6298, 248.5372, 248.6311, 
    248.1597, 248.3615, 247.9473, 246.3238, 246.7978, 245.3815, 244.5263, 
    243.9624, 243.5611, 243.6178, 243.7256, 244.2818, 244.8062, 245.2054, 
    245.472, 245.735, 246.5259, 246.9475, 247.898, 247.7295, 248.0161, 
    248.2919, 248.753, 248.6773, 248.8802, 248.0095, 248.5876, 247.6331, 
    247.894, 245.8008, 245.0126, 244.6725, 244.3792, 243.6613, 244.1567, 
    243.9613, 244.4275, 244.7229, 244.577, 245.4793, 245.1284, 246.9725, 
    246.1792, 248.2597, 247.7642, 248.3787, 248.0654, 248.6017, 248.119, 
    248.9561, 249.1378, 249.0135, 249.4928, 248.0921, 248.6293, 244.5727, 
    244.5964, 244.7078, 244.2182, 244.1886, 243.7417, 244.1399, 244.309, 
    244.7405, 244.9947, 245.2366, 245.7686, 246.3614, 247.1906, 247.7962, 
    248.196, 247.9512, 248.1673, 247.9255, 247.8125, 249.0694, 248.3631, 
    249.4238, 249.3653, 248.8848, 249.3719, 244.6132, 244.4763, 243.9992, 
    244.3726, 243.6932, 244.0727, 244.2906, 245.1345, 245.3212, 245.4925, 
    245.8323, 246.2674, 247.029, 247.7015, 248.3081, 248.2638, 248.2793, 
    248.4143, 248.0793, 248.4694, 248.5343, 248.3637, 249.3574, 249.0736, 
    249.3641, 249.1794, 244.521, 244.7516, 244.6269, 244.8611, 244.6956, 
    245.4295, 245.6494, 246.6793, 246.2585, 246.9297, 246.3271, 246.4336, 
    246.9492, 246.3601, 247.6639, 246.7749, 248.4196, 247.5294, 248.4746, 
    248.3055, 248.5861, 248.8368, 249.1533, 249.7356, 249.601, 250.0889, 
    245.0959, 245.3944, 245.3691, 245.6823, 245.9136, 246.4158, 247.2191, 
    246.9173, 247.4724, 247.5925, 246.7408, 247.2572, 245.5949, 245.8628, 
    245.7041, 245.1188, 246.9854, 246.0277, 247.8059, 247.2785, 248.8009, 
    248.0471, 249.5266, 250.1565, 250.7543, 251.4472, 245.5584, 245.3555, 
    245.7198, 246.2218, 246.6896, 247.3099, 247.3739, 247.4898, 247.8003, 
    248.0533, 247.5254, 248.1169, 245.9228, 247.069, 245.2778, 245.8163, 
    246.1927, 246.0288, 246.8831, 247.084, 247.9091, 247.4788, 250.0001, 
    248.8883, 251.9784, 251.114, 245.2843, 245.5582, 246.5092, 246.0574, 
    247.3519, 247.679, 247.9385, 248.2686, 248.305, 248.5008, 248.1799, 
    248.4885, 247.3112, 247.8424, 246.402, 246.7497, 246.5901, 246.4142, 
    246.9569, 247.5333, 247.5473, 247.7409, 248.2581, 247.3571, 250.1405, 
    248.424, 245.8568, 246.3816, 246.4585, 246.2551, 247.647, 247.1368, 
    248.4962, 248.1316, 248.7295, 248.4322, 248.3884, 248.007, 247.7691, 
    247.1594, 246.6712, 246.2848, 246.3748, 246.7992, 247.569, 248.3076, 
    248.1475, 248.6841, 247.258, 247.8603, 247.6304, 248.2301, 246.9089, 
    248.0302, 246.6241, 246.7469, 247.1268, 247.8994, 248.0708, 248.2509, 
    248.1401, 247.5979, 247.5008, 247.118, 247.0115, 246.7203, 246.4784, 
    246.699, 246.9303, 247.5988, 248.1923, 248.8401, 248.9993, 249.7521, 
    249.137, 250.1497, 249.2852, 250.7836, 248.0971, 249.2632, 247.1447, 
    247.3723, 247.7912, 248.7352, 248.2273, 248.8221, 247.4975, 246.813, 
    246.638, 246.308, 246.6456, 246.6182, 246.941, 246.8374, 247.6207, 
    247.1959, 248.3869, 248.8178, 250.0372, 250.7838, 251.5465, 251.8824, 
    251.9848, 252.0275 ;

 FSH_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSH_V =
  -13.26599, -13.26692, -13.26674, -13.26748, -13.26708, -13.26756, 
    -13.26618, -13.26695, -13.26647, -13.26608, -13.26891, -13.26752, 
    -13.27039, -13.26952, -13.27173, -13.27024, -13.27204, -13.27171, 
    -13.27275, -13.27245, -13.27375, -13.27289, -13.27446, -13.27355, 
    -13.27369, -13.27285, -13.26782, -13.26873, -13.26776, -13.26789, 
    -13.26783, -13.26708, -13.26669, -13.26593, -13.26607, -13.26664, 
    -13.26795, -13.26751, -13.26864, -13.26862, -13.26985, -13.2693, 
    -13.27135, -13.27077, -13.27246, -13.27203, -13.27244, -13.27232, 
    -13.27244, -13.27181, -13.27208, -13.27153, -13.2694, -13.27002, 
    -13.26813, -13.26695, -13.26621, -13.26568, -13.26576, -13.2659, 
    -13.26664, -13.26736, -13.2679, -13.26826, -13.26861, -13.26964, 
    -13.27021, -13.27145, -13.27124, -13.27161, -13.27199, -13.2726, 
    -13.2725, -13.27277, -13.27162, -13.27238, -13.27112, -13.27146, 
    -13.26865, -13.26763, -13.26715, -13.26677, -13.26581, -13.26647, 
    -13.26621, -13.26685, -13.26724, -13.26705, -13.26827, -13.26779, 
    -13.27024, -13.2692, -13.27195, -13.27129, -13.27211, -13.27169, 
    -13.2724, -13.27176, -13.27287, -13.27311, -13.27295, -13.27359, 
    -13.27172, -13.27243, -13.26704, -13.26707, -13.26723, -13.26655, 
    -13.26652, -13.26592, -13.26646, -13.26668, -13.26727, -13.26761, 
    -13.26793, -13.26865, -13.26944, -13.27054, -13.27133, -13.27186, 
    -13.27154, -13.27183, -13.2715, -13.27136, -13.27302, -13.27208, 
    -13.2735, -13.27342, -13.27277, -13.27343, -13.2671, -13.26691, 
    -13.26627, -13.26677, -13.26586, -13.26636, -13.26665, -13.26779, 
    -13.26805, -13.26828, -13.26874, -13.26933, -13.27033, -13.2712, 
    -13.27201, -13.27196, -13.27198, -13.27215, -13.27171, -13.27223, 
    -13.27231, -13.27209, -13.27341, -13.27303, -13.27342, -13.27318, 
    -13.26697, -13.26728, -13.26711, -13.26743, -13.2672, -13.26818, 
    -13.26848, -13.26985, -13.26931, -13.27019, -13.26941, -13.26954, 
    -13.2702, -13.26945, -13.27114, -13.26997, -13.27216, -13.27097, 
    -13.27223, -13.27201, -13.27238, -13.27271, -13.27314, -13.27391, 
    -13.27373, -13.27439, -13.26775, -13.26814, -13.26812, -13.26854, 
    -13.26885, -13.26953, -13.27058, -13.27019, -13.27093, -13.27106, 
    -13.26996, -13.27063, -13.26841, -13.26877, -13.26857, -13.26777, 
    -13.27026, -13.26899, -13.27134, -13.27066, -13.27267, -13.27165, 
    -13.27363, -13.27446, -13.27529, -13.27621, -13.26837, -13.2681, 
    -13.26859, -13.26925, -13.26988, -13.2707, -13.27079, -13.27094, 
    -13.27134, -13.27167, -13.27098, -13.27176, -13.26882, -13.27038, 
    -13.26799, -13.2687, -13.26922, -13.26901, -13.27015, -13.27041, 
    -13.27147, -13.27093, -13.27424, -13.27277, -13.27695, -13.27576, 
    -13.268, -13.26837, -13.26964, -13.26905, -13.27077, -13.27117, 
    -13.27152, -13.27195, -13.27201, -13.27226, -13.27184, -13.27225, 
    -13.27071, -13.27139, -13.26951, -13.26996, -13.26976, -13.26953, 
    -13.27024, -13.27099, -13.27102, -13.27125, -13.27188, -13.27077, 
    -13.2744, -13.27211, -13.26878, -13.26946, -13.26958, -13.26931, 
    -13.27113, -13.27048, -13.27226, -13.27178, -13.27257, -13.27218, 
    -13.27212, -13.27161, -13.27129, -13.2705, -13.26986, -13.26936, 
    -13.26947, -13.27003, -13.27104, -13.27201, -13.27179, -13.27251, 
    -13.27064, -13.27141, -13.2711, -13.27191, -13.27017, -13.27159, 
    -13.2698, -13.26997, -13.27046, -13.27145, -13.2717, -13.27193, 
    -13.27179, -13.27106, -13.27096, -13.27046, -13.27031, -13.26993, 
    -13.26961, -13.2699, -13.2702, -13.27107, -13.27185, -13.27272, 
    -13.27293, -13.2739, -13.27309, -13.27441, -13.27325, -13.27529, 
    -13.2717, -13.27325, -13.27049, -13.27079, -13.27131, -13.27256, 
    -13.2719, -13.27268, -13.27095, -13.27003, -13.26982, -13.26938, 
    -13.26983, -13.2698, -13.27022, -13.27009, -13.2711, -13.27056, 
    -13.27211, -13.27268, -13.27431, -13.27531, -13.27637, -13.27683, 
    -13.27697, -13.27702 ;

 FSM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSNO_EFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSR =
  1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 1.081658, 
    1.081658, 1.081658 ;

 FSRND =
  0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 0.1614004, 
    0.1614004, 0.1614004 ;

 FSRNDLN =
  0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 0.2604372, 
    0.2604372, 0.2604372 ;

 FSRNI =
  0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 0.3794284, 
    0.3794284, 0.3794284 ;

 FSRVD =
  0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 0.09660081, 
    0.09660081, 0.09660081 ;

 FSRVDLN =
  0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 0.1560678, 
    0.1560678, 0.1560678 ;

 FSRVI =
  0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 0.444228, 
    0.444228, 0.444228 ;

 FUELC =
  0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806 ;

 F_DENIT =
  1.095188e-14, 1.099342e-14, 1.09853e-14, 1.101883e-14, 1.10002e-14, 
    1.102213e-14, 1.09602e-14, 1.099496e-14, 1.097274e-14, 1.095546e-14, 
    1.108377e-14, 1.102018e-14, 1.114976e-14, 1.110917e-14, 1.121104e-14, 
    1.114341e-14, 1.122466e-14, 1.120902e-14, 1.125594e-14, 1.124247e-14, 
    1.130251e-14, 1.12621e-14, 1.133359e-14, 1.129282e-14, 1.129918e-14, 
    1.126068e-14, 1.103308e-14, 1.107599e-14, 1.103051e-14, 1.103663e-14, 
    1.103386e-14, 1.100052e-14, 1.098373e-14, 1.094853e-14, 1.095489e-14, 
    1.098072e-14, 1.103925e-14, 1.101933e-14, 1.10694e-14, 1.106828e-14, 
    1.112404e-14, 1.109888e-14, 1.119266e-14, 1.116596e-14, 1.124301e-14, 
    1.12236e-14, 1.124207e-14, 1.123643e-14, 1.124209e-14, 1.121367e-14, 
    1.12258e-14, 1.12008e-14, 1.110381e-14, 1.11324e-14, 1.104706e-14, 
    1.099576e-14, 1.096165e-14, 1.093749e-14, 1.094087e-14, 1.094739e-14, 
    1.098084e-14, 1.101227e-14, 1.103625e-14, 1.105227e-14, 1.106806e-14, 
    1.111598e-14, 1.114129e-14, 1.119802e-14, 1.118775e-14, 1.120509e-14, 
    1.122165e-14, 1.124947e-14, 1.124487e-14, 1.125712e-14, 1.120452e-14, 
    1.123947e-14, 1.118175e-14, 1.119753e-14, 1.10726e-14, 1.102478e-14, 
    1.10045e-14, 1.09867e-14, 1.094348e-14, 1.097332e-14, 1.096153e-14, 
    1.098947e-14, 1.100724e-14, 1.099842e-14, 1.105269e-14, 1.103156e-14, 
    1.114276e-14, 1.109485e-14, 1.121974e-14, 1.118981e-14, 1.122686e-14, 
    1.120794e-14, 1.124032e-14, 1.121115e-14, 1.126164e-14, 1.127266e-14, 
    1.12651e-14, 1.129398e-14, 1.120942e-14, 1.124189e-14, 1.099828e-14, 
    1.099972e-14, 1.100638e-14, 1.097699e-14, 1.097519e-14, 1.094825e-14, 
    1.097216e-14, 1.098237e-14, 1.100822e-14, 1.102351e-14, 1.103805e-14, 
    1.107007e-14, 1.110582e-14, 1.115581e-14, 1.119173e-14, 1.121579e-14, 
    1.120101e-14, 1.121403e-14, 1.119944e-14, 1.119257e-14, 1.126848e-14, 
    1.122585e-14, 1.128978e-14, 1.128624e-14, 1.125727e-14, 1.128658e-14, 
    1.100069e-14, 1.099241e-14, 1.096376e-14, 1.098615e-14, 1.094528e-14, 
    1.096815e-14, 1.098128e-14, 1.103199e-14, 1.10431e-14, 1.105345e-14, 
    1.107384e-14, 1.110003e-14, 1.114602e-14, 1.118601e-14, 1.122254e-14, 
    1.121983e-14, 1.122077e-14, 1.122891e-14, 1.120868e-14, 1.123219e-14, 
    1.123612e-14, 1.122579e-14, 1.128571e-14, 1.126858e-14, 1.128609e-14, 
    1.12749e-14, 1.099507e-14, 1.100893e-14, 1.10014e-14, 1.101552e-14, 
    1.100554e-14, 1.104976e-14, 1.1063e-14, 1.112502e-14, 1.109951e-14, 
    1.114006e-14, 1.110359e-14, 1.111005e-14, 1.114134e-14, 1.110551e-14, 
    1.118376e-14, 1.113069e-14, 1.12292e-14, 1.117622e-14, 1.123249e-14, 
    1.122223e-14, 1.123914e-14, 1.125431e-14, 1.127334e-14, 1.130856e-14, 
    1.130037e-14, 1.132981e-14, 1.102961e-14, 1.104761e-14, 1.1046e-14, 
    1.106483e-14, 1.107876e-14, 1.110899e-14, 1.115746e-14, 1.113919e-14, 
    1.117265e-14, 1.117938e-14, 1.112847e-14, 1.115971e-14, 1.105948e-14, 
    1.107565e-14, 1.106599e-14, 1.103076e-14, 1.114326e-14, 1.108549e-14, 
    1.119211e-14, 1.116079e-14, 1.125209e-14, 1.120668e-14, 1.129586e-14, 
    1.133405e-14, 1.136991e-14, 1.141187e-14, 1.105741e-14, 1.104514e-14, 
    1.106704e-14, 1.109739e-14, 1.112549e-14, 1.116292e-14, 1.116672e-14, 
    1.11737e-14, 1.119184e-14, 1.120712e-14, 1.117589e-14, 1.12109e-14, 
    1.10794e-14, 1.114826e-14, 1.104028e-14, 1.10728e-14, 1.109534e-14, 
    1.108543e-14, 1.113687e-14, 1.114897e-14, 1.119827e-14, 1.117277e-14, 
    1.132458e-14, 1.125739e-14, 1.144378e-14, 1.139168e-14, 1.104084e-14, 
    1.105729e-14, 1.111464e-14, 1.108734e-14, 1.116536e-14, 1.118458e-14, 
    1.120016e-14, 1.122015e-14, 1.122226e-14, 1.123411e-14, 1.121466e-14, 
    1.12333e-14, 1.11628e-14, 1.119429e-14, 1.110786e-14, 1.112887e-14, 
    1.111918e-14, 1.110854e-14, 1.114126e-14, 1.117618e-14, 1.117688e-14, 
    1.118805e-14, 1.121963e-14, 1.116533e-14, 1.133321e-14, 1.122952e-14, 
    1.107524e-14, 1.110698e-14, 1.111147e-14, 1.109917e-14, 1.11826e-14, 
    1.115236e-14, 1.123381e-14, 1.121176e-14, 1.124782e-14, 1.122989e-14, 
    1.122722e-14, 1.120419e-14, 1.118981e-14, 1.115361e-14, 1.11241e-14, 
    1.110074e-14, 1.110613e-14, 1.11318e-14, 1.117825e-14, 1.122224e-14, 
    1.121258e-14, 1.124485e-14, 1.115932e-14, 1.119518e-14, 1.118129e-14, 
    1.121741e-14, 1.113864e-14, 1.12061e-14, 1.112138e-14, 1.112877e-14, 
    1.115171e-14, 1.119791e-14, 1.120806e-14, 1.121898e-14, 1.12122e-14, 
    1.117957e-14, 1.117419e-14, 1.115102e-14, 1.114462e-14, 1.112699e-14, 
    1.111236e-14, 1.11257e-14, 1.113967e-14, 1.117943e-14, 1.121525e-14, 
    1.12543e-14, 1.126385e-14, 1.130953e-14, 1.127234e-14, 1.13337e-14, 
    1.128153e-14, 1.137178e-14, 1.120993e-14, 1.128034e-14, 1.115275e-14, 
    1.116646e-14, 1.119131e-14, 1.124829e-14, 1.121747e-14, 1.125348e-14, 
    1.117397e-14, 1.113273e-14, 1.112202e-14, 1.110213e-14, 1.112244e-14, 
    1.112079e-14, 1.114024e-14, 1.113395e-14, 1.11807e-14, 1.115558e-14, 
    1.122691e-14, 1.125297e-14, 1.132652e-14, 1.137161e-14, 1.141751e-14, 
    1.143776e-14, 1.144392e-14, 1.144648e-14 ;

 F_DENIT_vr =
  6.253638e-13, 6.277359e-13, 6.272722e-13, 6.291864e-13, 6.281229e-13, 
    6.293749e-13, 6.25839e-13, 6.278233e-13, 6.265548e-13, 6.255678e-13, 
    6.328945e-13, 6.292634e-13, 6.366629e-13, 6.343449e-13, 6.401619e-13, 
    6.363001e-13, 6.409394e-13, 6.400468e-13, 6.427261e-13, 6.419566e-13, 
    6.453852e-13, 6.430776e-13, 6.471599e-13, 6.448317e-13, 6.451949e-13, 
    6.429966e-13, 6.300004e-13, 6.324504e-13, 6.298535e-13, 6.302029e-13, 
    6.300447e-13, 6.281408e-13, 6.271824e-13, 6.251723e-13, 6.255354e-13, 
    6.270105e-13, 6.303524e-13, 6.292152e-13, 6.320744e-13, 6.3201e-13, 
    6.351939e-13, 6.337575e-13, 6.391122e-13, 6.375878e-13, 6.419874e-13, 
    6.408793e-13, 6.419336e-13, 6.41612e-13, 6.419347e-13, 6.40312e-13, 
    6.41005e-13, 6.39577e-13, 6.34039e-13, 6.356717e-13, 6.307983e-13, 
    6.278693e-13, 6.259218e-13, 6.24542e-13, 6.247349e-13, 6.251072e-13, 
    6.27017e-13, 6.288121e-13, 6.301812e-13, 6.310961e-13, 6.319977e-13, 
    6.34734e-13, 6.36179e-13, 6.394183e-13, 6.388321e-13, 6.398221e-13, 
    6.407679e-13, 6.423563e-13, 6.42094e-13, 6.427931e-13, 6.397898e-13, 
    6.417853e-13, 6.384894e-13, 6.393905e-13, 6.322568e-13, 6.295261e-13, 
    6.283686e-13, 6.27352e-13, 6.248842e-13, 6.265878e-13, 6.25915e-13, 
    6.275102e-13, 6.28525e-13, 6.280211e-13, 6.311199e-13, 6.299134e-13, 
    6.362631e-13, 6.335272e-13, 6.406589e-13, 6.389499e-13, 6.410651e-13, 
    6.399851e-13, 6.41834e-13, 6.401681e-13, 6.430515e-13, 6.436805e-13, 
    6.432486e-13, 6.448981e-13, 6.400693e-13, 6.419233e-13, 6.280133e-13, 
    6.280955e-13, 6.284755e-13, 6.267977e-13, 6.266946e-13, 6.251562e-13, 
    6.265219e-13, 6.271047e-13, 6.285808e-13, 6.29454e-13, 6.302839e-13, 
    6.321123e-13, 6.341536e-13, 6.37008e-13, 6.390594e-13, 6.404335e-13, 
    6.395892e-13, 6.403326e-13, 6.394995e-13, 6.391074e-13, 6.434421e-13, 
    6.410077e-13, 6.446578e-13, 6.444558e-13, 6.428017e-13, 6.444756e-13, 
    6.281509e-13, 6.276779e-13, 6.26042e-13, 6.273202e-13, 6.249868e-13, 
    6.262927e-13, 6.270425e-13, 6.299378e-13, 6.305723e-13, 6.311632e-13, 
    6.323277e-13, 6.33823e-13, 6.364492e-13, 6.387329e-13, 6.408186e-13, 
    6.40664e-13, 6.407175e-13, 6.411822e-13, 6.400269e-13, 6.413697e-13, 
    6.415943e-13, 6.410042e-13, 6.444257e-13, 6.434477e-13, 6.444473e-13, 
    6.438086e-13, 6.278299e-13, 6.286213e-13, 6.281915e-13, 6.289977e-13, 
    6.284278e-13, 6.30953e-13, 6.317088e-13, 6.3525e-13, 6.337937e-13, 
    6.361087e-13, 6.340265e-13, 6.343954e-13, 6.361821e-13, 6.341359e-13, 
    6.386042e-13, 6.355739e-13, 6.411991e-13, 6.381737e-13, 6.413866e-13, 
    6.408009e-13, 6.417663e-13, 6.426327e-13, 6.437196e-13, 6.457306e-13, 
    6.452625e-13, 6.46944e-13, 6.298023e-13, 6.308299e-13, 6.307382e-13, 
    6.318133e-13, 6.326085e-13, 6.343347e-13, 6.371027e-13, 6.360594e-13, 
    6.379698e-13, 6.383541e-13, 6.35447e-13, 6.372312e-13, 6.315075e-13, 
    6.324308e-13, 6.318793e-13, 6.298678e-13, 6.362915e-13, 6.329928e-13, 
    6.390808e-13, 6.372924e-13, 6.425062e-13, 6.399133e-13, 6.450055e-13, 
    6.471857e-13, 6.492333e-13, 6.516297e-13, 6.313898e-13, 6.306889e-13, 
    6.319392e-13, 6.336725e-13, 6.352767e-13, 6.374141e-13, 6.376311e-13, 
    6.380301e-13, 6.390657e-13, 6.399382e-13, 6.381548e-13, 6.401538e-13, 
    6.326454e-13, 6.365772e-13, 6.304114e-13, 6.322683e-13, 6.335553e-13, 
    6.329893e-13, 6.359266e-13, 6.366179e-13, 6.39433e-13, 6.379769e-13, 
    6.466451e-13, 6.428088e-13, 6.534515e-13, 6.504769e-13, 6.304436e-13, 
    6.313827e-13, 6.346572e-13, 6.330986e-13, 6.375534e-13, 6.386513e-13, 
    6.395409e-13, 6.406823e-13, 6.408027e-13, 6.414791e-13, 6.403689e-13, 
    6.41433e-13, 6.374073e-13, 6.392053e-13, 6.342705e-13, 6.354698e-13, 
    6.349167e-13, 6.343093e-13, 6.361776e-13, 6.381712e-13, 6.382114e-13, 
    6.388492e-13, 6.406525e-13, 6.375521e-13, 6.471382e-13, 6.412172e-13, 
    6.324076e-13, 6.342198e-13, 6.344764e-13, 6.337742e-13, 6.385383e-13, 
    6.368114e-13, 6.414624e-13, 6.40203e-13, 6.422622e-13, 6.412386e-13, 
    6.410857e-13, 6.397707e-13, 6.389499e-13, 6.368825e-13, 6.351977e-13, 
    6.338635e-13, 6.341714e-13, 6.356375e-13, 6.382899e-13, 6.408013e-13, 
    6.4025e-13, 6.420924e-13, 6.372088e-13, 6.392566e-13, 6.384631e-13, 
    6.40526e-13, 6.360276e-13, 6.3988e-13, 6.350424e-13, 6.354646e-13, 
    6.367741e-13, 6.39412e-13, 6.399918e-13, 6.406155e-13, 6.402283e-13, 
    6.383649e-13, 6.380578e-13, 6.36735e-13, 6.363694e-13, 6.353628e-13, 
    6.345274e-13, 6.35289e-13, 6.360865e-13, 6.38357e-13, 6.404023e-13, 
    6.426322e-13, 6.431775e-13, 6.457861e-13, 6.436622e-13, 6.471661e-13, 
    6.441872e-13, 6.493407e-13, 6.400988e-13, 6.441192e-13, 6.368336e-13, 
    6.376163e-13, 6.390356e-13, 6.422888e-13, 6.405291e-13, 6.425853e-13, 
    6.38045e-13, 6.356903e-13, 6.35079e-13, 6.339434e-13, 6.351029e-13, 
    6.350086e-13, 6.361192e-13, 6.357602e-13, 6.384293e-13, 6.36995e-13, 
    6.410682e-13, 6.425563e-13, 6.46756e-13, 6.493308e-13, 6.519517e-13, 
    6.53108e-13, 6.534599e-13, 6.53606e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 F_N2O_DENIT =
  3.320056e-16, 3.321001e-16, 3.320807e-16, 3.321552e-16, 3.321133e-16, 
    3.321609e-16, 3.32022e-16, 3.321002e-16, 3.320496e-16, 3.320091e-16, 
    3.322893e-16, 3.321541e-16, 3.324182e-16, 3.323378e-16, 3.325298e-16, 
    3.324049e-16, 3.325532e-16, 3.325244e-16, 3.326057e-16, 3.325819e-16, 
    3.326819e-16, 3.326148e-16, 3.327294e-16, 3.326649e-16, 3.326747e-16, 
    3.326099e-16, 3.321853e-16, 3.322771e-16, 3.321787e-16, 3.321922e-16, 
    3.321854e-16, 3.32112e-16, 3.320747e-16, 3.319927e-16, 3.320068e-16, 
    3.320663e-16, 3.321942e-16, 3.321501e-16, 3.322557e-16, 3.322535e-16, 
    3.323651e-16, 3.323151e-16, 3.324942e-16, 3.32444e-16, 3.325822e-16, 
    3.325478e-16, 3.325797e-16, 3.325691e-16, 3.325782e-16, 3.325287e-16, 
    3.32549e-16, 3.325045e-16, 3.323312e-16, 3.323869e-16, 3.322133e-16, 
    3.321018e-16, 3.320233e-16, 3.319671e-16, 3.319739e-16, 3.319894e-16, 
    3.320655e-16, 3.321343e-16, 3.321859e-16, 3.322192e-16, 3.322515e-16, 
    3.323499e-16, 3.323982e-16, 3.325031e-16, 3.324838e-16, 3.325148e-16, 
    3.325437e-16, 3.325913e-16, 3.325831e-16, 3.326033e-16, 3.325107e-16, 
    3.325727e-16, 3.324681e-16, 3.324973e-16, 3.322678e-16, 3.321642e-16, 
    3.321205e-16, 3.320795e-16, 3.319797e-16, 3.320487e-16, 3.320211e-16, 
    3.320834e-16, 3.321227e-16, 3.321023e-16, 3.322195e-16, 3.321738e-16, 
    3.324002e-16, 3.323056e-16, 3.325411e-16, 3.324865e-16, 3.32552e-16, 
    3.325186e-16, 3.325746e-16, 3.325233e-16, 3.326099e-16, 3.326286e-16, 
    3.326147e-16, 3.326623e-16, 3.325171e-16, 3.325744e-16, 3.321051e-16, 
    3.321084e-16, 3.321224e-16, 3.320563e-16, 3.320519e-16, 3.319891e-16, 
    3.320434e-16, 3.320668e-16, 3.321234e-16, 3.321561e-16, 3.321867e-16, 
    3.322543e-16, 3.323267e-16, 3.324231e-16, 3.324894e-16, 3.325318e-16, 
    3.325051e-16, 3.325276e-16, 3.325012e-16, 3.324879e-16, 3.326202e-16, 
    3.325472e-16, 3.32654e-16, 3.326483e-16, 3.325997e-16, 3.326474e-16, 
    3.321095e-16, 3.320902e-16, 3.320254e-16, 3.320752e-16, 3.319811e-16, 
    3.320342e-16, 3.320635e-16, 3.321744e-16, 3.321971e-16, 3.322192e-16, 
    3.322609e-16, 3.323136e-16, 3.324038e-16, 3.32478e-16, 3.325431e-16, 
    3.325375e-16, 3.32539e-16, 3.325526e-16, 3.325165e-16, 3.325573e-16, 
    3.325636e-16, 3.325455e-16, 3.32646e-16, 3.326177e-16, 3.32646e-16, 
    3.326267e-16, 3.320956e-16, 3.321255e-16, 3.321083e-16, 3.321396e-16, 
    3.321166e-16, 3.322125e-16, 3.322397e-16, 3.323643e-16, 3.323126e-16, 
    3.323927e-16, 3.323196e-16, 3.323328e-16, 3.323943e-16, 3.32322e-16, 
    3.324726e-16, 3.323715e-16, 3.325525e-16, 3.324573e-16, 3.325572e-16, 
    3.325384e-16, 3.325672e-16, 3.325935e-16, 3.326242e-16, 3.326819e-16, 
    3.326675e-16, 3.327141e-16, 3.3217e-16, 3.322079e-16, 3.322039e-16, 
    3.322428e-16, 3.32271e-16, 3.323321e-16, 3.324258e-16, 3.323899e-16, 
    3.324526e-16, 3.324653e-16, 3.323673e-16, 3.324278e-16, 3.322276e-16, 
    3.322607e-16, 3.3224e-16, 3.321648e-16, 3.323939e-16, 3.322788e-16, 
    3.32484e-16, 3.324251e-16, 3.325882e-16, 3.325093e-16, 3.326599e-16, 
    3.32721e-16, 3.327735e-16, 3.328335e-16, 3.322278e-16, 3.322009e-16, 
    3.322462e-16, 3.323091e-16, 3.323634e-16, 3.324353e-16, 3.324416e-16, 
    3.32454e-16, 3.324865e-16, 3.325143e-16, 3.324571e-16, 3.325196e-16, 
    3.322686e-16, 3.324032e-16, 3.321841e-16, 3.32253e-16, 3.322976e-16, 
    3.322774e-16, 3.323786e-16, 3.324012e-16, 3.324925e-16, 3.324454e-16, 
    3.32705e-16, 3.325954e-16, 3.328753e-16, 3.32804e-16, 3.321913e-16, 
    3.322252e-16, 3.323418e-16, 3.322869e-16, 3.324383e-16, 3.324742e-16, 
    3.325013e-16, 3.325374e-16, 3.325398e-16, 3.325608e-16, 3.325253e-16, 
    3.325582e-16, 3.324296e-16, 3.324878e-16, 3.323223e-16, 3.323632e-16, 
    3.323438e-16, 3.323219e-16, 3.323853e-16, 3.32452e-16, 3.324521e-16, 
    3.324722e-16, 3.325304e-16, 3.324287e-16, 3.327175e-16, 3.325458e-16, 
    3.32262e-16, 3.323262e-16, 3.32334e-16, 3.323093e-16, 3.324691e-16, 
    3.324126e-16, 3.325601e-16, 3.325204e-16, 3.325827e-16, 3.325519e-16, 
    3.325461e-16, 3.325053e-16, 3.324782e-16, 3.32411e-16, 3.323529e-16, 
    3.323064e-16, 3.323161e-16, 3.323671e-16, 3.324543e-16, 3.325336e-16, 
    3.325159e-16, 3.325712e-16, 3.324164e-16, 3.324832e-16, 3.324568e-16, 
    3.325219e-16, 3.323868e-16, 3.325141e-16, 3.323524e-16, 3.323661e-16, 
    3.324098e-16, 3.324963e-16, 3.325128e-16, 3.325326e-16, 3.325191e-16, 
    3.324604e-16, 3.324496e-16, 3.32405e-16, 3.323923e-16, 3.32358e-16, 
    3.323281e-16, 3.323546e-16, 3.323809e-16, 3.324559e-16, 3.325202e-16, 
    3.325872e-16, 3.326029e-16, 3.32678e-16, 3.32617e-16, 3.327158e-16, 
    3.326325e-16, 3.327714e-16, 3.325188e-16, 3.3264e-16, 3.324118e-16, 
    3.324368e-16, 3.324832e-16, 3.325832e-16, 3.325282e-16, 3.325914e-16, 
    3.324488e-16, 3.3237e-16, 3.323479e-16, 3.323086e-16, 3.323477e-16, 
    3.323445e-16, 3.323817e-16, 3.323687e-16, 3.324567e-16, 3.324097e-16, 
    3.325389e-16, 3.325843e-16, 3.327033e-16, 3.327709e-16, 3.328355e-16, 
    3.328622e-16, 3.328702e-16, 3.32873e-16 ;

 F_N2O_NIT =
  2.413928e-14, 2.434732e-14, 2.430679e-14, 2.447512e-14, 2.438167e-14, 
    2.449199e-14, 2.418137e-14, 2.435558e-14, 2.424429e-14, 2.415795e-14, 
    2.480347e-14, 2.448262e-14, 2.513901e-14, 2.493271e-14, 2.545261e-14, 
    2.510685e-14, 2.552262e-14, 2.544258e-14, 2.568383e-14, 2.561459e-14, 
    2.592445e-14, 2.571581e-14, 2.608582e-14, 2.587454e-14, 2.590753e-14, 
    2.570893e-14, 2.454703e-14, 2.476343e-14, 2.453423e-14, 2.456503e-14, 
    2.45512e-14, 2.438358e-14, 2.429935e-14, 2.412339e-14, 2.415528e-14, 
    2.428453e-14, 2.457886e-14, 2.447873e-14, 2.473145e-14, 2.472573e-14, 
    2.500862e-14, 2.488086e-14, 2.535883e-14, 2.52225e-14, 2.561748e-14, 
    2.551784e-14, 2.561279e-14, 2.558397e-14, 2.561315e-14, 2.546712e-14, 
    2.552963e-14, 2.540132e-14, 2.49048e-14, 2.505021e-14, 2.46178e-14, 
    2.435967e-14, 2.418899e-14, 2.406825e-14, 2.408529e-14, 2.411781e-14, 
    2.428529e-14, 2.444329e-14, 2.456405e-14, 2.4645e-14, 2.47249e-14, 
    2.496758e-14, 2.509651e-14, 2.538644e-14, 2.533398e-14, 2.542287e-14, 
    2.550794e-14, 2.565109e-14, 2.56275e-14, 2.569067e-14, 2.542051e-14, 
    2.559989e-14, 2.53041e-14, 2.538483e-14, 2.474669e-14, 2.450573e-14, 
    2.440371e-14, 2.431456e-14, 2.40984e-14, 2.424757e-14, 2.418871e-14, 
    2.432885e-14, 2.441812e-14, 2.437394e-14, 2.464721e-14, 2.454078e-14, 
    2.510416e-14, 2.486068e-14, 2.549801e-14, 2.534474e-14, 2.553481e-14, 
    2.543773e-14, 2.560419e-14, 2.545434e-14, 2.571419e-14, 2.577096e-14, 
    2.573216e-14, 2.588135e-14, 2.544603e-14, 2.561276e-14, 2.437272e-14, 
    2.437992e-14, 2.441348e-14, 2.426612e-14, 2.425712e-14, 2.41225e-14, 
    2.424226e-14, 2.429335e-14, 2.442329e-14, 2.450031e-14, 2.457365e-14, 
    2.473531e-14, 2.491649e-14, 2.517099e-14, 2.535465e-14, 2.547815e-14, 
    2.540238e-14, 2.546926e-14, 2.53945e-14, 2.535949e-14, 2.574968e-14, 
    2.55302e-14, 2.585986e-14, 2.584156e-14, 2.569215e-14, 2.584362e-14, 
    2.438497e-14, 2.434354e-14, 2.419998e-14, 2.431228e-14, 2.410786e-14, 
    2.422218e-14, 2.428803e-14, 2.4543e-14, 2.45992e-14, 2.465138e-14, 
    2.475459e-14, 2.488737e-14, 2.512121e-14, 2.532557e-14, 2.551288e-14, 
    2.549913e-14, 2.550396e-14, 2.55459e-14, 2.544209e-14, 2.556295e-14, 
    2.558327e-14, 2.553017e-14, 2.58391e-14, 2.575065e-14, 2.584116e-14, 
    2.578354e-14, 2.4357e-14, 2.442674e-14, 2.438904e-14, 2.445996e-14, 
    2.440998e-14, 2.463262e-14, 2.469957e-14, 2.50141e-14, 2.488476e-14, 
    2.509076e-14, 2.490564e-14, 2.493839e-14, 2.50975e-14, 2.491561e-14, 
    2.531428e-14, 2.504364e-14, 2.554753e-14, 2.527599e-14, 2.556458e-14, 
    2.551204e-14, 2.559905e-14, 2.567711e-14, 2.577548e-14, 2.595752e-14, 
    2.59153e-14, 2.606791e-14, 2.453092e-14, 2.462174e-14, 2.461373e-14, 
    2.470894e-14, 2.477948e-14, 2.493273e-14, 2.517954e-14, 2.508657e-14, 
    2.525736e-14, 2.529172e-14, 2.503229e-14, 2.519142e-14, 2.468259e-14, 
    2.476444e-14, 2.471568e-14, 2.453804e-14, 2.510796e-14, 2.481463e-14, 
    2.535766e-14, 2.519772e-14, 2.566597e-14, 2.543254e-14, 2.589207e-14, 
    2.608983e-14, 2.627664e-14, 2.649585e-14, 2.467137e-14, 2.460957e-14, 
    2.472027e-14, 2.487387e-14, 2.50168e-14, 2.520749e-14, 2.522704e-14, 
    2.526286e-14, 2.535576e-14, 2.543402e-14, 2.527419e-14, 2.545364e-14, 
    2.478344e-14, 2.51335e-14, 2.45862e-14, 2.475036e-14, 2.486476e-14, 
    2.481453e-14, 2.507592e-14, 2.513773e-14, 2.538973e-14, 2.52593e-14, 
    2.604095e-14, 2.56936e-14, 2.666337e-14, 2.639049e-14, 2.4588e-14, 
    2.467115e-14, 2.496169e-14, 2.482323e-14, 2.522024e-14, 2.531846e-14, 
    2.539845e-14, 2.55009e-14, 2.551197e-14, 2.557278e-14, 2.547316e-14, 
    2.556884e-14, 2.520787e-14, 2.536885e-14, 2.492835e-14, 2.50352e-14, 
    2.498601e-14, 2.493212e-14, 2.509863e-14, 2.527667e-14, 2.528047e-14, 
    2.53377e-14, 2.549935e-14, 2.52218e-14, 2.608596e-14, 2.555051e-14, 
    2.476198e-14, 2.492287e-14, 2.494589e-14, 2.488347e-14, 2.53086e-14, 
    2.515413e-14, 2.55713e-14, 2.54582e-14, 2.564364e-14, 2.55514e-14, 
    2.553784e-14, 2.541966e-14, 2.534622e-14, 2.516118e-14, 2.501114e-14, 
    2.489248e-14, 2.492004e-14, 2.505047e-14, 2.528757e-14, 2.551294e-14, 
    2.546348e-14, 2.562949e-14, 2.519129e-14, 2.537456e-14, 2.530364e-14, 
    2.548876e-14, 2.508409e-14, 2.542855e-14, 2.499644e-14, 2.503417e-14, 
    2.515106e-14, 2.538706e-14, 2.543941e-14, 2.549539e-14, 2.546083e-14, 
    2.529362e-14, 2.526628e-14, 2.51482e-14, 2.511564e-14, 2.502592e-14, 
    2.495176e-14, 2.501951e-14, 2.509076e-14, 2.529367e-14, 2.547726e-14, 
    2.567819e-14, 2.572749e-14, 2.596355e-14, 2.577131e-14, 2.608895e-14, 
    2.581878e-14, 2.628736e-14, 2.544856e-14, 2.581089e-14, 2.515639e-14, 
    2.522647e-14, 2.535351e-14, 2.564611e-14, 2.548792e-14, 2.567297e-14, 
    2.526521e-14, 2.505498e-14, 2.500073e-14, 2.489969e-14, 2.500304e-14, 
    2.499462e-14, 2.509371e-14, 2.506184e-14, 2.530041e-14, 2.517212e-14, 
    2.553746e-14, 2.567147e-14, 2.605186e-14, 2.628649e-14, 2.652643e-14, 
    2.663272e-14, 2.666511e-14, 2.667866e-14 ;

 F_NIT =
  4.023214e-11, 4.057886e-11, 4.051132e-11, 4.079187e-11, 4.063611e-11, 
    4.081998e-11, 4.030228e-11, 4.059263e-11, 4.040715e-11, 4.026324e-11, 
    4.133912e-11, 4.080437e-11, 4.189836e-11, 4.155451e-11, 4.242101e-11, 
    4.184475e-11, 4.25377e-11, 4.240431e-11, 4.280638e-11, 4.269099e-11, 
    4.320742e-11, 4.285968e-11, 4.347637e-11, 4.312423e-11, 4.317922e-11, 
    4.284821e-11, 4.091171e-11, 4.127238e-11, 4.089039e-11, 4.094171e-11, 
    4.091867e-11, 4.063931e-11, 4.049891e-11, 4.020565e-11, 4.02588e-11, 
    4.047422e-11, 4.096476e-11, 4.079789e-11, 4.121908e-11, 4.120955e-11, 
    4.168104e-11, 4.146811e-11, 4.226472e-11, 4.20375e-11, 4.269579e-11, 
    4.252973e-11, 4.268798e-11, 4.263995e-11, 4.268859e-11, 4.24452e-11, 
    4.254938e-11, 4.233553e-11, 4.1508e-11, 4.175035e-11, 4.102967e-11, 
    4.059946e-11, 4.031498e-11, 4.011375e-11, 4.014215e-11, 4.019636e-11, 
    4.047548e-11, 4.073881e-11, 4.094008e-11, 4.1075e-11, 4.120816e-11, 
    4.161264e-11, 4.182751e-11, 4.231073e-11, 4.22233e-11, 4.237145e-11, 
    4.251323e-11, 4.275182e-11, 4.27125e-11, 4.281778e-11, 4.236751e-11, 
    4.266649e-11, 4.21735e-11, 4.230805e-11, 4.124449e-11, 4.084289e-11, 
    4.067284e-11, 4.052426e-11, 4.016401e-11, 4.041261e-11, 4.031451e-11, 
    4.054808e-11, 4.069686e-11, 4.062323e-11, 4.107869e-11, 4.09013e-11, 
    4.184026e-11, 4.143447e-11, 4.249669e-11, 4.224123e-11, 4.255802e-11, 
    4.239621e-11, 4.267365e-11, 4.24239e-11, 4.285699e-11, 4.29516e-11, 
    4.288693e-11, 4.313559e-11, 4.241006e-11, 4.268794e-11, 4.062119e-11, 
    4.06332e-11, 4.068913e-11, 4.044353e-11, 4.042853e-11, 4.020417e-11, 
    4.040376e-11, 4.048891e-11, 4.070548e-11, 4.083386e-11, 4.095609e-11, 
    4.122551e-11, 4.152749e-11, 4.195166e-11, 4.225776e-11, 4.246358e-11, 
    4.23373e-11, 4.244877e-11, 4.232417e-11, 4.226582e-11, 4.291613e-11, 
    4.255034e-11, 4.309977e-11, 4.306927e-11, 4.282025e-11, 4.307269e-11, 
    4.064162e-11, 4.057256e-11, 4.03333e-11, 4.052047e-11, 4.017977e-11, 
    4.03703e-11, 4.048006e-11, 4.090501e-11, 4.099867e-11, 4.108563e-11, 
    4.125765e-11, 4.147896e-11, 4.186868e-11, 4.220928e-11, 4.252147e-11, 
    4.249854e-11, 4.250661e-11, 4.257649e-11, 4.240348e-11, 4.260492e-11, 
    4.263878e-11, 4.255028e-11, 4.306517e-11, 4.291774e-11, 4.30686e-11, 
    4.297257e-11, 4.059499e-11, 4.071124e-11, 4.064839e-11, 4.076661e-11, 
    4.06833e-11, 4.105436e-11, 4.116595e-11, 4.169017e-11, 4.14746e-11, 
    4.181794e-11, 4.15094e-11, 4.156398e-11, 4.182917e-11, 4.152603e-11, 
    4.219046e-11, 4.17394e-11, 4.257921e-11, 4.212665e-11, 4.260764e-11, 
    4.252007e-11, 4.266509e-11, 4.279519e-11, 4.295914e-11, 4.326253e-11, 
    4.319216e-11, 4.344651e-11, 4.088486e-11, 4.103623e-11, 4.102288e-11, 
    4.118157e-11, 4.129914e-11, 4.155455e-11, 4.196589e-11, 4.181095e-11, 
    4.20956e-11, 4.215286e-11, 4.172048e-11, 4.198569e-11, 4.113765e-11, 
    4.127406e-11, 4.11928e-11, 4.089673e-11, 4.18466e-11, 4.135771e-11, 
    4.226277e-11, 4.19962e-11, 4.277662e-11, 4.238757e-11, 4.315346e-11, 
    4.348306e-11, 4.37944e-11, 4.415975e-11, 4.111896e-11, 4.101595e-11, 
    4.120045e-11, 4.145645e-11, 4.169467e-11, 4.201249e-11, 4.204507e-11, 
    4.210476e-11, 4.22596e-11, 4.239003e-11, 4.212365e-11, 4.242274e-11, 
    4.130574e-11, 4.188917e-11, 4.0977e-11, 4.125059e-11, 4.144127e-11, 
    4.135756e-11, 4.17932e-11, 4.189622e-11, 4.231622e-11, 4.209883e-11, 
    4.340158e-11, 4.282267e-11, 4.443895e-11, 4.398416e-11, 4.098e-11, 
    4.111858e-11, 4.160281e-11, 4.137205e-11, 4.203373e-11, 4.219744e-11, 
    4.233075e-11, 4.25015e-11, 4.251995e-11, 4.262131e-11, 4.245526e-11, 
    4.261473e-11, 4.201312e-11, 4.228141e-11, 4.154726e-11, 4.172533e-11, 
    4.164335e-11, 4.155353e-11, 4.183105e-11, 4.212779e-11, 4.213412e-11, 
    4.22295e-11, 4.249891e-11, 4.203634e-11, 4.34766e-11, 4.258418e-11, 
    4.126998e-11, 4.153812e-11, 4.157647e-11, 4.147245e-11, 4.2181e-11, 
    4.192355e-11, 4.261883e-11, 4.243033e-11, 4.27394e-11, 4.258567e-11, 
    4.256306e-11, 4.23661e-11, 4.22437e-11, 4.19353e-11, 4.168523e-11, 
    4.148747e-11, 4.15334e-11, 4.175078e-11, 4.214596e-11, 4.252157e-11, 
    4.243914e-11, 4.271581e-11, 4.198548e-11, 4.229093e-11, 4.217273e-11, 
    4.248127e-11, 4.180683e-11, 4.238091e-11, 4.166073e-11, 4.172361e-11, 
    4.191843e-11, 4.231177e-11, 4.239901e-11, 4.249231e-11, 4.243472e-11, 
    4.215604e-11, 4.211047e-11, 4.191366e-11, 4.185941e-11, 4.170987e-11, 
    4.158628e-11, 4.169919e-11, 4.181793e-11, 4.215612e-11, 4.246209e-11, 
    4.279699e-11, 4.287915e-11, 4.327258e-11, 4.295218e-11, 4.348158e-11, 
    4.303129e-11, 4.381227e-11, 4.241427e-11, 4.301816e-11, 4.192731e-11, 
    4.204412e-11, 4.225585e-11, 4.274352e-11, 4.247986e-11, 4.278828e-11, 
    4.210868e-11, 4.175831e-11, 4.166788e-11, 4.149948e-11, 4.167173e-11, 
    4.16577e-11, 4.182285e-11, 4.176973e-11, 4.216736e-11, 4.195353e-11, 
    4.256244e-11, 4.278579e-11, 4.341977e-11, 4.381081e-11, 4.421071e-11, 
    4.438786e-11, 4.444185e-11, 4.446443e-11 ;

 F_NIT_vr =
  2.390771e-10, 2.401292e-10, 2.39924e-10, 2.407732e-10, 2.403018e-10, 
    2.408575e-10, 2.39289e-10, 2.401692e-10, 2.396069e-10, 2.391696e-10, 
    2.424208e-10, 2.408091e-10, 2.440969e-10, 2.43067e-10, 2.456546e-10, 
    2.43936e-10, 2.460011e-10, 2.456043e-10, 2.467978e-10, 2.464554e-10, 
    2.47983e-10, 2.469551e-10, 2.487753e-10, 2.47737e-10, 2.47899e-10, 
    2.469199e-10, 2.41135e-10, 2.422219e-10, 2.410702e-10, 2.412251e-10, 
    2.411553e-10, 2.403104e-10, 2.39885e-10, 2.389944e-10, 2.391556e-10, 
    2.398096e-10, 2.41293e-10, 2.407887e-10, 2.420587e-10, 2.4203e-10, 
    2.434453e-10, 2.428068e-10, 2.451885e-10, 2.445107e-10, 2.464693e-10, 
    2.45976e-10, 2.464457e-10, 2.463028e-10, 2.464468e-10, 2.45724e-10, 
    2.460331e-10, 2.453973e-10, 2.429293e-10, 2.436554e-10, 2.4149e-10, 
    2.401896e-10, 2.393266e-10, 2.387149e-10, 2.388008e-10, 2.389657e-10, 
    2.398129e-10, 2.406099e-10, 2.412179e-10, 2.416244e-10, 2.420252e-10, 
    2.432402e-10, 2.438833e-10, 2.45325e-10, 2.450645e-10, 2.455052e-10, 
    2.459267e-10, 2.466344e-10, 2.465178e-10, 2.468294e-10, 2.454922e-10, 
    2.463806e-10, 2.449139e-10, 2.453148e-10, 2.421368e-10, 2.409257e-10, 
    2.404114e-10, 2.399612e-10, 2.388671e-10, 2.396224e-10, 2.393243e-10, 
    2.400324e-10, 2.404827e-10, 2.402596e-10, 2.416352e-10, 2.410998e-10, 
    2.439211e-10, 2.427049e-10, 2.458778e-10, 2.451173e-10, 2.460594e-10, 
    2.455785e-10, 2.464021e-10, 2.456604e-10, 2.469451e-10, 2.472252e-10, 
    2.470332e-10, 2.477686e-10, 2.456177e-10, 2.464431e-10, 2.402548e-10, 
    2.402912e-10, 2.404602e-10, 2.397158e-10, 2.396702e-10, 2.389885e-10, 
    2.395943e-10, 2.398527e-10, 2.405082e-10, 2.408959e-10, 2.412647e-10, 
    2.420766e-10, 2.429837e-10, 2.442533e-10, 2.451663e-10, 2.457785e-10, 
    2.454027e-10, 2.457339e-10, 2.453631e-10, 2.45189e-10, 2.471195e-10, 
    2.46035e-10, 2.476621e-10, 2.47572e-10, 2.468349e-10, 2.475814e-10, 
    2.403162e-10, 2.401067e-10, 2.39381e-10, 2.399484e-10, 2.389138e-10, 
    2.394927e-10, 2.398253e-10, 2.411106e-10, 2.41393e-10, 2.416552e-10, 
    2.421728e-10, 2.428375e-10, 2.44005e-10, 2.450213e-10, 2.459502e-10, 
    2.458817e-10, 2.459056e-10, 2.461128e-10, 2.455985e-10, 2.461967e-10, 
    2.462969e-10, 2.460342e-10, 2.475592e-10, 2.471232e-10, 2.475691e-10, 
    2.472847e-10, 2.401744e-10, 2.405258e-10, 2.403354e-10, 2.40693e-10, 
    2.404405e-10, 2.415612e-10, 2.418971e-10, 2.434712e-10, 2.428244e-10, 
    2.438534e-10, 2.429284e-10, 2.430922e-10, 2.438861e-10, 2.429777e-10, 
    2.449644e-10, 2.436167e-10, 2.461206e-10, 2.447734e-10, 2.462045e-10, 
    2.459441e-10, 2.463743e-10, 2.467601e-10, 2.47245e-10, 2.481413e-10, 
    2.479331e-10, 2.48683e-10, 2.410503e-10, 2.415067e-10, 2.414663e-10, 
    2.419441e-10, 2.422975e-10, 2.430647e-10, 2.442957e-10, 2.438321e-10, 
    2.446823e-10, 2.44853e-10, 2.435606e-10, 2.443537e-10, 2.418098e-10, 
    2.4222e-10, 2.419755e-10, 2.410825e-10, 2.439368e-10, 2.424706e-10, 
    2.451783e-10, 2.44383e-10, 2.467044e-10, 2.455492e-10, 2.478187e-10, 
    2.487904e-10, 2.497052e-10, 2.50775e-10, 2.417558e-10, 2.414449e-10, 
    2.420005e-10, 2.427701e-10, 2.43484e-10, 2.444346e-10, 2.445315e-10, 
    2.447093e-10, 2.451704e-10, 2.455587e-10, 2.44765e-10, 2.456554e-10, 
    2.42315e-10, 2.44064e-10, 2.413242e-10, 2.421486e-10, 2.427212e-10, 
    2.424698e-10, 2.437759e-10, 2.440837e-10, 2.453361e-10, 2.446885e-10, 
    2.485498e-10, 2.468397e-10, 2.515899e-10, 2.502606e-10, 2.413362e-10, 
    2.417536e-10, 2.432086e-10, 2.42516e-10, 2.444973e-10, 2.449856e-10, 
    2.453821e-10, 2.4589e-10, 2.459443e-10, 2.462454e-10, 2.457516e-10, 
    2.462254e-10, 2.444338e-10, 2.452339e-10, 2.430393e-10, 2.435727e-10, 
    2.43327e-10, 2.430573e-10, 2.438883e-10, 2.447746e-10, 2.447932e-10, 
    2.450771e-10, 2.458785e-10, 2.445006e-10, 2.487697e-10, 2.46131e-10, 
    2.422091e-10, 2.430142e-10, 2.43129e-10, 2.428169e-10, 2.449359e-10, 
    2.441676e-10, 2.46238e-10, 2.456776e-10, 2.46595e-10, 2.461389e-10, 
    2.460713e-10, 2.454858e-10, 2.451208e-10, 2.442008e-10, 2.434521e-10, 
    2.428591e-10, 2.429965e-10, 2.43648e-10, 2.448281e-10, 2.459461e-10, 
    2.457008e-10, 2.46522e-10, 2.443483e-10, 2.452591e-10, 2.449064e-10, 
    2.458249e-10, 2.438188e-10, 2.455315e-10, 2.433811e-10, 2.435691e-10, 
    2.441516e-10, 2.453248e-10, 2.45584e-10, 2.458614e-10, 2.456897e-10, 
    2.448599e-10, 2.447238e-10, 2.441358e-10, 2.439732e-10, 2.435258e-10, 
    2.431549e-10, 2.434933e-10, 2.438482e-10, 2.448582e-10, 2.457689e-10, 
    2.467625e-10, 2.470057e-10, 2.481679e-10, 2.472213e-10, 2.487831e-10, 
    2.474547e-10, 2.497545e-10, 2.4563e-10, 2.474209e-10, 2.441782e-10, 
    2.445267e-10, 2.451578e-10, 2.466067e-10, 2.458237e-10, 2.467391e-10, 
    2.447183e-10, 2.436709e-10, 2.433998e-10, 2.428948e-10, 2.434108e-10, 
    2.433689e-10, 2.43863e-10, 2.437037e-10, 2.448911e-10, 2.44253e-10, 
    2.460662e-10, 2.467288e-10, 2.486015e-10, 2.497506e-10, 2.509216e-10, 
    2.514385e-10, 2.515959e-10, 2.516615e-10,
  1.335429e-10, 1.345507e-10, 1.343546e-10, 1.351691e-10, 1.34717e-10, 
    1.352507e-10, 1.33747e-10, 1.345908e-10, 1.340519e-10, 1.336335e-10, 
    1.367547e-10, 1.352054e-10, 1.38371e-10, 1.373779e-10, 1.398775e-10, 
    1.382162e-10, 1.402133e-10, 1.398295e-10, 1.40986e-10, 1.406543e-10, 
    1.421371e-10, 1.411391e-10, 1.42908e-10, 1.418986e-10, 1.420563e-10, 
    1.411062e-10, 1.355167e-10, 1.365615e-10, 1.354549e-10, 1.356037e-10, 
    1.355369e-10, 1.347264e-10, 1.343185e-10, 1.33466e-10, 1.336207e-10, 
    1.342469e-10, 1.356706e-10, 1.351867e-10, 1.364075e-10, 1.363799e-10, 
    1.377436e-10, 1.371281e-10, 1.394275e-10, 1.387726e-10, 1.406681e-10, 
    1.401906e-10, 1.406457e-10, 1.405076e-10, 1.406475e-10, 1.399473e-10, 
    1.402471e-10, 1.396316e-10, 1.372433e-10, 1.379437e-10, 1.358587e-10, 
    1.346106e-10, 1.33784e-10, 1.331985e-10, 1.332813e-10, 1.33439e-10, 
    1.342506e-10, 1.350153e-10, 1.355992e-10, 1.359902e-10, 1.363759e-10, 
    1.375458e-10, 1.381666e-10, 1.3956e-10, 1.393082e-10, 1.397349e-10, 
    1.401431e-10, 1.408292e-10, 1.407162e-10, 1.410188e-10, 1.397237e-10, 
    1.405839e-10, 1.391648e-10, 1.395525e-10, 1.364808e-10, 1.353172e-10, 
    1.348237e-10, 1.343923e-10, 1.333449e-10, 1.340679e-10, 1.337827e-10, 
    1.344616e-10, 1.348936e-10, 1.346798e-10, 1.360009e-10, 1.354867e-10, 
    1.382034e-10, 1.370308e-10, 1.400954e-10, 1.393599e-10, 1.40272e-10, 
    1.398063e-10, 1.406045e-10, 1.39886e-10, 1.411315e-10, 1.414032e-10, 
    1.412175e-10, 1.419313e-10, 1.398462e-10, 1.406457e-10, 1.346738e-10, 
    1.347087e-10, 1.348711e-10, 1.341577e-10, 1.341142e-10, 1.334618e-10, 
    1.340422e-10, 1.342897e-10, 1.349186e-10, 1.352911e-10, 1.356456e-10, 
    1.364262e-10, 1.372999e-10, 1.38525e-10, 1.394075e-10, 1.400002e-10, 
    1.396367e-10, 1.399576e-10, 1.395989e-10, 1.394308e-10, 1.413013e-10, 
    1.402499e-10, 1.418286e-10, 1.41741e-10, 1.41026e-10, 1.417509e-10, 
    1.347332e-10, 1.345326e-10, 1.338373e-10, 1.343814e-10, 1.333908e-10, 
    1.339449e-10, 1.342639e-10, 1.354975e-10, 1.357691e-10, 1.360211e-10, 
    1.365193e-10, 1.371596e-10, 1.382855e-10, 1.392679e-10, 1.401668e-10, 
    1.401009e-10, 1.401241e-10, 1.403252e-10, 1.398273e-10, 1.40407e-10, 
    1.405043e-10, 1.402498e-10, 1.417293e-10, 1.413061e-10, 1.417392e-10, 
    1.414635e-10, 1.345978e-10, 1.349353e-10, 1.347529e-10, 1.35096e-10, 
    1.348543e-10, 1.359304e-10, 1.362536e-10, 1.3777e-10, 1.37147e-10, 
    1.38139e-10, 1.372476e-10, 1.374054e-10, 1.381714e-10, 1.372958e-10, 
    1.392136e-10, 1.379123e-10, 1.40333e-10, 1.390297e-10, 1.404148e-10, 
    1.401629e-10, 1.405801e-10, 1.40954e-10, 1.41425e-10, 1.422954e-10, 
    1.420937e-10, 1.428227e-10, 1.354391e-10, 1.358779e-10, 1.358392e-10, 
    1.36299e-10, 1.366394e-10, 1.373782e-10, 1.385661e-10, 1.381189e-10, 
    1.389402e-10, 1.391053e-10, 1.378577e-10, 1.386232e-10, 1.361719e-10, 
    1.365668e-10, 1.363316e-10, 1.354736e-10, 1.382219e-10, 1.36809e-10, 
    1.394221e-10, 1.386537e-10, 1.409007e-10, 1.397815e-10, 1.419827e-10, 
    1.429273e-10, 1.438185e-10, 1.448622e-10, 1.361176e-10, 1.358192e-10, 
    1.363537e-10, 1.370944e-10, 1.377831e-10, 1.387005e-10, 1.387945e-10, 
    1.389667e-10, 1.394129e-10, 1.397886e-10, 1.390211e-10, 1.398828e-10, 
    1.366584e-10, 1.383448e-10, 1.357064e-10, 1.364989e-10, 1.370507e-10, 
    1.368086e-10, 1.380679e-10, 1.383653e-10, 1.395761e-10, 1.389497e-10, 
    1.426939e-10, 1.41033e-10, 1.456588e-10, 1.443608e-10, 1.35715e-10, 
    1.361166e-10, 1.375177e-10, 1.368504e-10, 1.387618e-10, 1.392338e-10, 
    1.396179e-10, 1.401094e-10, 1.401625e-10, 1.404541e-10, 1.399764e-10, 
    1.404352e-10, 1.387025e-10, 1.394758e-10, 1.373573e-10, 1.378718e-10, 
    1.37635e-10, 1.373754e-10, 1.381772e-10, 1.390332e-10, 1.390515e-10, 
    1.393263e-10, 1.401019e-10, 1.387696e-10, 1.429088e-10, 1.403473e-10, 
    1.36555e-10, 1.373306e-10, 1.374416e-10, 1.371409e-10, 1.391864e-10, 
    1.38444e-10, 1.40447e-10, 1.399046e-10, 1.407937e-10, 1.403516e-10, 
    1.402866e-10, 1.397197e-10, 1.393672e-10, 1.38478e-10, 1.37756e-10, 
    1.371845e-10, 1.373173e-10, 1.379454e-10, 1.390856e-10, 1.401673e-10, 
    1.399301e-10, 1.40726e-10, 1.386229e-10, 1.395034e-10, 1.391628e-10, 
    1.400514e-10, 1.381071e-10, 1.397621e-10, 1.376851e-10, 1.378668e-10, 
    1.384293e-10, 1.395631e-10, 1.398145e-10, 1.40083e-10, 1.399173e-10, 
    1.391145e-10, 1.389832e-10, 1.384156e-10, 1.38259e-10, 1.378272e-10, 
    1.374701e-10, 1.377964e-10, 1.381393e-10, 1.391149e-10, 1.399962e-10, 
    1.409593e-10, 1.411954e-10, 1.423243e-10, 1.41405e-10, 1.42923e-10, 
    1.41632e-10, 1.438695e-10, 1.398582e-10, 1.415942e-10, 1.384549e-10, 
    1.387919e-10, 1.394021e-10, 1.408055e-10, 1.400473e-10, 1.409341e-10, 
    1.389781e-10, 1.379671e-10, 1.377059e-10, 1.372192e-10, 1.377171e-10, 
    1.376766e-10, 1.381535e-10, 1.380002e-10, 1.391473e-10, 1.385307e-10, 
    1.40285e-10, 1.409271e-10, 1.427462e-10, 1.438654e-10, 1.450079e-10, 
    1.455133e-10, 1.456672e-10, 1.457316e-10,
  1.249127e-10, 1.260166e-10, 1.258017e-10, 1.266944e-10, 1.261989e-10, 
    1.267839e-10, 1.251362e-10, 1.260605e-10, 1.254701e-10, 1.250119e-10, 
    1.284345e-10, 1.267343e-10, 1.302107e-10, 1.29119e-10, 1.318688e-10, 
    1.300406e-10, 1.322387e-10, 1.318159e-10, 1.330902e-10, 1.327246e-10, 
    1.3436e-10, 1.332591e-10, 1.35211e-10, 1.340967e-10, 1.342708e-10, 
    1.332228e-10, 1.270757e-10, 1.282223e-10, 1.270079e-10, 1.271711e-10, 
    1.270979e-10, 1.262091e-10, 1.257622e-10, 1.248285e-10, 1.249978e-10, 
    1.256837e-10, 1.272445e-10, 1.267138e-10, 1.280532e-10, 1.280229e-10, 
    1.295209e-10, 1.288446e-10, 1.313733e-10, 1.306525e-10, 1.327399e-10, 
    1.322136e-10, 1.327151e-10, 1.32563e-10, 1.327171e-10, 1.319456e-10, 
    1.32276e-10, 1.31598e-10, 1.289712e-10, 1.297408e-10, 1.274509e-10, 
    1.260822e-10, 1.251766e-10, 1.245357e-10, 1.246262e-10, 1.247989e-10, 
    1.256877e-10, 1.265258e-10, 1.271662e-10, 1.275952e-10, 1.280186e-10, 
    1.293036e-10, 1.299859e-10, 1.315192e-10, 1.31242e-10, 1.317118e-10, 
    1.321613e-10, 1.329174e-10, 1.327929e-10, 1.331264e-10, 1.316994e-10, 
    1.326471e-10, 1.310842e-10, 1.315109e-10, 1.281337e-10, 1.268569e-10, 
    1.263158e-10, 1.25843e-10, 1.246958e-10, 1.254876e-10, 1.251752e-10, 
    1.259189e-10, 1.263924e-10, 1.261581e-10, 1.27607e-10, 1.270428e-10, 
    1.300264e-10, 1.287377e-10, 1.321089e-10, 1.312989e-10, 1.323033e-10, 
    1.317904e-10, 1.326698e-10, 1.318782e-10, 1.332506e-10, 1.335503e-10, 
    1.333455e-10, 1.341329e-10, 1.318344e-10, 1.327151e-10, 1.261515e-10, 
    1.261897e-10, 1.263677e-10, 1.25586e-10, 1.255383e-10, 1.248238e-10, 
    1.254595e-10, 1.257305e-10, 1.264199e-10, 1.268283e-10, 1.272171e-10, 
    1.280737e-10, 1.290333e-10, 1.303801e-10, 1.313513e-10, 1.32004e-10, 
    1.316036e-10, 1.319571e-10, 1.31562e-10, 1.31377e-10, 1.33438e-10, 
    1.32279e-10, 1.340195e-10, 1.339229e-10, 1.331343e-10, 1.339338e-10, 
    1.262166e-10, 1.259968e-10, 1.252351e-10, 1.25831e-10, 1.247461e-10, 
    1.253529e-10, 1.257023e-10, 1.270546e-10, 1.273525e-10, 1.27629e-10, 
    1.281759e-10, 1.288792e-10, 1.301168e-10, 1.311976e-10, 1.321875e-10, 
    1.321149e-10, 1.321404e-10, 1.323619e-10, 1.318135e-10, 1.324521e-10, 
    1.325594e-10, 1.322789e-10, 1.3391e-10, 1.334432e-10, 1.339209e-10, 
    1.336168e-10, 1.260682e-10, 1.264382e-10, 1.262382e-10, 1.266143e-10, 
    1.263493e-10, 1.275296e-10, 1.278843e-10, 1.2955e-10, 1.288653e-10, 
    1.299557e-10, 1.289759e-10, 1.291493e-10, 1.299912e-10, 1.290288e-10, 
    1.311379e-10, 1.297064e-10, 1.323706e-10, 1.309354e-10, 1.324607e-10, 
    1.321832e-10, 1.326428e-10, 1.33055e-10, 1.335743e-10, 1.345347e-10, 
    1.34312e-10, 1.351169e-10, 1.269905e-10, 1.274719e-10, 1.274295e-10, 
    1.279341e-10, 1.283078e-10, 1.291193e-10, 1.304253e-10, 1.299336e-10, 
    1.30837e-10, 1.310186e-10, 1.296464e-10, 1.304882e-10, 1.277946e-10, 
    1.282281e-10, 1.279699e-10, 1.270285e-10, 1.300468e-10, 1.28494e-10, 
    1.313674e-10, 1.305217e-10, 1.329962e-10, 1.317631e-10, 1.341895e-10, 
    1.352324e-10, 1.362169e-10, 1.373711e-10, 1.27735e-10, 1.274075e-10, 
    1.279942e-10, 1.288076e-10, 1.295643e-10, 1.305732e-10, 1.306766e-10, 
    1.30866e-10, 1.313572e-10, 1.317708e-10, 1.309259e-10, 1.318746e-10, 
    1.283287e-10, 1.301819e-10, 1.272838e-10, 1.281536e-10, 1.287596e-10, 
    1.284936e-10, 1.298774e-10, 1.302044e-10, 1.315369e-10, 1.308474e-10, 
    1.349747e-10, 1.331421e-10, 1.382527e-10, 1.368165e-10, 1.272932e-10, 
    1.277339e-10, 1.292726e-10, 1.285395e-10, 1.306407e-10, 1.3116e-10, 
    1.315829e-10, 1.321242e-10, 1.321828e-10, 1.32504e-10, 1.319777e-10, 
    1.324832e-10, 1.305754e-10, 1.314265e-10, 1.290964e-10, 1.296619e-10, 
    1.294016e-10, 1.291163e-10, 1.299976e-10, 1.309392e-10, 1.309594e-10, 
    1.312619e-10, 1.32116e-10, 1.306492e-10, 1.352119e-10, 1.323863e-10, 
    1.282152e-10, 1.290671e-10, 1.29189e-10, 1.288586e-10, 1.311079e-10, 
    1.30291e-10, 1.324962e-10, 1.318987e-10, 1.328782e-10, 1.323911e-10, 
    1.323195e-10, 1.316951e-10, 1.313069e-10, 1.303284e-10, 1.295346e-10, 
    1.289065e-10, 1.290524e-10, 1.297427e-10, 1.309969e-10, 1.32188e-10, 
    1.319267e-10, 1.328037e-10, 1.304878e-10, 1.314568e-10, 1.310819e-10, 
    1.320604e-10, 1.299205e-10, 1.317417e-10, 1.294567e-10, 1.296564e-10, 
    1.302748e-10, 1.315226e-10, 1.317994e-10, 1.320952e-10, 1.319126e-10, 
    1.310288e-10, 1.308843e-10, 1.302598e-10, 1.300876e-10, 1.296129e-10, 
    1.292204e-10, 1.295789e-10, 1.29956e-10, 1.310292e-10, 1.319995e-10, 
    1.330609e-10, 1.333211e-10, 1.345666e-10, 1.335523e-10, 1.352277e-10, 
    1.338027e-10, 1.362734e-10, 1.318476e-10, 1.337609e-10, 1.30303e-10, 
    1.306737e-10, 1.313454e-10, 1.328912e-10, 1.320558e-10, 1.330331e-10, 
    1.308786e-10, 1.297666e-10, 1.294795e-10, 1.289446e-10, 1.294918e-10, 
    1.294472e-10, 1.299716e-10, 1.29803e-10, 1.310649e-10, 1.303864e-10, 
    1.323177e-10, 1.330254e-10, 1.350324e-10, 1.362689e-10, 1.375323e-10, 
    1.380916e-10, 1.382621e-10, 1.383333e-10,
  1.281122e-10, 1.293279e-10, 1.290912e-10, 1.300749e-10, 1.295287e-10, 
    1.301735e-10, 1.283583e-10, 1.293763e-10, 1.28726e-10, 1.282214e-10, 
    1.319941e-10, 1.301188e-10, 1.339555e-10, 1.327496e-10, 1.357889e-10, 
    1.337675e-10, 1.361982e-10, 1.357303e-10, 1.371408e-10, 1.36736e-10, 
    1.385476e-10, 1.373278e-10, 1.394912e-10, 1.382558e-10, 1.384488e-10, 
    1.372876e-10, 1.304952e-10, 1.317599e-10, 1.304204e-10, 1.306004e-10, 
    1.305196e-10, 1.2954e-10, 1.290477e-10, 1.280195e-10, 1.282059e-10, 
    1.289612e-10, 1.306813e-10, 1.300962e-10, 1.315733e-10, 1.315398e-10, 
    1.331934e-10, 1.324466e-10, 1.352407e-10, 1.344437e-10, 1.367529e-10, 
    1.361704e-10, 1.367255e-10, 1.36557e-10, 1.367277e-10, 1.358739e-10, 
    1.362394e-10, 1.354892e-10, 1.325863e-10, 1.334364e-10, 1.309089e-10, 
    1.294003e-10, 1.284028e-10, 1.276973e-10, 1.277969e-10, 1.27987e-10, 
    1.289656e-10, 1.29889e-10, 1.305948e-10, 1.31068e-10, 1.31535e-10, 
    1.329535e-10, 1.337072e-10, 1.354021e-10, 1.350955e-10, 1.356152e-10, 
    1.361125e-10, 1.369495e-10, 1.368115e-10, 1.371809e-10, 1.356014e-10, 
    1.366502e-10, 1.349209e-10, 1.353929e-10, 1.316622e-10, 1.302539e-10, 
    1.296576e-10, 1.291367e-10, 1.278736e-10, 1.287452e-10, 1.284013e-10, 
    1.292202e-10, 1.297419e-10, 1.294838e-10, 1.310809e-10, 1.304589e-10, 
    1.337519e-10, 1.323287e-10, 1.360544e-10, 1.351584e-10, 1.362696e-10, 
    1.35702e-10, 1.366753e-10, 1.357992e-10, 1.373185e-10, 1.376503e-10, 
    1.374235e-10, 1.382958e-10, 1.357507e-10, 1.367255e-10, 1.294766e-10, 
    1.295186e-10, 1.297148e-10, 1.288536e-10, 1.288011e-10, 1.280144e-10, 
    1.287142e-10, 1.290128e-10, 1.297722e-10, 1.302224e-10, 1.30651e-10, 
    1.315959e-10, 1.32655e-10, 1.341427e-10, 1.352164e-10, 1.359384e-10, 
    1.354955e-10, 1.358865e-10, 1.354494e-10, 1.352448e-10, 1.375259e-10, 
    1.362428e-10, 1.381702e-10, 1.380632e-10, 1.371897e-10, 1.380753e-10, 
    1.295482e-10, 1.293061e-10, 1.284672e-10, 1.291235e-10, 1.279289e-10, 
    1.285969e-10, 1.289818e-10, 1.304719e-10, 1.308004e-10, 1.311053e-10, 
    1.317086e-10, 1.324848e-10, 1.338517e-10, 1.350464e-10, 1.361415e-10, 
    1.360611e-10, 1.360894e-10, 1.363345e-10, 1.357276e-10, 1.364343e-10, 
    1.365531e-10, 1.362426e-10, 1.380489e-10, 1.375317e-10, 1.380609e-10, 
    1.377241e-10, 1.293848e-10, 1.297924e-10, 1.29572e-10, 1.299865e-10, 
    1.296945e-10, 1.309957e-10, 1.31387e-10, 1.332255e-10, 1.324695e-10, 
    1.336737e-10, 1.325916e-10, 1.32783e-10, 1.337131e-10, 1.326499e-10, 
    1.349804e-10, 1.333983e-10, 1.363441e-10, 1.347566e-10, 1.364439e-10, 
    1.361367e-10, 1.366454e-10, 1.371018e-10, 1.37677e-10, 1.387412e-10, 
    1.384944e-10, 1.393867e-10, 1.304012e-10, 1.309321e-10, 1.308853e-10, 
    1.314418e-10, 1.318541e-10, 1.327499e-10, 1.341926e-10, 1.336492e-10, 
    1.346476e-10, 1.348485e-10, 1.33332e-10, 1.342621e-10, 1.312879e-10, 
    1.317663e-10, 1.314813e-10, 1.304431e-10, 1.337744e-10, 1.320597e-10, 
    1.352342e-10, 1.342991e-10, 1.370367e-10, 1.35672e-10, 1.383587e-10, 
    1.395149e-10, 1.406072e-10, 1.41889e-10, 1.312222e-10, 1.30861e-10, 
    1.315081e-10, 1.324058e-10, 1.332414e-10, 1.343561e-10, 1.344704e-10, 
    1.346798e-10, 1.35223e-10, 1.356804e-10, 1.347461e-10, 1.357952e-10, 
    1.318774e-10, 1.339237e-10, 1.307246e-10, 1.31684e-10, 1.323528e-10, 
    1.320592e-10, 1.335872e-10, 1.339485e-10, 1.354217e-10, 1.346592e-10, 
    1.392291e-10, 1.371983e-10, 1.428686e-10, 1.41273e-10, 1.307349e-10, 
    1.31221e-10, 1.329192e-10, 1.321099e-10, 1.344307e-10, 1.350049e-10, 
    1.354725e-10, 1.360715e-10, 1.361362e-10, 1.364918e-10, 1.359094e-10, 
    1.364687e-10, 1.343585e-10, 1.352995e-10, 1.327245e-10, 1.333491e-10, 
    1.330616e-10, 1.327466e-10, 1.3372e-10, 1.347608e-10, 1.34783e-10, 
    1.351176e-10, 1.360626e-10, 1.344401e-10, 1.394923e-10, 1.363617e-10, 
    1.317519e-10, 1.326923e-10, 1.328269e-10, 1.32462e-10, 1.349473e-10, 
    1.340442e-10, 1.364831e-10, 1.358219e-10, 1.369061e-10, 1.363668e-10, 
    1.362875e-10, 1.355966e-10, 1.351673e-10, 1.340856e-10, 1.332085e-10, 
    1.325149e-10, 1.32676e-10, 1.334384e-10, 1.348245e-10, 1.361421e-10, 
    1.35853e-10, 1.368235e-10, 1.342617e-10, 1.353331e-10, 1.349186e-10, 
    1.360008e-10, 1.336348e-10, 1.356484e-10, 1.331224e-10, 1.33343e-10, 
    1.340263e-10, 1.35406e-10, 1.357121e-10, 1.360393e-10, 1.358373e-10, 
    1.348598e-10, 1.347e-10, 1.340097e-10, 1.338194e-10, 1.332949e-10, 
    1.328615e-10, 1.332575e-10, 1.33674e-10, 1.348602e-10, 1.359335e-10, 
    1.371083e-10, 1.373965e-10, 1.387767e-10, 1.376527e-10, 1.395099e-10, 
    1.379302e-10, 1.406701e-10, 1.357655e-10, 1.378839e-10, 1.340575e-10, 
    1.344672e-10, 1.352099e-10, 1.369205e-10, 1.359957e-10, 1.370776e-10, 
    1.346937e-10, 1.334648e-10, 1.331477e-10, 1.32557e-10, 1.331612e-10, 
    1.33112e-10, 1.336913e-10, 1.33505e-10, 1.348997e-10, 1.341496e-10, 
    1.362856e-10, 1.37069e-10, 1.392931e-10, 1.40665e-10, 1.42068e-10, 
    1.426895e-10, 1.428789e-10, 1.429581e-10,
  1.381729e-10, 1.394607e-10, 1.392098e-10, 1.402524e-10, 1.396735e-10, 
    1.40357e-10, 1.384334e-10, 1.39512e-10, 1.388229e-10, 1.382885e-10, 
    1.422886e-10, 1.40299e-10, 1.443719e-10, 1.430906e-10, 1.463217e-10, 
    1.441721e-10, 1.467573e-10, 1.462593e-10, 1.477609e-10, 1.473298e-10, 
    1.492604e-10, 1.479601e-10, 1.502667e-10, 1.489492e-10, 1.491549e-10, 
    1.479174e-10, 1.40698e-10, 1.4204e-10, 1.406188e-10, 1.408096e-10, 
    1.407239e-10, 1.396854e-10, 1.391638e-10, 1.380747e-10, 1.38272e-10, 
    1.390721e-10, 1.408955e-10, 1.40275e-10, 1.418417e-10, 1.418062e-10, 
    1.43562e-10, 1.427688e-10, 1.457384e-10, 1.448908e-10, 1.473478e-10, 
    1.467277e-10, 1.473187e-10, 1.471393e-10, 1.47321e-10, 1.464121e-10, 
    1.468011e-10, 1.460028e-10, 1.429172e-10, 1.438201e-10, 1.411368e-10, 
    1.395374e-10, 1.384806e-10, 1.377336e-10, 1.37839e-10, 1.380402e-10, 
    1.390768e-10, 1.400553e-10, 1.408037e-10, 1.413056e-10, 1.418011e-10, 
    1.433073e-10, 1.441079e-10, 1.459102e-10, 1.455839e-10, 1.461368e-10, 
    1.46666e-10, 1.475572e-10, 1.474103e-10, 1.478037e-10, 1.461221e-10, 
    1.472385e-10, 1.453982e-10, 1.459002e-10, 1.419363e-10, 1.404422e-10, 
    1.398101e-10, 1.39258e-10, 1.379202e-10, 1.388433e-10, 1.38479e-10, 
    1.393465e-10, 1.398994e-10, 1.396258e-10, 1.413193e-10, 1.406596e-10, 
    1.441555e-10, 1.426436e-10, 1.466043e-10, 1.456508e-10, 1.468333e-10, 
    1.462292e-10, 1.472652e-10, 1.463326e-10, 1.479502e-10, 1.483039e-10, 
    1.480622e-10, 1.489918e-10, 1.46281e-10, 1.473187e-10, 1.396182e-10, 
    1.396628e-10, 1.398706e-10, 1.389582e-10, 1.389024e-10, 1.380693e-10, 
    1.388104e-10, 1.391268e-10, 1.399315e-10, 1.404088e-10, 1.408633e-10, 
    1.418657e-10, 1.429901e-10, 1.445708e-10, 1.457125e-10, 1.464807e-10, 
    1.460094e-10, 1.464255e-10, 1.459604e-10, 1.457427e-10, 1.481713e-10, 
    1.468048e-10, 1.488579e-10, 1.487438e-10, 1.478131e-10, 1.487567e-10, 
    1.396941e-10, 1.394375e-10, 1.385488e-10, 1.39244e-10, 1.379788e-10, 
    1.386862e-10, 1.390939e-10, 1.406734e-10, 1.410217e-10, 1.413452e-10, 
    1.419853e-10, 1.428093e-10, 1.442614e-10, 1.455317e-10, 1.466968e-10, 
    1.466113e-10, 1.466414e-10, 1.469024e-10, 1.462564e-10, 1.470086e-10, 
    1.471351e-10, 1.468046e-10, 1.487286e-10, 1.481774e-10, 1.487414e-10, 
    1.483824e-10, 1.395208e-10, 1.399529e-10, 1.397193e-10, 1.401587e-10, 
    1.398491e-10, 1.412289e-10, 1.416441e-10, 1.435961e-10, 1.427931e-10, 
    1.440723e-10, 1.429227e-10, 1.431261e-10, 1.441143e-10, 1.429847e-10, 
    1.454615e-10, 1.437798e-10, 1.469126e-10, 1.452236e-10, 1.470188e-10, 
    1.466918e-10, 1.472334e-10, 1.477194e-10, 1.483322e-10, 1.494667e-10, 
    1.492036e-10, 1.501552e-10, 1.405984e-10, 1.411614e-10, 1.411118e-10, 
    1.417022e-10, 1.421398e-10, 1.430908e-10, 1.446238e-10, 1.440462e-10, 
    1.451076e-10, 1.453212e-10, 1.437091e-10, 1.446978e-10, 1.415389e-10, 
    1.420466e-10, 1.417442e-10, 1.406428e-10, 1.441793e-10, 1.423581e-10, 
    1.457314e-10, 1.447371e-10, 1.476501e-10, 1.461973e-10, 1.490588e-10, 
    1.502921e-10, 1.514579e-10, 1.528272e-10, 1.414692e-10, 1.41086e-10, 
    1.417725e-10, 1.427255e-10, 1.436129e-10, 1.447976e-10, 1.449191e-10, 
    1.451418e-10, 1.457195e-10, 1.462062e-10, 1.452123e-10, 1.463284e-10, 
    1.421647e-10, 1.44338e-10, 1.409414e-10, 1.419594e-10, 1.426692e-10, 
    1.423575e-10, 1.439803e-10, 1.443643e-10, 1.45931e-10, 1.451198e-10, 
    1.499872e-10, 1.478223e-10, 1.538745e-10, 1.52169e-10, 1.409523e-10, 
    1.414679e-10, 1.432707e-10, 1.424113e-10, 1.448768e-10, 1.454875e-10, 
    1.45985e-10, 1.466224e-10, 1.466913e-10, 1.470698e-10, 1.464498e-10, 
    1.470453e-10, 1.448001e-10, 1.45801e-10, 1.430639e-10, 1.437274e-10, 
    1.434219e-10, 1.430873e-10, 1.441214e-10, 1.452279e-10, 1.452515e-10, 
    1.456074e-10, 1.466132e-10, 1.448869e-10, 1.502682e-10, 1.469316e-10, 
    1.420313e-10, 1.430298e-10, 1.431726e-10, 1.427851e-10, 1.454262e-10, 
    1.444661e-10, 1.470606e-10, 1.463567e-10, 1.475109e-10, 1.469367e-10, 
    1.468524e-10, 1.46117e-10, 1.456603e-10, 1.4451e-10, 1.43578e-10, 
    1.428413e-10, 1.430124e-10, 1.438223e-10, 1.452957e-10, 1.466976e-10, 
    1.463898e-10, 1.47423e-10, 1.446973e-10, 1.458367e-10, 1.453957e-10, 
    1.465472e-10, 1.440309e-10, 1.461724e-10, 1.434865e-10, 1.437208e-10, 
    1.444471e-10, 1.459143e-10, 1.462399e-10, 1.465882e-10, 1.463732e-10, 
    1.453332e-10, 1.451632e-10, 1.444293e-10, 1.442271e-10, 1.436698e-10, 
    1.432093e-10, 1.4363e-10, 1.440726e-10, 1.453336e-10, 1.464756e-10, 
    1.477264e-10, 1.480334e-10, 1.495047e-10, 1.483065e-10, 1.502869e-10, 
    1.486024e-10, 1.515252e-10, 1.462969e-10, 1.485528e-10, 1.444801e-10, 
    1.449157e-10, 1.457056e-10, 1.475265e-10, 1.465417e-10, 1.476937e-10, 
    1.451566e-10, 1.438503e-10, 1.435134e-10, 1.42886e-10, 1.435277e-10, 
    1.434755e-10, 1.440909e-10, 1.438929e-10, 1.453756e-10, 1.445781e-10, 
    1.468503e-10, 1.476846e-10, 1.500553e-10, 1.515196e-10, 1.530184e-10, 
    1.536829e-10, 1.538855e-10, 1.539703e-10,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GC_HEAT1 =
  24532.31, 24552.2, 24548.3, 24564.58, 24555.52, 24566.23, 24536.31, 24553, 
    24542.31, 24534.09, 24596.91, 24565.32, 24630.77, 24609.83, 24662.87, 
    24627.48, 24670.13, 24661.83, 24687.05, 24679.75, 24712.79, 24690.43, 
    24730.39, 24707.41, 24710.97, 24689.71, 24571.61, 24592.93, 24570.35, 
    24573.37, 24572.01, 24555.71, 24547.59, 24530.81, 24533.83, 24546.17, 
    24574.73, 24564.94, 24589.77, 24589.2, 24617.49, 24604.63, 24653.2, 
    24639.29, 24680.05, 24669.63, 24679.56, 24676.54, 24679.6, 24664.37, 
    24670.86, 24657.57, 24607.03, 24621.71, 24578.56, 24553.4, 24537.04, 
    24525.6, 24527.21, 24530.28, 24546.24, 24561.49, 24573.28, 24581.24, 
    24589.12, 24613.35, 24626.42, 24656.04, 24650.65, 24659.79, 24668.6, 
    24683.59, 24681.11, 24687.77, 24659.55, 24678.21, 24647.6, 24655.87, 
    24591.28, 24567.57, 24557.65, 24549.05, 24528.45, 24542.63, 24537.01, 
    24550.43, 24559.05, 24554.77, 24581.46, 24571, 24627.2, 24602.61, 
    24667.57, 24651.75, 24671.4, 24661.33, 24678.66, 24663.05, 24690.27, 
    24696.3, 24692.17, 24708.14, 24662.19, 24679.56, 24554.65, 24555.35, 
    24558.6, 24544.4, 24543.54, 24530.73, 24542.12, 24547.02, 24559.55, 
    24567.04, 24574.22, 24590.15, 24608.21, 24634.05, 24652.77, 24665.51, 
    24657.68, 24664.59, 24656.87, 24653.27, 24694.04, 24670.93, 24705.83, 
    24703.86, 24687.93, 24704.08, 24555.84, 24551.84, 24538.09, 24548.83, 
    24529.34, 24540.2, 24546.51, 24571.21, 24576.73, 24581.87, 24592.06, 
    24605.28, 24628.95, 24649.79, 24669.12, 24667.69, 24668.19, 24672.56, 
    24661.78, 24674.34, 24676.47, 24670.92, 24703.6, 24694.14, 24703.82, 
    24697.65, 24553.14, 24559.88, 24556.23, 24563.11, 24558.26, 24580.02, 
    24586.62, 24618.05, 24605.02, 24625.84, 24607.12, 24610.41, 24626.53, 
    24608.12, 24648.64, 24621.05, 24672.73, 24644.73, 24674.51, 24669.04, 
    24678.12, 24686.34, 24696.79, 24716.38, 24711.81, 24728.43, 24570.03, 
    24578.95, 24578.16, 24587.55, 24594.53, 24609.83, 24634.93, 24625.41, 
    24642.83, 24646.33, 24619.89, 24636.14, 24584.95, 24593.04, 24588.21, 
    24570.73, 24627.6, 24598.03, 24653.08, 24636.78, 24685.17, 24660.8, 
    24709.3, 24730.84, 24751.54, 24776.2, 24583.85, 24577.75, 24588.67, 
    24603.93, 24618.32, 24637.77, 24639.75, 24643.39, 24652.89, 24660.95, 
    24644.54, 24662.98, 24594.93, 24630.21, 24575.46, 24591.64, 24603.03, 
    24598.02, 24624.33, 24630.64, 24656.38, 24643.03, 24725.48, 24688.09, 
    24795.18, 24764.37, 24575.63, 24583.83, 24612.75, 24598.88, 24639.06, 
    24649.06, 24657.28, 24667.88, 24669.03, 24675.37, 24665, 24674.96, 
    24637.81, 24654.23, 24609.4, 24620.19, 24615.21, 24609.78, 24626.64, 
    24644.8, 24645.19, 24651.04, 24667.72, 24639.22, 24730.42, 24673.05, 
    24592.79, 24608.85, 24611.16, 24604.89, 24648.06, 24632.32, 24675.21, 
    24663.45, 24682.81, 24673.14, 24671.72, 24659.46, 24651.91, 24633.04, 
    24617.75, 24605.8, 24608.56, 24621.74, 24645.91, 24669.13, 24664, 
    24681.32, 24636.13, 24654.82, 24647.55, 24666.62, 24625.16, 24660.38, 
    24616.26, 24620.08, 24632, 24656.11, 24661.51, 24667.3, 24663.72, 
    24646.53, 24643.74, 24631.71, 24628.38, 24619.25, 24611.76, 24618.6, 
    24625.84, 24646.54, 24665.43, 24686.46, 24691.68, 24717.04, 24696.35, 
    24730.75, 24701.43, 24752.75, 24662.45, 24700.57, 24632.55, 24639.7, 
    24652.66, 24683.07, 24666.53, 24685.91, 24643.63, 24622.2, 24616.7, 
    24606.52, 24616.93, 24616.08, 24626.14, 24622.9, 24647.22, 24634.17, 
    24671.69, 24685.75, 24726.67, 24752.65, 24779.65, 24791.69, 24795.38, 
    24796.93 ;

 GC_ICE1 =
  17606.52, 17638.29, 17632.06, 17658.06, 17643.58, 17660.69, 17612.91, 
    17639.56, 17622.49, 17609.35, 17709.67, 17659.23, 17763.69, 17730.29, 
    17814.8, 17758.44, 17826.36, 17813.15, 17853.28, 17841.67, 17894.24, 
    17858.67, 17922.23, 17885.67, 17891.33, 17857.51, 17669.28, 17703.32, 
    17667.28, 17672.09, 17669.93, 17643.88, 17630.92, 17604.12, 17608.95, 
    17628.65, 17674.26, 17658.63, 17698.27, 17697.37, 17742.51, 17721.99, 
    17799.41, 17777.27, 17842.15, 17825.57, 17841.37, 17836.56, 17841.43, 
    17817.19, 17827.53, 17806.37, 17725.81, 17749.23, 17680.38, 17640.2, 
    17614.07, 17595.79, 17598.36, 17603.27, 17628.77, 17653.12, 17671.94, 
    17684.66, 17697.24, 17735.89, 17756.76, 17803.93, 17795.36, 17809.91, 
    17823.93, 17847.78, 17843.83, 17854.43, 17809.52, 17839.22, 17790.5, 
    17803.67, 17700.68, 17662.83, 17646.99, 17633.25, 17600.34, 17623, 
    17614.03, 17635.45, 17649.22, 17642.39, 17685.01, 17668.3, 17758, 
    17718.77, 17822.29, 17797.11, 17828.38, 17812.35, 17839.93, 17815.09, 
    17858.4, 17868.01, 17861.44, 17886.84, 17813.72, 17841.37, 17642.2, 
    17643.31, 17648.5, 17625.83, 17624.46, 17603.98, 17622.19, 17630, 
    17650.02, 17661.99, 17673.45, 17698.88, 17727.69, 17768.92, 17798.73, 
    17819.01, 17806.55, 17817.55, 17805.26, 17799.53, 17864.4, 17827.62, 
    17883.16, 17880.03, 17854.69, 17880.38, 17644.1, 17637.71, 17615.74, 
    17632.91, 17601.77, 17619.12, 17629.19, 17668.65, 17677.46, 17685.67, 
    17701.93, 17723.03, 17760.79, 17793.99, 17824.75, 17822.48, 17823.28, 
    17830.23, 17813.07, 17833.06, 17836.45, 17827.62, 17879.61, 17864.57, 
    17879.96, 17870.15, 17639.78, 17650.56, 17644.73, 17655.71, 17647.96, 
    17682.71, 17693.26, 17743.4, 17722.61, 17755.83, 17725.95, 17731.2, 
    17756.93, 17727.55, 17792.15, 17748.18, 17830.5, 17785.94, 17833.34, 
    17824.62, 17839.08, 17852.16, 17868.78, 17899.95, 17892.68, 17919.11, 
    17666.76, 17681, 17679.74, 17694.73, 17705.87, 17730.29, 17770.32, 
    17755.14, 17782.91, 17788.48, 17746.34, 17772.27, 17690.59, 17703.49, 
    17695.8, 17667.88, 17758.63, 17711.45, 17799.23, 17773.28, 17850.29, 
    17811.51, 17888.69, 17922.95, 17955.87, 17995.02, 17688.83, 17679.09, 
    17696.52, 17720.88, 17743.83, 17774.85, 17778.01, 17783.8, 17798.92, 
    17811.74, 17785.64, 17814.98, 17706.5, 17762.79, 17675.42, 17701.27, 
    17719.43, 17711.43, 17753.42, 17763.49, 17804.48, 17783.23, 17914.42, 
    17854.94, 18025.1, 17976.25, 17675.7, 17688.79, 17734.95, 17712.81, 
    17776.91, 17792.83, 17805.9, 17822.77, 17824.6, 17834.7, 17818.19, 
    17834.04, 17774.92, 17801.06, 17729.6, 17746.81, 17738.87, 17730.2, 
    17757.11, 17786.05, 17786.66, 17795.98, 17822.53, 17777.17, 17922.28, 
    17831.01, 17703.1, 17728.72, 17732.41, 17722.41, 17791.23, 17766.16, 
    17834.45, 17815.73, 17846.54, 17831.14, 17828.89, 17809.39, 17797.36, 
    17767.32, 17742.92, 17723.85, 17728.27, 17749.29, 17787.82, 17824.77, 
    17816.6, 17844.17, 17772.25, 17802, 17790.43, 17820.77, 17754.74, 
    17810.85, 17740.54, 17746.64, 17765.66, 17804.04, 17812.63, 17821.86, 
    17816.16, 17788.8, 17784.36, 17765.2, 17759.88, 17745.31, 17733.36, 
    17744.28, 17755.83, 17788.81, 17818.88, 17852.35, 17860.65, 17901, 
    17868.08, 17922.8, 17876.16, 17957.79, 17814.14, 17874.8, 17766.54, 
    17777.92, 17798.55, 17846.96, 17820.63, 17851.46, 17784.19, 17750.02, 
    17741.24, 17725.01, 17741.62, 17740.26, 17756.31, 17751.13, 17789.91, 
    17769.12, 17828.84, 17851.22, 17916.32, 17957.62, 18000.49, 18019.57, 
    18025.42, 18027.87 ;

 GC_LIQ1 =
  5232.788, 5234.817, 5234.419, 5236.08, 5235.155, 5236.248, 5233.196, 
    5234.898, 5233.808, 5232.969, 5239.389, 5236.155, 5242.869, 5240.717, 
    5246.218, 5242.53, 5246.98, 5246.11, 5248.753, 5247.988, 5251.455, 
    5249.108, 5253.304, 5250.889, 5251.263, 5249.032, 5236.797, 5238.98, 
    5236.669, 5236.977, 5236.839, 5235.174, 5234.346, 5232.634, 5232.943, 
    5234.201, 5237.116, 5236.116, 5238.655, 5238.597, 5241.504, 5240.182, 
    5245.206, 5243.751, 5248.02, 5246.928, 5247.969, 5247.652, 5247.973, 
    5246.376, 5247.057, 5245.664, 5240.428, 5241.937, 5237.506, 5234.938, 
    5233.27, 5232.103, 5232.267, 5232.581, 5234.208, 5235.765, 5236.967, 
    5237.781, 5238.589, 5241.078, 5242.422, 5245.503, 5244.939, 5245.896, 
    5246.82, 5248.391, 5248.131, 5248.83, 5245.871, 5247.827, 5244.62, 
    5245.486, 5238.811, 5236.385, 5235.373, 5234.495, 5232.394, 5233.84, 
    5233.267, 5234.635, 5235.515, 5235.079, 5237.803, 5236.735, 5242.502, 
    5239.975, 5246.712, 5245.055, 5247.113, 5246.057, 5247.874, 5246.237, 
    5249.091, 5249.724, 5249.291, 5250.966, 5246.147, 5247.969, 5235.067, 
    5235.138, 5235.469, 5234.021, 5233.933, 5232.626, 5233.788, 5234.288, 
    5235.566, 5236.331, 5237.064, 5238.694, 5240.549, 5243.206, 5245.162, 
    5246.496, 5245.675, 5246.399, 5245.59, 5245.213, 5249.486, 5247.063, 
    5250.723, 5250.517, 5248.846, 5250.54, 5235.188, 5234.78, 5233.376, 
    5234.473, 5232.485, 5233.593, 5234.236, 5236.757, 5237.32, 5237.845, 
    5238.891, 5240.25, 5242.682, 5244.85, 5246.874, 5246.724, 5246.777, 
    5247.235, 5246.104, 5247.421, 5247.645, 5247.063, 5250.489, 5249.497, 
    5250.513, 5249.865, 5234.912, 5235.601, 5235.228, 5235.93, 5235.435, 
    5237.656, 5238.332, 5241.561, 5240.223, 5242.362, 5240.438, 5240.776, 
    5242.433, 5240.541, 5244.729, 5241.87, 5247.252, 5244.32, 5247.439, 
    5246.865, 5247.818, 5248.68, 5249.775, 5251.832, 5251.351, 5253.098, 
    5236.636, 5237.546, 5237.466, 5238.427, 5239.144, 5240.717, 5243.296, 
    5242.318, 5244.122, 5244.488, 5241.75, 5243.422, 5238.161, 5238.991, 
    5238.496, 5236.708, 5242.542, 5239.503, 5245.194, 5243.489, 5248.556, 
    5246.002, 5251.088, 5253.351, 5255.533, 5258.151, 5238.047, 5237.424, 
    5238.542, 5240.11, 5241.589, 5243.592, 5243.799, 5244.18, 5245.173, 
    5246.017, 5244.301, 5246.23, 5239.185, 5242.811, 5237.19, 5238.848, 
    5240.017, 5239.502, 5242.207, 5242.855, 5245.54, 5244.143, 5252.788, 
    5248.863, 5260.196, 5256.885, 5237.208, 5238.044, 5241.017, 5239.591, 
    5243.727, 5244.773, 5245.633, 5246.744, 5246.864, 5247.529, 5246.442, 
    5247.486, 5243.596, 5245.314, 5240.672, 5241.781, 5241.27, 5240.711, 
    5242.445, 5244.328, 5244.368, 5244.98, 5246.728, 5243.744, 5253.307, 
    5247.286, 5238.966, 5240.616, 5240.854, 5240.209, 5244.668, 5243.028, 
    5247.513, 5246.279, 5248.309, 5247.295, 5247.146, 5245.862, 5245.071, 
    5243.103, 5241.531, 5240.302, 5240.586, 5241.941, 5244.444, 5246.875, 
    5246.337, 5248.153, 5243.421, 5245.376, 5244.616, 5246.612, 5242.292, 
    5245.958, 5241.377, 5241.771, 5242.996, 5245.511, 5246.076, 5246.684, 
    5246.308, 5244.508, 5244.217, 5242.966, 5242.624, 5241.685, 5240.915, 
    5241.618, 5242.362, 5244.509, 5246.487, 5248.692, 5249.239, 5251.901, 
    5249.729, 5253.341, 5250.262, 5255.66, 5246.175, 5250.172, 5243.052, 
    5243.793, 5245.15, 5248.337, 5246.603, 5248.634, 5244.205, 5241.988, 
    5241.422, 5240.376, 5241.446, 5241.359, 5242.393, 5242.06, 5244.581, 
    5243.218, 5247.143, 5248.618, 5252.913, 5255.649, 5258.521, 5259.819, 
    5260.218, 5260.385 ;

 GPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GROSS_NMIN =
  8.957596e-09, 8.996981e-09, 8.989325e-09, 9.021091e-09, 9.003469e-09, 
    9.02427e-09, 8.965581e-09, 8.998545e-09, 8.977501e-09, 8.961142e-09, 
    9.082739e-09, 9.022508e-09, 9.145298e-09, 9.106886e-09, 9.203375e-09, 
    9.139321e-09, 9.21629e-09, 9.201526e-09, 9.24596e-09, 9.23323e-09, 
    9.290067e-09, 9.251836e-09, 9.319527e-09, 9.280936e-09, 9.286974e-09, 
    9.250575e-09, 9.034628e-09, 9.075241e-09, 9.032222e-09, 9.038014e-09, 
    9.035415e-09, 9.003833e-09, 8.987919e-09, 8.954586e-09, 8.960638e-09, 
    8.985119e-09, 9.040618e-09, 9.021778e-09, 9.069256e-09, 9.068184e-09, 
    9.121042e-09, 9.09721e-09, 9.186048e-09, 9.160799e-09, 9.233762e-09, 
    9.215412e-09, 9.2329e-09, 9.227597e-09, 9.232969e-09, 9.206058e-09, 
    9.217588e-09, 9.193908e-09, 9.101673e-09, 9.128781e-09, 9.047932e-09, 
    8.99932e-09, 8.967027e-09, 8.944113e-09, 8.947352e-09, 8.953528e-09, 
    8.985262e-09, 9.015098e-09, 9.037835e-09, 9.053045e-09, 9.06803e-09, 
    9.113394e-09, 9.1374e-09, 9.191155e-09, 9.181453e-09, 9.197888e-09, 
    9.213587e-09, 9.239947e-09, 9.235608e-09, 9.247222e-09, 9.197453e-09, 
    9.23053e-09, 9.175927e-09, 9.190861e-09, 9.072108e-09, 9.02686e-09, 
    9.007631e-09, 8.990797e-09, 8.949843e-09, 8.978125e-09, 8.966976e-09, 
    8.993499e-09, 9.010352e-09, 9.002017e-09, 9.05346e-09, 9.033461e-09, 
    9.138823e-09, 9.093441e-09, 9.211756e-09, 9.183444e-09, 9.218542e-09, 
    9.200632e-09, 9.23132e-09, 9.203701e-09, 9.251543e-09, 9.261961e-09, 
    9.254842e-09, 9.282187e-09, 9.202171e-09, 9.232901e-09, 9.001783e-09, 
    9.003143e-09, 9.009476e-09, 8.981637e-09, 8.979933e-09, 8.95442e-09, 
    8.977121e-09, 8.986789e-09, 9.011329e-09, 9.025845e-09, 9.039644e-09, 
    9.069982e-09, 9.103865e-09, 9.151243e-09, 9.185279e-09, 9.208095e-09, 
    9.194104e-09, 9.206456e-09, 9.192648e-09, 9.186177e-09, 9.258057e-09, 
    9.217696e-09, 9.278255e-09, 9.274904e-09, 9.247498e-09, 9.275281e-09, 
    9.004098e-09, 8.996274e-09, 8.969113e-09, 8.990369e-09, 8.951641e-09, 
    8.97332e-09, 8.985785e-09, 9.033879e-09, 9.044445e-09, 9.054244e-09, 
    9.073595e-09, 9.09843e-09, 9.141995e-09, 9.1799e-09, 9.2145e-09, 
    9.211965e-09, 9.212858e-09, 9.220588e-09, 9.20144e-09, 9.223731e-09, 
    9.227473e-09, 9.217691e-09, 9.274455e-09, 9.258238e-09, 9.274832e-09, 
    9.264273e-09, 8.998817e-09, 9.01198e-09, 9.004868e-09, 9.018244e-09, 
    9.00882e-09, 9.050722e-09, 9.063284e-09, 9.122066e-09, 9.097941e-09, 
    9.136334e-09, 9.101841e-09, 9.107954e-09, 9.137589e-09, 9.103704e-09, 
    9.17781e-09, 9.127571e-09, 9.220888e-09, 9.170721e-09, 9.224032e-09, 
    9.214351e-09, 9.230379e-09, 9.244736e-09, 9.262795e-09, 9.296119e-09, 
    9.288402e-09, 9.31627e-09, 9.031604e-09, 9.048678e-09, 9.047175e-09, 
    9.065042e-09, 9.078255e-09, 9.106896e-09, 9.15283e-09, 9.135556e-09, 
    9.167266e-09, 9.173632e-09, 9.125456e-09, 9.155037e-09, 9.060105e-09, 
    9.075444e-09, 9.06631e-09, 9.032951e-09, 9.139538e-09, 9.084839e-09, 
    9.185842e-09, 9.156211e-09, 9.242688e-09, 9.199683e-09, 9.284155e-09, 
    9.320267e-09, 9.354251e-09, 9.393969e-09, 9.057996e-09, 9.046395e-09, 
    9.067167e-09, 9.095906e-09, 9.122569e-09, 9.158018e-09, 9.161645e-09, 
    9.168286e-09, 9.185487e-09, 9.19995e-09, 9.170386e-09, 9.203576e-09, 
    9.079002e-09, 9.144285e-09, 9.042009e-09, 9.072808e-09, 9.094212e-09, 
    9.084822e-09, 9.133582e-09, 9.145074e-09, 9.191774e-09, 9.167632e-09, 
    9.311355e-09, 9.247769e-09, 9.424208e-09, 9.374903e-09, 9.042341e-09, 
    9.057955e-09, 9.112298e-09, 9.086443e-09, 9.160384e-09, 9.178585e-09, 
    9.193379e-09, 9.212294e-09, 9.214335e-09, 9.225541e-09, 9.207178e-09, 
    9.224816e-09, 9.158094e-09, 9.18791e-09, 9.106087e-09, 9.126002e-09, 
    9.11684e-09, 9.10679e-09, 9.137807e-09, 9.170853e-09, 9.171557e-09, 
    9.182153e-09, 9.212014e-09, 9.160684e-09, 9.319565e-09, 9.221447e-09, 
    9.074982e-09, 9.105059e-09, 9.109353e-09, 9.097702e-09, 9.17676e-09, 
    9.148115e-09, 9.225268e-09, 9.204416e-09, 9.238581e-09, 9.221604e-09, 
    9.219106e-09, 9.197302e-09, 9.183726e-09, 9.149429e-09, 9.121522e-09, 
    9.099392e-09, 9.104538e-09, 9.128847e-09, 9.172873e-09, 9.214521e-09, 
    9.205397e-09, 9.235984e-09, 9.155023e-09, 9.188972e-09, 9.175851e-09, 
    9.210064e-09, 9.135097e-09, 9.198939e-09, 9.118779e-09, 9.125807e-09, 
    9.147547e-09, 9.191276e-09, 9.200948e-09, 9.211279e-09, 9.204904e-09, 
    9.17399e-09, 9.168925e-09, 9.147018e-09, 9.14097e-09, 9.124276e-09, 
    9.110457e-09, 9.123084e-09, 9.136345e-09, 9.174003e-09, 9.20794e-09, 
    9.24494e-09, 9.253994e-09, 9.297228e-09, 9.262036e-09, 9.320111e-09, 
    9.270739e-09, 9.356204e-09, 9.202637e-09, 9.269284e-09, 9.148535e-09, 
    9.161544e-09, 9.185073e-09, 9.239038e-09, 9.209903e-09, 9.243975e-09, 
    9.168727e-09, 9.129686e-09, 9.119584e-09, 9.100738e-09, 9.120015e-09, 
    9.118446e-09, 9.136893e-09, 9.130965e-09, 9.175253e-09, 9.151464e-09, 
    9.219044e-09, 9.243706e-09, 9.31335e-09, 9.356044e-09, 9.399502e-09, 
    9.418687e-09, 9.424527e-09, 9.426969e-09 ;

 H2OCAN =
  0.07672504, 0.0767098, 0.0767127, 0.07670052, 0.07670717, 0.07669927, 
    0.07672182, 0.07670932, 0.07671723, 0.07672349, 0.07667714, 0.07669994, 
    0.07665227, 0.07666692, 0.07662957, 0.07665474, 0.07662441, 0.07662998, 
    0.07661238, 0.07661742, 0.07659543, 0.07661005, 0.07658342, 0.07659876, 
    0.07659648, 0.07661058, 0.07669507, 0.07668009, 0.07669602, 0.07669388, 
    0.07669477, 0.07670714, 0.07671355, 0.07672599, 0.07672368, 0.07671443, 
    0.07669291, 0.07670002, 0.07668144, 0.07668184, 0.07666141, 0.07667059, 
    0.07663606, 0.07664583, 0.0766172, 0.07662448, 0.0766176, 0.07661965, 
    0.07661757, 0.07662822, 0.07662369, 0.07663293, 0.07666892, 0.07665848, 
    0.07668996, 0.07670932, 0.07672133, 0.07673005, 0.07672882, 0.07672653, 
    0.07671438, 0.07670262, 0.07669372, 0.07668781, 0.07668191, 0.07666495, 
    0.07665534, 0.07663423, 0.07663778, 0.07663155, 0.07662519, 0.07661485, 
    0.07661651, 0.07661201, 0.07663152, 0.07661867, 0.07663987, 0.07663412, 
    0.07668138, 0.07669806, 0.07670603, 0.07671218, 0.0767279, 0.07671711, 
    0.07672139, 0.07671097, 0.07670448, 0.07670765, 0.07668764, 0.07669548, 
    0.07665477, 0.07667221, 0.07662594, 0.07663703, 0.07662322, 0.07663023, 
    0.07661831, 0.07662904, 0.07661024, 0.07660625, 0.076609, 0.07659806, 
    0.07662966, 0.0766177, 0.07670779, 0.07670728, 0.07670478, 0.07671577, 
    0.07671639, 0.07672611, 0.07671736, 0.07671372, 0.07670402, 0.07669847, 
    0.0766931, 0.07668126, 0.07666822, 0.07664979, 0.07663633, 0.07662731, 
    0.07663277, 0.07662795, 0.07663338, 0.07663587, 0.07660782, 0.07662371, 
    0.07659964, 0.07660093, 0.07661194, 0.07660078, 0.0767069, 0.07670987, 
    0.07672049, 0.07671218, 0.07672714, 0.07671891, 0.07671425, 0.07669555, 
    0.07669117, 0.07668743, 0.07667978, 0.07667012, 0.07665335, 0.07663853, 
    0.07662478, 0.07662576, 0.07662543, 0.07662246, 0.07662997, 0.07662121, 
    0.07661984, 0.07662358, 0.07660112, 0.07660754, 0.07660096, 0.07660513, 
    0.07670888, 0.07670383, 0.07670657, 0.07670147, 0.07670516, 0.07668904, 
    0.0766842, 0.07666128, 0.07667037, 0.0766556, 0.07666878, 0.0766665, 
    0.07665557, 0.076668, 0.07663956, 0.07665927, 0.07662234, 0.07664257, 
    0.07662109, 0.07662484, 0.07661852, 0.07661296, 0.07660575, 0.07659271, 
    0.07659569, 0.07658456, 0.07669619, 0.07668971, 0.07669008, 0.07668313, 
    0.07667803, 0.07666678, 0.07664904, 0.07665566, 0.07664328, 0.07664087, 
    0.07665955, 0.07664827, 0.07668521, 0.07667942, 0.07668272, 0.07669579, 
    0.07665441, 0.0766757, 0.07663614, 0.07664768, 0.07661378, 0.07663091, 
    0.07659738, 0.07658342, 0.07656925, 0.0765537, 0.07668594, 0.07669038, 
    0.07668225, 0.07667136, 0.0766608, 0.07664701, 0.07664549, 0.07664296, 
    0.07663616, 0.07663051, 0.07664236, 0.07662907, 0.07667848, 0.07665247, 
    0.07669224, 0.0766805, 0.07667191, 0.07667546, 0.07665637, 0.07665193, 
    0.07663393, 0.07664313, 0.07658705, 0.07661208, 0.0765411, 0.07656129, 
    0.07669198, 0.07668586, 0.0766649, 0.07667479, 0.07664599, 0.07663896, 
    0.07663305, 0.07662581, 0.07662488, 0.07662055, 0.07662766, 0.07662075, 
    0.07664698, 0.07663527, 0.07666704, 0.07665946, 0.07666288, 0.07666677, 
    0.07665475, 0.07664222, 0.07664163, 0.07663766, 0.076627, 0.07664586, 
    0.07658441, 0.07662313, 0.0766792, 0.07666788, 0.07666589, 0.07667031, 
    0.07663967, 0.07665084, 0.07662061, 0.07662875, 0.0766153, 0.07662202, 
    0.07662303, 0.07663155, 0.07663693, 0.0766504, 0.07666123, 0.07666963, 
    0.07666765, 0.07665841, 0.07664138, 0.07662494, 0.0766286, 0.07661632, 
    0.07664809, 0.076635, 0.07664017, 0.07662659, 0.07665592, 0.07663195, 
    0.07666212, 0.07665942, 0.07665106, 0.07663433, 0.07663012, 0.07662621, 
    0.07662856, 0.07664089, 0.07664275, 0.07665119, 0.07665367, 0.07665998, 
    0.07666535, 0.07666053, 0.07665552, 0.07664075, 0.07662755, 0.07661293, 
    0.07660922, 0.07659282, 0.07660663, 0.07658426, 0.07660397, 0.0765694, 
    0.07663007, 0.07660388, 0.07665057, 0.07664551, 0.07663668, 0.07661557, 
    0.07662665, 0.07661353, 0.0766428, 0.07665826, 0.07666183, 0.07666918, 
    0.07666167, 0.07666226, 0.07665509, 0.07665738, 0.07664026, 0.07664944, 
    0.07662314, 0.07661355, 0.07658584, 0.0765689, 0.07655099, 0.07654322, 
    0.07654082, 0.07653984 ;

 H2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO_TOP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSOI =
  3.85672, 3.869828, 3.867278, 3.877869, 3.871993, 3.878931, 3.859377, 
    3.870348, 3.863343, 3.857902, 3.898485, 3.878343, 3.919517, 3.906602, 
    3.939118, 3.917503, 3.943489, 3.938498, 3.953546, 3.949231, 3.968518, 
    3.955539, 3.978554, 3.965418, 3.967469, 3.955111, 3.882394, 3.895971, 
    3.88159, 3.883523, 3.882657, 3.872113, 3.866805, 3.855723, 3.857734, 
    3.865876, 3.884393, 3.878102, 3.893982, 3.893623, 3.91136, 3.903354, 
    3.933267, 3.924748, 3.949411, 3.943196, 3.949118, 3.947322, 3.949141, 
    3.94003, 3.943931, 3.935923, 3.904851, 3.913961, 3.886841, 3.870601, 
    3.859857, 3.852244, 3.85332, 3.85537, 3.865924, 3.875873, 3.883467, 
    3.888553, 3.893571, 3.908779, 3.916858, 3.934989, 3.931716, 3.937265, 
    3.942578, 3.951505, 3.950036, 3.953972, 3.937122, 3.948313, 3.929852, 
    3.934894, 3.89492, 3.879799, 3.873374, 3.867768, 3.854146, 3.863548, 
    3.859839, 3.868671, 3.874289, 3.87151, 3.888693, 3.882004, 3.917338, 
    3.902086, 3.941958, 3.932388, 3.944255, 3.938197, 3.948581, 3.939235, 
    3.955439, 3.958972, 3.956557, 3.965847, 3.938717, 3.949116, 3.871432, 
    3.871885, 3.873997, 3.864717, 3.86415, 3.855668, 3.863216, 3.866433, 
    3.874616, 3.87946, 3.88407, 3.894223, 3.905585, 3.921523, 3.933008, 
    3.940721, 3.935991, 3.940166, 3.935498, 3.933313, 3.957647, 3.943967, 
    3.96451, 3.963371, 3.954065, 3.9635, 3.872203, 3.869596, 3.860551, 
    3.867628, 3.854745, 3.86195, 3.866097, 3.882141, 3.885677, 3.888953, 
    3.895435, 3.903764, 3.918408, 3.931189, 3.942888, 3.94203, 3.942332, 
    3.944947, 3.93847, 3.946012, 3.947278, 3.943967, 3.963219, 3.957711, 
    3.963347, 3.959761, 3.870444, 3.874833, 3.87246, 3.876921, 3.873777, 
    3.887771, 3.891975, 3.9117, 3.903599, 3.916502, 3.904909, 3.90696, 
    3.916917, 3.905536, 3.930481, 3.913549, 3.945049, 3.928085, 3.946114, 
    3.942837, 3.948265, 3.953129, 3.959258, 3.970582, 3.967959, 3.977446, 
    3.881384, 3.88709, 3.88659, 3.892569, 3.896996, 3.906607, 3.922059, 
    3.916244, 3.926929, 3.929076, 3.912846, 3.922802, 3.890914, 3.896049, 
    3.892993, 3.881833, 3.917579, 3.899199, 3.933197, 3.9232, 3.952435, 
    3.937871, 3.966514, 3.978801, 3.990406, 4.003985, 3.890209, 3.886329, 
    3.893282, 3.902912, 3.911874, 3.923808, 3.925033, 3.927272, 3.933079, 
    3.937966, 3.927977, 3.939192, 3.897234, 3.919179, 3.884861, 3.895165, 
    3.902345, 3.899197, 3.91558, 3.919449, 3.935199, 3.927052, 3.975763, 
    3.954153, 4.014358, 3.99746, 3.884974, 3.890198, 3.908419, 3.899741, 
    3.924608, 3.930747, 3.935746, 3.942139, 3.942832, 3.946624, 3.940411, 
    3.94638, 3.923834, 3.933897, 3.906336, 3.913028, 3.909949, 3.906573, 
    3.917002, 3.928133, 3.928376, 3.93195, 3.942027, 3.924709, 3.978551, 
    3.945222, 3.8959, 3.905984, 3.907432, 3.903521, 3.930131, 3.920472, 
    3.946532, 3.939476, 3.951044, 3.945292, 3.944446, 3.937071, 3.932483, 
    3.920913, 3.911521, 3.904088, 3.905816, 3.913984, 3.928816, 3.942892, 
    3.939805, 3.950164, 3.9228, 3.934253, 3.929822, 3.941386, 3.916088, 
    3.937608, 3.910601, 3.912964, 3.92028, 3.935028, 3.938304, 3.941796, 
    3.939642, 3.929194, 3.927487, 3.920103, 3.918064, 3.91245, 3.907804, 
    3.912048, 3.916507, 3.9292, 3.940666, 3.953198, 3.956271, 3.970951, 
    3.958992, 3.978736, 3.961935, 3.991059, 3.938865, 3.961451, 3.920615, 
    3.924999, 3.932934, 3.951192, 3.941332, 3.952867, 3.92742, 3.914264, 
    3.910872, 3.904539, 3.911016, 3.91049, 3.916695, 3.9147, 3.929623, 
    3.921601, 3.944424, 3.952777, 3.976449, 3.991013, 4.005888, 4.012465, 
    4.01447, 4.015307,
  3.29179, 3.304526, 3.302049, 3.312307, 3.306631, 3.313312, 3.294372, 
    3.305029, 3.298225, 3.292939, 3.331818, 3.312756, 3.351753, 3.33952, 
    3.37033, 3.349842, 3.374475, 3.369747, 3.384017, 3.379924, 3.398208, 
    3.385907, 3.407732, 3.395272, 3.397215, 3.3855, 3.316594, 3.329437, 
    3.315832, 3.317661, 3.316842, 3.306746, 3.301585, 3.290823, 3.292777, 
    3.300685, 3.318484, 3.312531, 3.327569, 3.327229, 3.344028, 3.336445, 
    3.364789, 3.356715, 3.380095, 3.374202, 3.379817, 3.378114, 3.379839, 
    3.371199, 3.374898, 3.367307, 3.337862, 3.346491, 3.320803, 3.305271, 
    3.294837, 3.287443, 3.288488, 3.290478, 3.300731, 3.310401, 3.317612, 
    3.322428, 3.32718, 3.341574, 3.349233, 3.366418, 3.36332, 3.368577, 
    3.373616, 3.38208, 3.380687, 3.384418, 3.368444, 3.379051, 3.361554, 
    3.366331, 3.328441, 3.314138, 3.307966, 3.302524, 3.28929, 3.298423, 
    3.29482, 3.303403, 3.308862, 3.306162, 3.32256, 3.316226, 3.349687, 
    3.335242, 3.373028, 3.363956, 3.375207, 3.369464, 3.379306, 3.370447, 
    3.38581, 3.389159, 3.38687, 3.395682, 3.369956, 3.379813, 3.306085, 
    3.306525, 3.308579, 3.299558, 3.299009, 3.290768, 3.298102, 3.301227, 
    3.309181, 3.313816, 3.318182, 3.327796, 3.338555, 3.353656, 3.364543, 
    3.371856, 3.367373, 3.37133, 3.366905, 3.364834, 3.387902, 3.374931, 
    3.394413, 3.393334, 3.384506, 3.393456, 3.306835, 3.304302, 3.295513, 
    3.30239, 3.289872, 3.296871, 3.300898, 3.316351, 3.319704, 3.322805, 
    3.328944, 3.336832, 3.350705, 3.362818, 3.373911, 3.373098, 3.373384, 
    3.375862, 3.369721, 3.376872, 3.37807, 3.374933, 3.393189, 3.387966, 
    3.393311, 3.38991, 3.305126, 3.30939, 3.307085, 3.311412, 3.308363, 
    3.321681, 3.325662, 3.344346, 3.336675, 3.348898, 3.337918, 3.339859, 
    3.349284, 3.338512, 3.362143, 3.346096, 3.375959, 3.359869, 3.376968, 
    3.373863, 3.379009, 3.38362, 3.389433, 3.400171, 3.397683, 3.406684, 
    3.315639, 3.321038, 3.320569, 3.32623, 3.330421, 3.339527, 3.354166, 
    3.348657, 3.358783, 3.360817, 3.345438, 3.354868, 3.324661, 3.32952, 
    3.32663, 3.316061, 3.349918, 3.332504, 3.364722, 3.355248, 3.382961, 
    3.36915, 3.396313, 3.407963, 3.418983, 3.431864, 3.323995, 3.320322, 
    3.326906, 3.336022, 3.344515, 3.355824, 3.356986, 3.359107, 3.364613, 
    3.369245, 3.359772, 3.370407, 3.330636, 3.351435, 3.318929, 3.328682, 
    3.335487, 3.332506, 3.348029, 3.351694, 3.366619, 3.3589, 3.405079, 
    3.384586, 3.441717, 3.425672, 3.319038, 3.323985, 3.34124, 3.333022, 
    3.356583, 3.3624, 3.367141, 3.373198, 3.373857, 3.377451, 3.371562, 
    3.377221, 3.355848, 3.365386, 3.339271, 3.345609, 3.342694, 3.339495, 
    3.349376, 3.359919, 3.360154, 3.363539, 3.373075, 3.356679, 3.407714, 
    3.376107, 3.329386, 3.338931, 3.340307, 3.336604, 3.361816, 3.352662, 
    3.377365, 3.370677, 3.381644, 3.376189, 3.375387, 3.368396, 3.364046, 
    3.35308, 3.34418, 3.337142, 3.338778, 3.346514, 3.360567, 3.373912, 
    3.370984, 3.380809, 3.35487, 3.365722, 3.361521, 3.372486, 3.348509, 
    3.368889, 3.343312, 3.34555, 3.352481, 3.366453, 3.369565, 3.372873, 
    3.370833, 3.360927, 3.35931, 3.352314, 3.35038, 3.345063, 3.340662, 
    3.344681, 3.348904, 3.360934, 3.371801, 3.383684, 3.3866, 3.400512, 
    3.389171, 3.407889, 3.391951, 3.419588, 3.370087, 3.391501, 3.3528, 
    3.356954, 3.364469, 3.381777, 3.372434, 3.383367, 3.359247, 3.346776, 
    3.343567, 3.337568, 3.343705, 3.343206, 3.349085, 3.347195, 3.361335, 
    3.353734, 3.375365, 3.383283, 3.405736, 3.419553, 3.433677, 3.439922, 
    3.441826, 3.442621,
  3.019155, 3.033256, 3.030511, 3.041911, 3.035584, 3.043054, 3.02201, 
    3.033816, 3.026276, 3.020423, 3.064124, 3.042421, 3.086792, 3.072861, 
    3.107827, 3.08462, 3.1124, 3.107174, 3.122925, 3.118407, 3.138616, 
    3.125012, 3.149131, 3.135364, 3.137514, 3.124564, 3.04678, 3.061416, 
    3.045914, 3.047998, 3.047063, 3.035714, 3.030006, 3.01808, 3.020243, 
    3.029004, 3.048935, 3.042159, 3.059259, 3.058872, 3.07799, 3.069359, 
    3.101623, 3.092428, 3.118595, 3.112091, 3.118289, 3.116409, 3.118314, 
    3.108778, 3.112861, 3.10448, 3.070974, 3.080796, 3.051569, 3.034093, 
    3.022527, 3.014339, 3.015496, 3.017702, 3.029055, 3.039759, 3.047934, 
    3.053412, 3.058816, 3.075216, 3.083924, 3.103484, 3.099948, 3.105887, 
    3.111444, 3.12079, 3.11925, 3.123372, 3.105734, 3.117448, 3.097935, 
    3.103378, 3.060284, 3.043986, 3.037076, 3.031038, 3.016386, 3.026499, 
    3.022509, 3.032008, 3.038054, 3.035063, 3.053562, 3.04636, 3.08444, 
    3.067995, 3.110795, 3.100674, 3.113199, 3.106859, 3.117728, 3.107944, 
    3.124908, 3.12861, 3.12608, 3.13581, 3.107403, 3.118289, 3.034979, 
    3.035467, 3.03774, 3.027756, 3.027146, 3.018021, 3.02614, 3.029602, 
    3.038405, 3.043621, 3.048585, 3.05952, 3.071767, 3.088953, 3.101343, 
    3.109499, 3.10455, 3.108919, 3.10403, 3.10167, 3.127223, 3.112899, 
    3.134409, 3.133216, 3.12347, 3.133351, 3.035809, 3.033003, 3.023274, 
    3.030886, 3.017028, 3.024779, 3.029242, 3.04651, 3.050314, 3.053844, 
    3.060825, 3.069801, 3.085593, 3.099381, 3.111768, 3.11087, 3.111186, 
    3.113924, 3.107144, 3.115038, 3.116364, 3.112898, 3.133057, 3.127287, 
    3.133191, 3.129434, 3.033915, 3.038639, 3.036086, 3.040889, 3.037504, 
    3.052574, 3.057103, 3.07836, 3.069623, 3.083537, 3.071035, 3.073247, 
    3.083991, 3.07171, 3.09862, 3.080356, 3.11403, 3.096037, 3.115145, 
    3.111715, 3.117396, 3.12249, 3.128908, 3.140775, 3.138024, 3.147968, 
    3.045692, 3.051838, 3.051297, 3.057738, 3.062508, 3.072865, 3.08953, 
    3.083256, 3.094781, 3.097099, 3.079591, 3.090332, 3.055957, 3.061491, 
    3.058195, 3.046176, 3.0847, 3.064885, 3.101548, 3.090759, 3.121763, 
    3.106521, 3.136511, 3.149395, 3.161559, 3.175815, 3.055197, 3.051016, 
    3.058505, 3.068887, 3.078544, 3.091416, 3.092736, 3.095152, 3.101419, 
    3.106617, 3.095916, 3.1079, 3.062775, 3.086424, 3.049436, 3.060539, 
    3.068274, 3.06488, 3.082539, 3.086712, 3.10371, 3.094915, 3.14621, 
    3.123565, 3.186704, 3.168965, 3.049556, 3.055182, 3.074821, 3.065465, 
    3.092277, 3.098903, 3.104294, 3.110985, 3.111709, 3.11568, 3.109175, 
    3.115422, 3.091444, 3.102302, 3.072572, 3.079789, 3.076468, 3.072827, 
    3.084073, 3.096086, 3.096343, 3.100203, 3.110881, 3.092386, 3.14914, 
    3.114223, 3.061326, 3.072199, 3.073755, 3.069538, 3.098238, 3.087816, 
    3.115583, 3.108197, 3.120305, 3.114284, 3.113399, 3.10568, 3.100777, 
    3.088294, 3.078164, 3.070149, 3.072011, 3.08082, 3.096822, 3.111774, 
    3.108544, 3.119384, 3.090328, 3.102689, 3.097907, 3.110196, 3.083089, 
    3.106255, 3.07717, 3.079718, 3.08761, 3.103528, 3.106971, 3.110626, 
    3.10837, 3.097229, 3.095385, 3.087418, 3.085221, 3.079164, 3.074155, 
    3.078731, 3.083541, 3.097234, 3.109444, 3.122562, 3.125779, 3.141168, 
    3.128635, 3.149335, 3.131727, 3.162255, 3.107565, 3.131213, 3.08797, 
    3.092699, 3.101267, 3.120465, 3.110139, 3.122218, 3.095313, 3.081124, 
    3.077462, 3.070636, 3.077618, 3.07705, 3.083741, 3.08159, 3.097689, 
    3.089034, 3.113377, 3.122123, 3.146925, 3.1622, 3.177807, 3.184715, 
    3.18682, 3.1877,
  2.8934, 2.908718, 2.905735, 2.918126, 2.911247, 2.919368, 2.8965, 2.909328, 
    2.901133, 2.894776, 2.942291, 2.918679, 2.966968, 2.951795, 2.989996, 
    2.964603, 2.994976, 2.989283, 3.006442, 3.001518, 3.023554, 3.008717, 
    3.035026, 3.020005, 3.022352, 3.008229, 2.923418, 2.939343, 2.922477, 
    2.924743, 2.923726, 2.911389, 2.905188, 2.892231, 2.89458, 2.904098, 
    2.925762, 2.918394, 2.93699, 2.936569, 2.95738, 2.947983, 2.983129, 
    2.973107, 3.001724, 2.994637, 3.001391, 2.999341, 3.001417, 2.991029, 
    2.995476, 2.986253, 2.949741, 2.960436, 2.928627, 2.90963, 2.897062, 
    2.88817, 2.889426, 2.891821, 2.904153, 2.915784, 2.924673, 2.93063, 
    2.936509, 2.954363, 2.963844, 2.985159, 2.981303, 2.987837, 2.993932, 
    3.004115, 3.002437, 3.006931, 2.987664, 3.000475, 2.979108, 2.985042, 
    2.938113, 2.92038, 2.912871, 2.906308, 2.890391, 2.901376, 2.897042, 
    2.90736, 2.913932, 2.91068, 2.930793, 2.922961, 2.964406, 2.946499, 
    2.993226, 2.982094, 2.995845, 2.988929, 3.00078, 2.990121, 3.008604, 
    3.012641, 3.009882, 3.020491, 2.989531, 3.001391, 2.910589, 2.911119, 
    2.91359, 2.902742, 2.90208, 2.892167, 2.900985, 2.904747, 2.914313, 
    2.919983, 2.925381, 2.937276, 2.950605, 2.969321, 2.982823, 2.991814, 
    2.986331, 2.991182, 2.985753, 2.98318, 3.011128, 2.995518, 3.018963, 
    3.017662, 3.007038, 3.017808, 2.911492, 2.908442, 2.897872, 2.906141, 
    2.891089, 2.899508, 2.904357, 2.923126, 2.927261, 2.9311, 2.938694, 
    2.948463, 2.96566, 2.980686, 2.994285, 2.993307, 2.993651, 2.996634, 
    2.989249, 2.997848, 2.999293, 2.995516, 3.017488, 3.011197, 3.017634, 
    3.013537, 2.909433, 2.914567, 2.911792, 2.917013, 2.913334, 2.92972, 
    2.934647, 2.957784, 2.948271, 2.963422, 2.949807, 2.952216, 2.963919, 
    2.950541, 2.979857, 2.959959, 2.99675, 2.977043, 2.997964, 2.994227, 
    3.000416, 3.005968, 3.012964, 3.025908, 3.022906, 3.033756, 2.922235, 
    2.928919, 2.92833, 2.935336, 2.940526, 2.951799, 2.969949, 2.963113, 
    2.975671, 2.978197, 2.959122, 2.970824, 2.933399, 2.939421, 2.935834, 
    2.922762, 2.964689, 2.943115, 2.983047, 2.971288, 3.005176, 2.988552, 
    3.021255, 3.035315, 3.048592, 3.06417, 2.932572, 2.928024, 2.93617, 
    2.94747, 2.957983, 2.972005, 2.973442, 2.976076, 2.982905, 2.988657, 
    2.97691, 2.990072, 2.940821, 2.966567, 2.926307, 2.938386, 2.946803, 
    2.943108, 2.962333, 2.966878, 2.985405, 2.975816, 3.031841, 3.007143, 
    3.076071, 3.056684, 2.926437, 2.932556, 2.95393, 2.943745, 2.972942, 
    2.980164, 2.986043, 2.993434, 2.994221, 2.998547, 2.991461, 2.998267, 
    2.972035, 2.983869, 2.95148, 2.959338, 2.955721, 2.951757, 2.964003, 
    2.977094, 2.977373, 2.981581, 2.993328, 2.973061, 3.035043, 2.996968, 
    2.939239, 2.951076, 2.952768, 2.948176, 2.979439, 2.968082, 2.998441, 
    2.990396, 3.003587, 2.997027, 2.996063, 2.987603, 2.982206, 2.968602, 
    2.957569, 2.948842, 2.950869, 2.960462, 2.977896, 2.994293, 2.990775, 
    3.002583, 2.970818, 2.984291, 2.979079, 2.992573, 2.962932, 2.988258, 
    2.956486, 2.959261, 2.967857, 2.985208, 2.989055, 2.993042, 2.990584, 
    2.97834, 2.976329, 2.967648, 2.965255, 2.958656, 2.953203, 2.958185, 
    2.963426, 2.978344, 2.991755, 3.006048, 3.009553, 3.02634, 3.012671, 
    3.035256, 3.016048, 3.049358, 2.989712, 3.015482, 2.968248, 2.973402, 
    2.982742, 3.003765, 2.992512, 3.005675, 2.97625, 2.960794, 2.956804, 
    2.949372, 2.956974, 2.956355, 2.963642, 2.961298, 2.978841, 2.969408, 
    2.996038, 3.00557, 3.032618, 3.049294, 3.066343, 3.073895, 3.076196, 
    3.077159,
  2.944195, 2.960306, 2.957167, 2.970212, 2.962968, 2.97152, 2.947453, 
    2.960948, 2.952326, 2.945641, 2.995688, 2.970795, 3.021753, 3.00572, 
    3.04615, 3.019253, 3.051601, 3.045369, 3.064159, 3.058765, 3.082828, 
    3.066653, 3.095021, 3.079031, 3.08155, 3.066117, 2.975787, 2.992578, 
    2.974795, 2.977183, 2.976111, 2.963118, 2.956593, 2.942966, 2.945435, 
    2.955445, 2.978258, 2.970494, 2.990095, 2.989651, 3.011619, 3.001695, 
    3.03885, 3.028244, 3.05899, 3.051229, 3.058625, 3.05638, 3.058654, 
    3.047281, 3.052149, 3.042158, 3.003551, 3.014848, 2.981277, 2.961267, 
    2.948044, 2.938697, 2.940017, 2.942534, 2.955503, 2.967746, 2.977109, 
    2.983388, 2.989587, 3.008432, 3.01845, 3.041, 3.036917, 3.043836, 
    3.050458, 3.06161, 3.059772, 3.064695, 3.043652, 3.057622, 3.034594, 
    3.040876, 2.99128, 2.972586, 2.964679, 2.957771, 2.941032, 2.952582, 
    2.948024, 2.958878, 2.965795, 2.962372, 2.98356, 2.975306, 3.019045, 
    3.000129, 3.049685, 3.037755, 3.052551, 3.044992, 3.057956, 3.046286, 
    3.066529, 3.070955, 3.06793, 3.079564, 3.04564, 3.058625, 2.962276, 
    2.962834, 2.965435, 2.954019, 2.953322, 2.942898, 2.952171, 2.956129, 
    2.966197, 2.972168, 2.977855, 2.990396, 3.004464, 3.024241, 3.038527, 
    3.048139, 3.042241, 3.047448, 3.041628, 3.038904, 3.069296, 3.052194, 
    3.077888, 3.07646, 3.064812, 3.076621, 2.963226, 2.960016, 2.948897, 
    2.957595, 2.941765, 2.950616, 2.955718, 2.975479, 2.979836, 2.983884, 
    2.991893, 3.002202, 3.02037, 3.036264, 3.050844, 3.049773, 3.05015, 
    3.053416, 3.045333, 3.054745, 3.056328, 3.052192, 3.076269, 3.069371, 
    3.07643, 3.071937, 2.961059, 2.966465, 2.963542, 2.96904, 2.965166, 
    2.98243, 2.987624, 3.012047, 3.001999, 3.018004, 3.003621, 3.006165, 
    3.01853, 3.004396, 3.035387, 3.014344, 3.053543, 3.03241, 3.054872, 
    3.050781, 3.057558, 3.06364, 3.071309, 3.085328, 3.082139, 3.09367, 
    2.97454, 2.981585, 2.980963, 2.98835, 2.993825, 3.005724, 3.024905, 
    3.017678, 3.030957, 3.03363, 3.01346, 3.02583, 2.986308, 2.99266, 
    2.988876, 2.975096, 3.019343, 2.996557, 3.038763, 3.026321, 3.062773, 
    3.044593, 3.080385, 3.095329, 3.109456, 3.126053, 2.985435, 2.980641, 
    2.98923, 3.001154, 3.012256, 3.027079, 3.028599, 3.031385, 3.038613, 
    3.044704, 3.032268, 3.046233, 2.994137, 3.021328, 2.978831, 2.991568, 
    3.000449, 2.996549, 3.016852, 3.021657, 3.04126, 3.031111, 3.091635, 
    3.064928, 3.138747, 3.118074, 2.978968, 2.985418, 3.007975, 2.997222, 
    3.02807, 3.035711, 3.041936, 3.049912, 3.050774, 3.055511, 3.047753, 
    3.055204, 3.027111, 3.039633, 3.005387, 3.013688, 3.009866, 3.00568, 
    3.018618, 3.032464, 3.032758, 3.037212, 3.049798, 3.028196, 3.09504, 
    3.053783, 2.992467, 3.004961, 3.006747, 3.001899, 3.034945, 3.022931, 
    3.055395, 3.046587, 3.061031, 3.053846, 3.05279, 3.043588, 3.037873, 
    3.023481, 3.011819, 3.002602, 3.004742, 3.014876, 3.033312, 3.050853, 
    3.047002, 3.059931, 3.025823, 3.040081, 3.034563, 3.048971, 3.017486, 
    3.044282, 3.010674, 3.013606, 3.022693, 3.041052, 3.045125, 3.049484, 
    3.046793, 3.033781, 3.031654, 3.022471, 3.019941, 3.012968, 3.007206, 
    3.01247, 3.018008, 3.033786, 3.048075, 3.063727, 3.067569, 3.085788, 
    3.070988, 3.095267, 3.074692, 3.110272, 3.04584, 3.074071, 3.023106, 
    3.028557, 3.038441, 3.061226, 3.048903, 3.063319, 3.03157, 3.015227, 
    3.01101, 3.003162, 3.01119, 3.010536, 3.018236, 3.015759, 3.034311, 
    3.024332, 3.052764, 3.063205, 3.09246, 3.110204, 3.12837, 3.136424, 
    3.13888, 3.139907,
  2.969919, 2.988319, 2.984731, 2.999652, 2.991363, 3.001151, 2.973637, 
    2.989053, 2.9792, 2.971568, 3.028875, 3.00032, 3.058885, 3.040413, 
    3.087081, 3.056003, 3.093395, 3.086177, 3.10796, 3.1017, 3.129779, 
    3.110855, 3.144458, 3.125246, 3.128242, 3.110234, 3.006038, 3.025302, 
    3.004902, 3.007638, 3.00641, 2.991535, 2.984074, 2.968517, 2.971334, 
    2.982763, 3.00887, 2.999975, 3.02245, 3.021941, 3.047204, 3.035781, 
    3.078634, 3.066377, 3.101961, 3.092964, 3.101538, 3.098935, 3.101572, 
    3.08839, 3.094029, 3.082461, 3.037916, 3.050925, 3.012331, 2.989418, 
    2.974312, 2.96365, 2.965154, 2.968025, 2.98283, 2.99683, 3.007553, 
    3.014753, 3.021867, 3.043535, 3.055076, 3.08112, 3.076398, 3.084402, 
    3.092071, 3.105001, 3.102868, 3.108582, 3.084189, 3.100375, 3.073713, 
    3.080977, 3.023812, 3.002371, 2.99332, 2.98542, 2.966312, 2.979492, 
    2.974288, 2.986686, 2.994597, 2.990681, 3.01495, 3.005486, 3.055762, 
    3.03398, 3.091175, 3.077367, 3.094496, 3.08574, 3.100762, 3.087238, 
    3.110712, 3.115854, 3.112339, 3.125865, 3.086491, 3.101539, 2.990571, 
    2.99121, 2.994185, 2.981134, 2.980337, 2.96844, 2.979023, 2.983544, 
    2.995056, 3.001892, 3.008408, 3.022796, 3.038966, 3.061756, 3.078259, 
    3.089385, 3.082556, 3.088584, 3.081847, 3.078696, 3.113926, 3.094082, 
    3.123915, 3.122255, 3.108718, 3.122442, 2.991658, 2.987987, 2.975284, 
    2.985219, 2.967148, 2.977248, 2.983075, 3.005685, 3.010679, 3.015322, 
    3.024515, 3.036364, 3.057291, 3.075644, 3.092517, 3.091277, 3.091713, 
    3.095498, 3.086135, 3.097039, 3.098874, 3.094079, 3.122032, 3.114014, 
    3.12222, 3.116995, 2.989179, 2.995363, 2.99202, 2.998311, 2.993877, 
    3.013653, 3.019614, 3.047697, 3.036131, 3.054562, 3.037996, 3.040924, 
    3.055168, 3.038888, 3.07463, 3.050344, 3.095645, 3.071189, 3.097186, 
    3.092444, 3.1003, 3.107358, 3.116265, 3.132787, 3.128951, 3.14283, 
    3.00461, 3.012685, 3.011971, 3.020447, 3.026735, 3.040416, 3.062522, 
    3.054186, 3.069511, 3.072599, 3.049325, 3.06359, 3.018103, 3.025396, 
    3.02105, 3.005246, 3.056106, 3.029874, 3.078533, 3.064157, 3.106351, 
    3.085278, 3.126842, 3.14483, 3.161399, 3.180833, 3.017102, 3.011602, 
    3.021457, 3.035159, 3.047937, 3.065032, 3.066787, 3.070005, 3.07836, 
    3.085407, 3.071025, 3.087177, 3.027093, 3.058396, 3.009527, 3.024142, 
    3.034348, 3.029865, 3.053234, 3.058775, 3.081422, 3.069688, 3.140379, 
    3.108853, 3.195733, 3.171485, 3.009684, 3.017082, 3.043007, 3.030638, 
    3.066177, 3.075005, 3.082203, 3.091438, 3.092436, 3.097927, 3.088937, 
    3.09757, 3.065068, 3.07954, 3.040029, 3.049588, 3.045185, 3.040366, 
    3.05527, 3.071251, 3.071592, 3.076739, 3.091306, 3.066322, 3.144481, 
    3.095923, 3.025175, 3.039538, 3.041594, 3.036016, 3.074118, 3.060244, 
    3.097792, 3.087587, 3.10433, 3.095996, 3.094772, 3.084115, 3.077504, 
    3.060879, 3.047434, 3.036824, 3.039287, 3.050956, 3.072232, 3.092528, 
    3.088068, 3.103053, 3.063582, 3.080057, 3.073677, 3.090347, 3.053965, 
    3.084919, 3.046116, 3.049493, 3.05997, 3.08118, 3.085895, 3.090942, 
    3.087826, 3.072774, 3.070316, 3.059714, 3.056796, 3.048757, 3.042123, 
    3.048184, 3.054566, 3.072779, 3.08931, 3.107459, 3.11192, 3.133341, 
    3.115892, 3.144755, 3.120199, 3.162355, 3.086721, 3.119477, 3.060447, 
    3.066738, 3.078161, 3.104556, 3.090269, 3.106985, 3.070219, 3.051361, 
    3.046503, 3.037468, 3.04671, 3.045957, 3.05483, 3.051975, 3.073386, 
    3.061862, 3.094742, 3.106852, 3.141372, 3.162275, 3.18355, 3.193005, 
    3.195889, 3.197097,
  3.25474, 3.278216, 3.273628, 3.292736, 3.282112, 3.294659, 3.259475, 
    3.279155, 3.266567, 3.25684, 3.329905, 3.293593, 3.36768, 3.344389, 
    3.403475, 3.364037, 3.411532, 3.402323, 3.430178, 3.422154, 3.458264, 
    3.433893, 3.477266, 3.452412, 3.456279, 3.433096, 3.300937, 3.32543, 
    3.299477, 3.302995, 3.301415, 3.282331, 3.272789, 3.252956, 3.256541, 
    3.271114, 3.304579, 3.29315, 3.321861, 3.321223, 3.352937, 3.338568, 
    3.39272, 3.377162, 3.422488, 3.410982, 3.421946, 3.418614, 3.42199, 
    3.405144, 3.412343, 3.397589, 3.341251, 3.357627, 3.309035, 3.279622, 
    3.260334, 3.246769, 3.248681, 3.252331, 3.2712, 3.289115, 3.302885, 
    3.312154, 3.321131, 3.348316, 3.362867, 3.395883, 3.389878, 3.400062, 
    3.409841, 3.426383, 3.42365, 3.430976, 3.399791, 3.420457, 3.386467, 
    3.3957, 3.323564, 3.296226, 3.284618, 3.27451, 3.250152, 3.266939, 
    3.260304, 3.276128, 3.286254, 3.281238, 3.312408, 3.300228, 3.363733, 
    3.336308, 3.408698, 3.391109, 3.412939, 3.401766, 3.420953, 3.403676, 
    3.433709, 3.440316, 3.435799, 3.453212, 3.402723, 3.421947, 3.281098, 
    3.281915, 3.285726, 3.269035, 3.268018, 3.252858, 3.26634, 3.272112, 
    3.286842, 3.295611, 3.303986, 3.322293, 3.342571, 3.371311, 3.392244, 
    3.406413, 3.397711, 3.405391, 3.396808, 3.392798, 3.437838, 3.41241, 
    3.450697, 3.448557, 3.43115, 3.448798, 3.282489, 3.277791, 3.261574, 
    3.274253, 3.251215, 3.264076, 3.271513, 3.300484, 3.306908, 3.312887, 
    3.324444, 3.339301, 3.365664, 3.388919, 3.410411, 3.408828, 3.409385, 
    3.41422, 3.402269, 3.416189, 3.418537, 3.412406, 3.44827, 3.437951, 
    3.448511, 3.441785, 3.279317, 3.287235, 3.282952, 3.291014, 3.285331, 
    3.310737, 3.318314, 3.353558, 3.339008, 3.362218, 3.341351, 3.345032, 
    3.362983, 3.342472, 3.387631, 3.356895, 3.414408, 3.383263, 3.416378, 
    3.410318, 3.420361, 3.429405, 3.440845, 3.46215, 3.457194, 3.475154, 
    3.299102, 3.30949, 3.308571, 3.319355, 3.327223, 3.344393, 3.37228, 
    3.361742, 3.381134, 3.385053, 3.35561, 3.373632, 3.316426, 3.325547, 
    3.32011, 3.29992, 3.364168, 3.331157, 3.392592, 3.37435, 3.428113, 
    3.401177, 3.454472, 3.477748, 3.499923, 3.526196, 3.315175, 3.308096, 
    3.320618, 3.337787, 3.353861, 3.375458, 3.377681, 3.381761, 3.392371, 
    3.401342, 3.383055, 3.403597, 3.327673, 3.367061, 3.305425, 3.323977, 
    3.33677, 3.331146, 3.360542, 3.367541, 3.396266, 3.381359, 3.471977, 
    3.431324, 3.546063, 3.513536, 3.305627, 3.31515, 3.347653, 3.332115, 
    3.376908, 3.388107, 3.397261, 3.409034, 3.410308, 3.417325, 3.405841, 
    3.416869, 3.375504, 3.393872, 3.343906, 3.355941, 3.350394, 3.34433, 
    3.363112, 3.383342, 3.383774, 3.390311, 3.408866, 3.377091, 3.477296, 
    3.414763, 3.32527, 3.34329, 3.345875, 3.338864, 3.386981, 3.369398, 
    3.417153, 3.404121, 3.425522, 3.414856, 3.413292, 3.399696, 3.391283, 
    3.370201, 3.353227, 3.339879, 3.342974, 3.357667, 3.384586, 3.410425, 
    3.404733, 3.423887, 3.373622, 3.394531, 3.386421, 3.407641, 3.361464, 
    3.40072, 3.351566, 3.355822, 3.369051, 3.395959, 3.401963, 3.408401, 
    3.404425, 3.385274, 3.382155, 3.368728, 3.365039, 3.354895, 3.34654, 
    3.354172, 3.362223, 3.385281, 3.406317, 3.429534, 3.435261, 3.462866, 
    3.440366, 3.477651, 3.445909, 3.501211, 3.403017, 3.444978, 3.369654, 
    3.377619, 3.392118, 3.425813, 3.407541, 3.428927, 3.382033, 3.358178, 
    3.352053, 3.340688, 3.352314, 3.351366, 3.362556, 3.358952, 3.386052, 
    3.371444, 3.413254, 3.428756, 3.473264, 3.501102, 3.529882, 3.542461, 
    3.54627, 3.547865,
  3.812393, 3.852924, 3.844952, 3.878324, 3.859713, 3.881707, 3.820515, 
    3.854559, 3.83273, 3.815992, 3.945428, 3.879831, 4.016907, 3.972589, 
    4.084889, 4.009922, 4.100391, 4.08268, 4.136661, 4.120984, 4.192374, 
    4.143956, 4.230835, 4.180657, 4.188393, 4.142387, 3.892786, 3.937095, 
    3.890205, 3.896428, 3.893631, 3.860096, 3.843497, 3.80934, 3.815479, 
    3.840594, 3.899235, 3.879052, 3.93047, 3.929288, 3.988761, 3.961638, 
    4.064354, 4.034963, 4.121634, 4.099329, 4.12058, 4.114101, 4.120664, 
    4.088093, 4.101956, 4.073629, 3.96668, 3.997681, 3.907147, 3.855371, 
    3.821991, 3.798779, 3.802038, 3.808271, 3.840742, 3.871965, 3.896233, 
    3.912702, 3.929118, 3.980006, 4.007683, 4.070376, 4.058958, 4.078353, 
    4.097129, 4.129234, 4.123899, 4.138225, 4.077835, 4.117682, 4.052496, 
    4.070027, 3.933629, 3.884468, 3.86409, 3.846481, 3.804549, 3.833373, 
    3.82194, 3.849291, 3.866952, 3.858189, 3.913155, 3.891532, 4.00934, 
    3.957397, 4.094926, 4.061294, 4.103108, 4.081614, 4.118647, 4.085274, 
    4.143593, 4.15662, 4.147705, 4.182254, 4.083448, 4.120581, 3.857945, 
    3.85937, 3.866028, 3.836994, 3.835237, 3.809173, 3.832339, 3.842322, 
    3.867982, 3.883384, 3.898182, 3.931272, 3.969163, 4.023889, 4.06345, 
    4.09053, 4.073862, 4.088568, 4.072139, 4.064504, 4.151726, 4.102087, 
    4.177233, 4.172968, 4.138568, 4.173448, 3.860372, 3.852184, 3.824124, 
    3.846035, 3.806363, 3.828434, 3.841284, 3.891984, 3.903368, 3.91401, 
    3.935263, 3.963014, 4.01304, 4.05714, 4.098228, 4.095177, 4.096251, 
    4.105585, 4.082578, 4.109397, 4.113951, 4.102079, 4.172398, 4.151948, 
    4.172878, 4.159524, 3.85484, 3.86867, 3.86118, 3.875299, 3.865339, 
    3.910178, 3.923903, 3.989941, 3.962463, 4.006441, 3.966868, 3.973802, 
    4.007906, 3.968978, 4.0547, 3.996286, 4.105948, 4.046445, 4.109763, 
    4.098048, 4.117496, 4.135146, 4.157666, 4.200188, 4.190227, 4.226528, 
    3.889542, 3.907957, 3.906323, 3.92583, 3.940431, 3.972598, 4.025756, 
    4.005533, 4.042431, 4.049824, 3.99384, 4.028343, 3.920414, 3.937314, 
    3.927225, 3.890987, 4.010172, 3.947763, 4.064112, 4.029688, 4.132617, 
    4.080487, 4.184773, 4.231818, 4.277538, 4.332246, 3.918106, 3.905478, 
    3.928166, 3.960172, 3.990517, 4.031764, 4.035937, 4.043613, 4.063693, 
    4.080802, 4.046052, 4.085124, 3.941267, 4.015718, 3.900735, 3.934397, 
    3.958264, 3.947742, 4.003239, 4.01664, 4.071107, 4.042855, 4.220065, 
    4.138907, 4.374605, 4.306057, 3.901093, 3.918061, 3.978752, 3.949552, 
    4.034485, 4.055602, 4.073004, 4.095573, 4.09803, 4.111598, 4.089432, 
    4.110715, 4.031851, 4.066545, 3.971679, 3.994471, 3.983939, 3.972478, 
    4.008152, 4.046594, 4.047409, 4.05978, 4.09525, 4.03483, 4.230896, 
    4.106637, 3.936798, 3.970517, 3.975393, 3.962193, 4.053471, 4.020208, 
    4.111266, 4.086128, 4.127552, 4.106816, 4.103791, 4.077653, 4.061625, 
    4.021753, 3.989313, 3.964099, 3.969922, 3.997757, 4.048943, 4.098255, 
    4.087304, 4.124361, 4.028325, 4.067799, 4.052412, 4.092893, 4.005001, 
    4.079612, 3.986161, 3.994245, 4.019541, 4.070521, 4.081992, 4.094354, 
    4.086712, 4.050242, 4.044355, 4.018919, 4.011842, 3.99248, 3.976649, 
    3.991108, 4.006452, 4.050256, 4.090347, 4.1354, 4.146646, 4.201631, 
    4.156718, 4.231621, 4.167703, 4.280221, 4.084012, 4.165855, 4.020701, 
    4.03582, 4.06321, 4.128119, 4.0927, 4.134209, 4.044125, 3.99873, 
    3.987085, 3.965621, 3.98758, 3.985781, 4.007088, 4.000206, 4.051713, 
    4.024145, 4.103716, 4.133875, 4.222682, 4.279996, 4.339895, 4.366773, 
    4.375056, 4.378533,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HC =
  24814.35, 24834.79, 24830.78, 24847.51, 24838.19, 24849.2, 24818.46, 
    24835.61, 24824.62, 24816.17, 24880.72, 24848.26, 24915.51, 24894, 
    24948.5, 24912.13, 24955.97, 24947.43, 24973.35, 24965.85, 24999.81, 
    24976.83, 25017.9, 24994.28, 24997.93, 24976.08, 24854.72, 24876.64, 
    24853.44, 24856.54, 24855.14, 24838.38, 24830.05, 24812.81, 24815.91, 
    24828.59, 24857.93, 24847.87, 24873.38, 24872.8, 24901.87, 24888.66, 
    24938.56, 24924.27, 24966.16, 24955.46, 24965.66, 24962.55, 24965.7, 
    24950.04, 24956.72, 24943.06, 24891.12, 24906.2, 24861.87, 24836.01, 
    24819.21, 24807.45, 24809.1, 24812.26, 24828.66, 24844.33, 24856.44, 
    24864.62, 24872.72, 24897.61, 24911.05, 24941.48, 24935.95, 24945.34, 
    24954.4, 24969.8, 24967.25, 24974.1, 24945.09, 24964.27, 24932.81, 
    24941.31, 24874.94, 24850.57, 24840.39, 24831.55, 24810.38, 24824.95, 
    24819.18, 24832.96, 24841.82, 24837.43, 24864.85, 24854.1, 24911.85, 
    24886.58, 24953.34, 24937.08, 24957.27, 24946.92, 24964.73, 24948.69, 
    24976.66, 24982.87, 24978.62, 24995.03, 24947.8, 24965.66, 24837.31, 
    24838.02, 24841.36, 24826.77, 24825.89, 24812.72, 24824.43, 24829.46, 
    24842.34, 24850.04, 24857.41, 24873.78, 24892.33, 24918.88, 24938.12, 
    24951.22, 24943.17, 24950.27, 24942.34, 24938.64, 24980.54, 24956.78, 
    24992.65, 24990.63, 24974.26, 24990.86, 24838.52, 24834.41, 24820.28, 
    24831.32, 24811.3, 24822.46, 24828.93, 24854.32, 24859.99, 24865.27, 
    24875.74, 24889.33, 24913.64, 24935.06, 24954.93, 24953.46, 24953.97, 
    24958.46, 24947.38, 24960.29, 24962.48, 24956.78, 24990.36, 24980.64, 
    24990.59, 24984.25, 24835.75, 24842.68, 24838.93, 24846, 24841.01, 
    24863.37, 24870.15, 24902.44, 24889.06, 24910.45, 24891.21, 24894.59, 
    24911.16, 24892.24, 24933.88, 24905.52, 24958.64, 24929.86, 24960.47, 
    24954.84, 24964.18, 24972.63, 24983.36, 25003.5, 24998.8, 25015.88, 
    24853.11, 24862.27, 24861.46, 24871.1, 24878.28, 24894, 24919.79, 
    24910.01, 24927.91, 24931.51, 24904.34, 24921.04, 24868.44, 24876.74, 
    24871.79, 24853.83, 24912.25, 24881.87, 24938.45, 24921.69, 24971.42, 
    24946.38, 24996.22, 25018.36, 25039.64, 25064.98, 24867.3, 24861.04, 
    24872.25, 24887.94, 24902.72, 24922.71, 24924.74, 24928.48, 24938.24, 
    24946.53, 24929.67, 24948.61, 24878.68, 24914.94, 24858.68, 24875.31, 
    24887.01, 24881.86, 24908.9, 24915.38, 24941.84, 24928.12, 25012.85, 
    24974.42, 25084.49, 25052.82, 24858.86, 24867.28, 24897, 24882.74, 
    24924.04, 24934.32, 24942.76, 24953.65, 24954.83, 24961.35, 24950.69, 
    24960.93, 24922.75, 24939.63, 24893.56, 24904.64, 24899.53, 24893.95, 
    24911.28, 24929.94, 24930.33, 24936.35, 24953.49, 24924.2, 25017.93, 
    24958.97, 24876.49, 24892.99, 24895.37, 24888.93, 24933.28, 24917.11, 
    24961.19, 24949.1, 24969, 24959.05, 24957.6, 24945.01, 24937.24, 
    24917.85, 24902.14, 24889.86, 24892.7, 24906.24, 24931.08, 24954.94, 
    24949.66, 24967.47, 24921.03, 24940.23, 24932.77, 24952.36, 24909.75, 
    24945.95, 24900.61, 24904.53, 24916.79, 24941.55, 24947.1, 24953.06, 
    24949.38, 24931.71, 24928.85, 24916.48, 24913.06, 24903.68, 24895.98, 
    24903.01, 24910.45, 24931.72, 24951.13, 24972.75, 24978.12, 25004.18, 
    24982.91, 25018.27, 24988.13, 25040.88, 24948.08, 24987.26, 24917.35, 
    24924.69, 24938.01, 24969.27, 24952.27, 24972.18, 24928.73, 24906.71, 
    24901.06, 24890.6, 24901.3, 24900.42, 24910.76, 24907.43, 24932.43, 
    24919.01, 24957.57, 24972.02, 25014.08, 25040.78, 25068.53, 25080.9, 
    25084.7, 25086.29 ;

 HCSOI =
  24814.35, 24834.79, 24830.78, 24847.51, 24838.19, 24849.2, 24818.46, 
    24835.61, 24824.62, 24816.17, 24880.72, 24848.26, 24915.51, 24894, 
    24948.5, 24912.13, 24955.97, 24947.43, 24973.35, 24965.85, 24999.81, 
    24976.83, 25017.9, 24994.28, 24997.93, 24976.08, 24854.72, 24876.64, 
    24853.44, 24856.54, 24855.14, 24838.38, 24830.05, 24812.81, 24815.91, 
    24828.59, 24857.93, 24847.87, 24873.38, 24872.8, 24901.87, 24888.66, 
    24938.56, 24924.27, 24966.16, 24955.46, 24965.66, 24962.55, 24965.7, 
    24950.04, 24956.72, 24943.06, 24891.12, 24906.2, 24861.87, 24836.01, 
    24819.21, 24807.45, 24809.1, 24812.26, 24828.66, 24844.33, 24856.44, 
    24864.62, 24872.72, 24897.61, 24911.05, 24941.48, 24935.95, 24945.34, 
    24954.4, 24969.8, 24967.25, 24974.1, 24945.09, 24964.27, 24932.81, 
    24941.31, 24874.94, 24850.57, 24840.39, 24831.55, 24810.38, 24824.95, 
    24819.18, 24832.96, 24841.82, 24837.43, 24864.85, 24854.1, 24911.85, 
    24886.58, 24953.34, 24937.08, 24957.27, 24946.92, 24964.73, 24948.69, 
    24976.66, 24982.87, 24978.62, 24995.03, 24947.8, 24965.66, 24837.31, 
    24838.02, 24841.36, 24826.77, 24825.89, 24812.72, 24824.43, 24829.46, 
    24842.34, 24850.04, 24857.41, 24873.78, 24892.33, 24918.88, 24938.12, 
    24951.22, 24943.17, 24950.27, 24942.34, 24938.64, 24980.54, 24956.78, 
    24992.65, 24990.63, 24974.26, 24990.86, 24838.52, 24834.41, 24820.28, 
    24831.32, 24811.3, 24822.46, 24828.93, 24854.32, 24859.99, 24865.27, 
    24875.74, 24889.33, 24913.64, 24935.06, 24954.93, 24953.46, 24953.97, 
    24958.46, 24947.38, 24960.29, 24962.48, 24956.78, 24990.36, 24980.64, 
    24990.59, 24984.25, 24835.75, 24842.68, 24838.93, 24846, 24841.01, 
    24863.37, 24870.15, 24902.44, 24889.06, 24910.45, 24891.21, 24894.59, 
    24911.16, 24892.24, 24933.88, 24905.52, 24958.64, 24929.86, 24960.47, 
    24954.84, 24964.18, 24972.63, 24983.36, 25003.5, 24998.8, 25015.88, 
    24853.11, 24862.27, 24861.46, 24871.1, 24878.28, 24894, 24919.79, 
    24910.01, 24927.91, 24931.51, 24904.34, 24921.04, 24868.44, 24876.74, 
    24871.79, 24853.83, 24912.25, 24881.87, 24938.45, 24921.69, 24971.42, 
    24946.38, 24996.22, 25018.36, 25039.64, 25064.98, 24867.3, 24861.04, 
    24872.25, 24887.94, 24902.72, 24922.71, 24924.74, 24928.48, 24938.24, 
    24946.53, 24929.67, 24948.61, 24878.68, 24914.94, 24858.68, 24875.31, 
    24887.01, 24881.86, 24908.9, 24915.38, 24941.84, 24928.12, 25012.85, 
    24974.42, 25084.49, 25052.82, 24858.86, 24867.28, 24897, 24882.74, 
    24924.04, 24934.32, 24942.76, 24953.65, 24954.83, 24961.35, 24950.69, 
    24960.93, 24922.75, 24939.63, 24893.56, 24904.64, 24899.53, 24893.95, 
    24911.28, 24929.94, 24930.33, 24936.35, 24953.49, 24924.2, 25017.93, 
    24958.97, 24876.49, 24892.99, 24895.37, 24888.93, 24933.28, 24917.11, 
    24961.19, 24949.1, 24969, 24959.05, 24957.6, 24945.01, 24937.24, 
    24917.85, 24902.14, 24889.86, 24892.7, 24906.24, 24931.08, 24954.94, 
    24949.66, 24967.47, 24921.03, 24940.23, 24932.77, 24952.36, 24909.75, 
    24945.95, 24900.61, 24904.53, 24916.79, 24941.55, 24947.1, 24953.06, 
    24949.38, 24931.71, 24928.85, 24916.48, 24913.06, 24903.68, 24895.98, 
    24903.01, 24910.45, 24931.72, 24951.13, 24972.75, 24978.12, 25004.18, 
    24982.91, 25018.27, 24988.13, 25040.88, 24948.08, 24987.26, 24917.35, 
    24924.69, 24938.01, 24969.27, 24952.27, 24972.18, 24928.73, 24906.71, 
    24901.06, 24890.6, 24901.3, 24900.42, 24910.76, 24907.43, 24932.43, 
    24919.01, 24957.57, 24972.02, 25014.08, 25040.78, 25068.53, 25080.9, 
    25084.7, 25086.29 ;

 HEAT_FROM_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HR =
  6.358388e-08, 6.386347e-08, 6.380911e-08, 6.403462e-08, 6.390952e-08, 
    6.405718e-08, 6.364056e-08, 6.387457e-08, 6.372518e-08, 6.360905e-08, 
    6.447225e-08, 6.404468e-08, 6.491634e-08, 6.464366e-08, 6.532863e-08, 
    6.487392e-08, 6.542031e-08, 6.53155e-08, 6.563094e-08, 6.554057e-08, 
    6.594404e-08, 6.567264e-08, 6.615318e-08, 6.587923e-08, 6.592209e-08, 
    6.566369e-08, 6.413072e-08, 6.441902e-08, 6.411364e-08, 6.415475e-08, 
    6.41363e-08, 6.391211e-08, 6.379913e-08, 6.356251e-08, 6.360547e-08, 
    6.377926e-08, 6.417324e-08, 6.403949e-08, 6.437654e-08, 6.436893e-08, 
    6.474416e-08, 6.457498e-08, 6.520563e-08, 6.502638e-08, 6.554434e-08, 
    6.541408e-08, 6.553822e-08, 6.550058e-08, 6.553871e-08, 6.534768e-08, 
    6.542952e-08, 6.526142e-08, 6.460666e-08, 6.47991e-08, 6.422516e-08, 
    6.388007e-08, 6.365083e-08, 6.348817e-08, 6.351116e-08, 6.3555e-08, 
    6.378028e-08, 6.399208e-08, 6.415348e-08, 6.426145e-08, 6.436783e-08, 
    6.468986e-08, 6.486028e-08, 6.524188e-08, 6.5173e-08, 6.528968e-08, 
    6.540112e-08, 6.558825e-08, 6.555744e-08, 6.563989e-08, 6.528659e-08, 
    6.55214e-08, 6.513378e-08, 6.52398e-08, 6.439678e-08, 6.407557e-08, 
    6.393907e-08, 6.381956e-08, 6.352884e-08, 6.372961e-08, 6.365047e-08, 
    6.383875e-08, 6.395839e-08, 6.389921e-08, 6.426441e-08, 6.412242e-08, 
    6.487038e-08, 6.454822e-08, 6.538812e-08, 6.518714e-08, 6.54363e-08, 
    6.530916e-08, 6.5527e-08, 6.533094e-08, 6.567057e-08, 6.574452e-08, 
    6.569399e-08, 6.588811e-08, 6.532007e-08, 6.553822e-08, 6.389756e-08, 
    6.390721e-08, 6.395216e-08, 6.375454e-08, 6.374245e-08, 6.356133e-08, 
    6.372249e-08, 6.379111e-08, 6.396532e-08, 6.406837e-08, 6.416632e-08, 
    6.438169e-08, 6.462222e-08, 6.495855e-08, 6.520017e-08, 6.536213e-08, 
    6.526282e-08, 6.53505e-08, 6.525248e-08, 6.520654e-08, 6.571682e-08, 
    6.543029e-08, 6.586019e-08, 6.58364e-08, 6.564185e-08, 6.583908e-08, 
    6.391399e-08, 6.385844e-08, 6.366564e-08, 6.381653e-08, 6.354161e-08, 
    6.36955e-08, 6.378399e-08, 6.41254e-08, 6.420041e-08, 6.426996e-08, 
    6.440733e-08, 6.458363e-08, 6.489289e-08, 6.516198e-08, 6.54076e-08, 
    6.538961e-08, 6.539594e-08, 6.545082e-08, 6.531489e-08, 6.547314e-08, 
    6.54997e-08, 6.543026e-08, 6.583321e-08, 6.571809e-08, 6.58359e-08, 
    6.576094e-08, 6.38765e-08, 6.396994e-08, 6.391945e-08, 6.40144e-08, 
    6.394751e-08, 6.424496e-08, 6.433414e-08, 6.475143e-08, 6.458016e-08, 
    6.485271e-08, 6.460785e-08, 6.465124e-08, 6.486162e-08, 6.462108e-08, 
    6.514714e-08, 6.47905e-08, 6.545295e-08, 6.509682e-08, 6.547527e-08, 
    6.540655e-08, 6.552033e-08, 6.562224e-08, 6.575045e-08, 6.598701e-08, 
    6.593223e-08, 6.613006e-08, 6.410925e-08, 6.423046e-08, 6.421978e-08, 
    6.434662e-08, 6.444042e-08, 6.464373e-08, 6.496981e-08, 6.484719e-08, 
    6.507229e-08, 6.511748e-08, 6.477549e-08, 6.498548e-08, 6.431157e-08, 
    6.442045e-08, 6.435562e-08, 6.411882e-08, 6.487545e-08, 6.448715e-08, 
    6.520416e-08, 6.499381e-08, 6.560771e-08, 6.530242e-08, 6.590207e-08, 
    6.615844e-08, 6.639969e-08, 6.668164e-08, 6.42966e-08, 6.421424e-08, 
    6.43617e-08, 6.456572e-08, 6.4755e-08, 6.500665e-08, 6.503239e-08, 
    6.507953e-08, 6.520164e-08, 6.530431e-08, 6.509445e-08, 6.533005e-08, 
    6.444572e-08, 6.490915e-08, 6.418311e-08, 6.440175e-08, 6.455369e-08, 
    6.448703e-08, 6.483317e-08, 6.491475e-08, 6.524627e-08, 6.507489e-08, 
    6.609517e-08, 6.564377e-08, 6.689631e-08, 6.654629e-08, 6.418547e-08, 
    6.429631e-08, 6.468208e-08, 6.449854e-08, 6.502344e-08, 6.515264e-08, 
    6.525767e-08, 6.539194e-08, 6.540643e-08, 6.548598e-08, 6.535562e-08, 
    6.548083e-08, 6.500718e-08, 6.521884e-08, 6.463799e-08, 6.477936e-08, 
    6.471433e-08, 6.464298e-08, 6.486317e-08, 6.509775e-08, 6.510275e-08, 
    6.517797e-08, 6.538995e-08, 6.502557e-08, 6.615345e-08, 6.545692e-08, 
    6.441718e-08, 6.463069e-08, 6.466117e-08, 6.457847e-08, 6.513969e-08, 
    6.493634e-08, 6.548404e-08, 6.533602e-08, 6.557855e-08, 6.545803e-08, 
    6.54403e-08, 6.528551e-08, 6.518914e-08, 6.494567e-08, 6.474756e-08, 
    6.459047e-08, 6.4627e-08, 6.479956e-08, 6.51121e-08, 6.540775e-08, 
    6.534299e-08, 6.556012e-08, 6.498538e-08, 6.522639e-08, 6.513324e-08, 
    6.537611e-08, 6.484393e-08, 6.529714e-08, 6.472809e-08, 6.477798e-08, 
    6.493231e-08, 6.524274e-08, 6.53114e-08, 6.538474e-08, 6.533948e-08, 
    6.512003e-08, 6.508407e-08, 6.492856e-08, 6.488562e-08, 6.476711e-08, 
    6.466901e-08, 6.475865e-08, 6.485278e-08, 6.512012e-08, 6.536104e-08, 
    6.562369e-08, 6.568797e-08, 6.599488e-08, 6.574506e-08, 6.615733e-08, 
    6.580684e-08, 6.641355e-08, 6.532339e-08, 6.579651e-08, 6.493933e-08, 
    6.503167e-08, 6.519871e-08, 6.558179e-08, 6.537497e-08, 6.561685e-08, 
    6.508266e-08, 6.480552e-08, 6.47338e-08, 6.460002e-08, 6.473686e-08, 
    6.472573e-08, 6.485668e-08, 6.48146e-08, 6.512899e-08, 6.496011e-08, 
    6.543986e-08, 6.561493e-08, 6.610933e-08, 6.641241e-08, 6.672092e-08, 
    6.685712e-08, 6.689857e-08, 6.69159e-08 ;

 HR_vr =
  2.668957e-07, 2.676048e-07, 2.67467e-07, 2.680385e-07, 2.677215e-07, 
    2.680956e-07, 2.670395e-07, 2.676329e-07, 2.672542e-07, 2.669595e-07, 
    2.691461e-07, 2.68064e-07, 2.702677e-07, 2.695792e-07, 2.713072e-07, 
    2.701607e-07, 2.715381e-07, 2.712741e-07, 2.720682e-07, 2.718408e-07, 
    2.728555e-07, 2.721731e-07, 2.733806e-07, 2.726925e-07, 2.728003e-07, 
    2.721506e-07, 2.682818e-07, 2.690115e-07, 2.682386e-07, 2.683427e-07, 
    2.68296e-07, 2.677281e-07, 2.674417e-07, 2.668415e-07, 2.669505e-07, 
    2.673913e-07, 2.683895e-07, 2.680508e-07, 2.689039e-07, 2.688846e-07, 
    2.69833e-07, 2.694056e-07, 2.709972e-07, 2.705453e-07, 2.718503e-07, 
    2.715224e-07, 2.718349e-07, 2.717402e-07, 2.718362e-07, 2.713552e-07, 
    2.715613e-07, 2.711378e-07, 2.694857e-07, 2.699718e-07, 2.685209e-07, 
    2.676469e-07, 2.670656e-07, 2.666527e-07, 2.667111e-07, 2.668224e-07, 
    2.673939e-07, 2.679307e-07, 2.683394e-07, 2.686127e-07, 2.688819e-07, 
    2.69696e-07, 2.701263e-07, 2.710886e-07, 2.70915e-07, 2.71209e-07, 
    2.714898e-07, 2.719608e-07, 2.718833e-07, 2.720907e-07, 2.712013e-07, 
    2.717926e-07, 2.708161e-07, 2.710833e-07, 2.689552e-07, 2.681422e-07, 
    2.677964e-07, 2.674935e-07, 2.66756e-07, 2.672654e-07, 2.670646e-07, 
    2.675421e-07, 2.678453e-07, 2.676954e-07, 2.686202e-07, 2.682608e-07, 
    2.701518e-07, 2.69338e-07, 2.71457e-07, 2.709506e-07, 2.715783e-07, 
    2.712581e-07, 2.718067e-07, 2.71313e-07, 2.721679e-07, 2.723539e-07, 
    2.722268e-07, 2.727149e-07, 2.712856e-07, 2.718349e-07, 2.676912e-07, 
    2.677156e-07, 2.678296e-07, 2.673286e-07, 2.67298e-07, 2.668385e-07, 
    2.672473e-07, 2.674214e-07, 2.678629e-07, 2.681239e-07, 2.68372e-07, 
    2.689169e-07, 2.69525e-07, 2.703742e-07, 2.709835e-07, 2.713915e-07, 
    2.711413e-07, 2.713622e-07, 2.711153e-07, 2.709995e-07, 2.722843e-07, 
    2.715632e-07, 2.726447e-07, 2.725849e-07, 2.720957e-07, 2.725916e-07, 
    2.677328e-07, 2.67592e-07, 2.671031e-07, 2.674858e-07, 2.667884e-07, 
    2.671789e-07, 2.674033e-07, 2.682684e-07, 2.684582e-07, 2.686343e-07, 
    2.689818e-07, 2.694275e-07, 2.702085e-07, 2.708872e-07, 2.715061e-07, 
    2.714607e-07, 2.714767e-07, 2.716149e-07, 2.712726e-07, 2.716711e-07, 
    2.717379e-07, 2.715631e-07, 2.725769e-07, 2.722875e-07, 2.725836e-07, 
    2.723952e-07, 2.676378e-07, 2.678746e-07, 2.677467e-07, 2.679872e-07, 
    2.678178e-07, 2.68571e-07, 2.687967e-07, 2.698514e-07, 2.694187e-07, 
    2.701071e-07, 2.694887e-07, 2.695983e-07, 2.701297e-07, 2.695221e-07, 
    2.708499e-07, 2.699501e-07, 2.716203e-07, 2.707231e-07, 2.716765e-07, 
    2.715034e-07, 2.717899e-07, 2.720463e-07, 2.723688e-07, 2.729634e-07, 
    2.728257e-07, 2.733226e-07, 2.682274e-07, 2.685343e-07, 2.685073e-07, 
    2.688282e-07, 2.690655e-07, 2.695793e-07, 2.704026e-07, 2.700932e-07, 
    2.706611e-07, 2.70775e-07, 2.699121e-07, 2.704422e-07, 2.687396e-07, 
    2.69015e-07, 2.68851e-07, 2.682517e-07, 2.701645e-07, 2.691837e-07, 
    2.709936e-07, 2.704632e-07, 2.720098e-07, 2.712412e-07, 2.7275e-07, 
    2.733939e-07, 2.73999e-07, 2.747055e-07, 2.687017e-07, 2.684932e-07, 
    2.688664e-07, 2.693823e-07, 2.698604e-07, 2.704955e-07, 2.705605e-07, 
    2.706794e-07, 2.709872e-07, 2.712459e-07, 2.70717e-07, 2.713107e-07, 
    2.69079e-07, 2.702496e-07, 2.684145e-07, 2.689677e-07, 2.693519e-07, 
    2.691833e-07, 2.700578e-07, 2.702637e-07, 2.710997e-07, 2.706677e-07, 
    2.73235e-07, 2.721006e-07, 2.752428e-07, 2.743665e-07, 2.684204e-07, 
    2.687009e-07, 2.696763e-07, 2.692124e-07, 2.705379e-07, 2.708637e-07, 
    2.711284e-07, 2.714667e-07, 2.715031e-07, 2.717034e-07, 2.713752e-07, 
    2.716905e-07, 2.704969e-07, 2.710305e-07, 2.695648e-07, 2.699219e-07, 
    2.697577e-07, 2.695775e-07, 2.701335e-07, 2.707254e-07, 2.707379e-07, 
    2.709275e-07, 2.714618e-07, 2.705433e-07, 2.733814e-07, 2.716304e-07, 
    2.690067e-07, 2.695465e-07, 2.696234e-07, 2.694144e-07, 2.70831e-07, 
    2.703182e-07, 2.716986e-07, 2.713258e-07, 2.719364e-07, 2.716331e-07, 
    2.715884e-07, 2.711985e-07, 2.709557e-07, 2.703417e-07, 2.698416e-07, 
    2.694447e-07, 2.695371e-07, 2.69973e-07, 2.707615e-07, 2.715065e-07, 
    2.713433e-07, 2.7189e-07, 2.704419e-07, 2.710496e-07, 2.708148e-07, 
    2.714268e-07, 2.700849e-07, 2.71228e-07, 2.697924e-07, 2.699184e-07, 
    2.70308e-07, 2.710908e-07, 2.712638e-07, 2.714485e-07, 2.713345e-07, 
    2.707815e-07, 2.706908e-07, 2.702985e-07, 2.701902e-07, 2.69891e-07, 
    2.696432e-07, 2.698696e-07, 2.701073e-07, 2.707817e-07, 2.713888e-07, 
    2.7205e-07, 2.722117e-07, 2.729832e-07, 2.723553e-07, 2.733912e-07, 
    2.725107e-07, 2.740339e-07, 2.71294e-07, 2.724847e-07, 2.703257e-07, 
    2.705587e-07, 2.709798e-07, 2.719446e-07, 2.714239e-07, 2.720328e-07, 
    2.706873e-07, 2.69988e-07, 2.698069e-07, 2.694689e-07, 2.698146e-07, 
    2.697865e-07, 2.701171e-07, 2.700109e-07, 2.70804e-07, 2.703782e-07, 
    2.715873e-07, 2.72028e-07, 2.732705e-07, 2.74031e-07, 2.748038e-07, 
    2.751447e-07, 2.752484e-07, 2.752918e-07,
  2.415169e-07, 2.424272e-07, 2.422503e-07, 2.42984e-07, 2.425771e-07, 
    2.430574e-07, 2.417015e-07, 2.424633e-07, 2.419771e-07, 2.415989e-07, 
    2.444062e-07, 2.430167e-07, 2.458473e-07, 2.449628e-07, 2.47183e-07, 
    2.457097e-07, 2.474798e-07, 2.471405e-07, 2.481612e-07, 2.478689e-07, 
    2.491731e-07, 2.482961e-07, 2.498484e-07, 2.489637e-07, 2.491022e-07, 
    2.482671e-07, 2.432965e-07, 2.442333e-07, 2.43241e-07, 2.433746e-07, 
    2.433147e-07, 2.425855e-07, 2.422178e-07, 2.414473e-07, 2.415872e-07, 
    2.421531e-07, 2.434347e-07, 2.429999e-07, 2.440954e-07, 2.440707e-07, 
    2.452889e-07, 2.447399e-07, 2.467848e-07, 2.462041e-07, 2.478811e-07, 
    2.474597e-07, 2.478614e-07, 2.477396e-07, 2.478629e-07, 2.472447e-07, 
    2.475096e-07, 2.469654e-07, 2.448427e-07, 2.454671e-07, 2.436036e-07, 
    2.424811e-07, 2.417349e-07, 2.412051e-07, 2.4128e-07, 2.414228e-07, 
    2.421564e-07, 2.428457e-07, 2.433706e-07, 2.437215e-07, 2.440672e-07, 
    2.451126e-07, 2.456655e-07, 2.469021e-07, 2.466791e-07, 2.470569e-07, 
    2.474177e-07, 2.480232e-07, 2.479235e-07, 2.481902e-07, 2.47047e-07, 
    2.478069e-07, 2.46552e-07, 2.468954e-07, 2.44161e-07, 2.431172e-07, 
    2.426731e-07, 2.422843e-07, 2.413376e-07, 2.419915e-07, 2.417338e-07, 
    2.423468e-07, 2.427361e-07, 2.425436e-07, 2.437311e-07, 2.432696e-07, 
    2.456982e-07, 2.446529e-07, 2.473757e-07, 2.467249e-07, 2.475316e-07, 
    2.4712e-07, 2.47825e-07, 2.471906e-07, 2.482894e-07, 2.485284e-07, 
    2.483651e-07, 2.489925e-07, 2.471554e-07, 2.478613e-07, 2.425382e-07, 
    2.425696e-07, 2.427159e-07, 2.420726e-07, 2.420333e-07, 2.414435e-07, 
    2.419683e-07, 2.421917e-07, 2.427586e-07, 2.430938e-07, 2.434123e-07, 
    2.441122e-07, 2.448932e-07, 2.459841e-07, 2.467671e-07, 2.472915e-07, 
    2.4697e-07, 2.472539e-07, 2.469365e-07, 2.467877e-07, 2.484389e-07, 
    2.475121e-07, 2.489023e-07, 2.488254e-07, 2.481965e-07, 2.488341e-07, 
    2.425916e-07, 2.424109e-07, 2.417832e-07, 2.422745e-07, 2.413792e-07, 
    2.418804e-07, 2.421685e-07, 2.432792e-07, 2.435231e-07, 2.437492e-07, 
    2.441955e-07, 2.44768e-07, 2.457713e-07, 2.466433e-07, 2.474387e-07, 
    2.473805e-07, 2.47401e-07, 2.475786e-07, 2.471386e-07, 2.476508e-07, 
    2.477367e-07, 2.47512e-07, 2.488151e-07, 2.48443e-07, 2.488238e-07, 
    2.485815e-07, 2.424696e-07, 2.427737e-07, 2.426094e-07, 2.429183e-07, 
    2.427007e-07, 2.436679e-07, 2.439576e-07, 2.453124e-07, 2.447567e-07, 
    2.45641e-07, 2.448465e-07, 2.449874e-07, 2.456698e-07, 2.448895e-07, 
    2.465952e-07, 2.454391e-07, 2.475855e-07, 2.464322e-07, 2.476577e-07, 
    2.474353e-07, 2.478035e-07, 2.481331e-07, 2.485476e-07, 2.493119e-07, 
    2.49135e-07, 2.497738e-07, 2.432267e-07, 2.436207e-07, 2.435861e-07, 
    2.439982e-07, 2.44303e-07, 2.44963e-07, 2.460207e-07, 2.456231e-07, 
    2.463528e-07, 2.464992e-07, 2.453906e-07, 2.460714e-07, 2.438843e-07, 
    2.44238e-07, 2.440275e-07, 2.432578e-07, 2.457147e-07, 2.444546e-07, 
    2.4678e-07, 2.460985e-07, 2.480861e-07, 2.470981e-07, 2.490376e-07, 
    2.498653e-07, 2.506436e-07, 2.515522e-07, 2.438357e-07, 2.435681e-07, 
    2.440472e-07, 2.447098e-07, 2.453241e-07, 2.461401e-07, 2.462235e-07, 
    2.463763e-07, 2.467719e-07, 2.471043e-07, 2.464246e-07, 2.471877e-07, 
    2.4432e-07, 2.45824e-07, 2.434669e-07, 2.441773e-07, 2.446707e-07, 
    2.444543e-07, 2.455776e-07, 2.458422e-07, 2.469164e-07, 2.463613e-07, 
    2.49661e-07, 2.482027e-07, 2.522434e-07, 2.511161e-07, 2.434745e-07, 
    2.438348e-07, 2.450874e-07, 2.444917e-07, 2.461945e-07, 2.466131e-07, 
    2.469533e-07, 2.47388e-07, 2.474349e-07, 2.476923e-07, 2.472705e-07, 
    2.476757e-07, 2.461418e-07, 2.468276e-07, 2.449444e-07, 2.454031e-07, 
    2.451921e-07, 2.449606e-07, 2.456749e-07, 2.464353e-07, 2.464515e-07, 
    2.466952e-07, 2.473814e-07, 2.462014e-07, 2.498491e-07, 2.475981e-07, 
    2.442275e-07, 2.449206e-07, 2.450196e-07, 2.447512e-07, 2.465712e-07, 
    2.459122e-07, 2.476861e-07, 2.47207e-07, 2.479918e-07, 2.476019e-07, 
    2.475445e-07, 2.470435e-07, 2.467314e-07, 2.459424e-07, 2.452999e-07, 
    2.447902e-07, 2.449087e-07, 2.454686e-07, 2.464818e-07, 2.474391e-07, 
    2.472295e-07, 2.479322e-07, 2.460712e-07, 2.46852e-07, 2.465502e-07, 
    2.473368e-07, 2.456125e-07, 2.470809e-07, 2.452368e-07, 2.453986e-07, 
    2.458991e-07, 2.469049e-07, 2.471273e-07, 2.473647e-07, 2.472182e-07, 
    2.465074e-07, 2.46391e-07, 2.458869e-07, 2.457477e-07, 2.453634e-07, 
    2.450451e-07, 2.453359e-07, 2.456412e-07, 2.465077e-07, 2.472879e-07, 
    2.481378e-07, 2.483456e-07, 2.493372e-07, 2.485301e-07, 2.498616e-07, 
    2.487296e-07, 2.506881e-07, 2.47166e-07, 2.486964e-07, 2.459219e-07, 
    2.462212e-07, 2.467623e-07, 2.480022e-07, 2.473331e-07, 2.481156e-07, 
    2.463864e-07, 2.454879e-07, 2.452553e-07, 2.448211e-07, 2.452652e-07, 
    2.452291e-07, 2.456539e-07, 2.455174e-07, 2.465365e-07, 2.459893e-07, 
    2.475431e-07, 2.481094e-07, 2.497068e-07, 2.506846e-07, 2.516788e-07, 
    2.521173e-07, 2.522507e-07, 2.523065e-07,
  2.260081e-07, 2.270054e-07, 2.268116e-07, 2.276156e-07, 2.271697e-07, 
    2.276961e-07, 2.262103e-07, 2.27045e-07, 2.265122e-07, 2.260979e-07, 
    2.291747e-07, 2.276515e-07, 2.307554e-07, 2.297851e-07, 2.322212e-07, 
    2.306044e-07, 2.32547e-07, 2.321746e-07, 2.332951e-07, 2.329742e-07, 
    2.344063e-07, 2.334432e-07, 2.351482e-07, 2.341764e-07, 2.343285e-07, 
    2.334114e-07, 2.279582e-07, 2.289851e-07, 2.278973e-07, 2.280438e-07, 
    2.279781e-07, 2.271789e-07, 2.26776e-07, 2.259318e-07, 2.260851e-07, 
    2.267051e-07, 2.281097e-07, 2.276331e-07, 2.28834e-07, 2.288069e-07, 
    2.301428e-07, 2.295406e-07, 2.317841e-07, 2.311468e-07, 2.329876e-07, 
    2.325249e-07, 2.329658e-07, 2.328322e-07, 2.329676e-07, 2.322889e-07, 
    2.325797e-07, 2.319824e-07, 2.296534e-07, 2.303383e-07, 2.282947e-07, 
    2.270645e-07, 2.26247e-07, 2.256665e-07, 2.257486e-07, 2.25905e-07, 
    2.267087e-07, 2.27464e-07, 2.280393e-07, 2.284241e-07, 2.28803e-07, 
    2.299494e-07, 2.305559e-07, 2.319129e-07, 2.316681e-07, 2.320828e-07, 
    2.324788e-07, 2.331435e-07, 2.330341e-07, 2.333269e-07, 2.320719e-07, 
    2.32906e-07, 2.315287e-07, 2.319055e-07, 2.289059e-07, 2.277617e-07, 
    2.272749e-07, 2.268489e-07, 2.258117e-07, 2.26528e-07, 2.262457e-07, 
    2.269173e-07, 2.273439e-07, 2.271329e-07, 2.284346e-07, 2.279287e-07, 
    2.305919e-07, 2.294453e-07, 2.324326e-07, 2.317184e-07, 2.326038e-07, 
    2.321521e-07, 2.32926e-07, 2.322295e-07, 2.334358e-07, 2.336983e-07, 
    2.335189e-07, 2.34208e-07, 2.321909e-07, 2.329658e-07, 2.27127e-07, 
    2.271614e-07, 2.273217e-07, 2.266169e-07, 2.265738e-07, 2.259276e-07, 
    2.265026e-07, 2.267474e-07, 2.273686e-07, 2.27736e-07, 2.280851e-07, 
    2.288524e-07, 2.297088e-07, 2.309055e-07, 2.317647e-07, 2.323403e-07, 
    2.319874e-07, 2.32299e-07, 2.319506e-07, 2.317874e-07, 2.336e-07, 
    2.325824e-07, 2.341089e-07, 2.340245e-07, 2.333338e-07, 2.34034e-07, 
    2.271856e-07, 2.269876e-07, 2.262998e-07, 2.268381e-07, 2.258572e-07, 
    2.264063e-07, 2.26722e-07, 2.279392e-07, 2.282066e-07, 2.284544e-07, 
    2.289437e-07, 2.295715e-07, 2.30672e-07, 2.316289e-07, 2.325019e-07, 
    2.324379e-07, 2.324605e-07, 2.326554e-07, 2.321724e-07, 2.327346e-07, 
    2.32829e-07, 2.325823e-07, 2.340132e-07, 2.336045e-07, 2.340227e-07, 
    2.337566e-07, 2.27052e-07, 2.273851e-07, 2.272051e-07, 2.275436e-07, 
    2.273051e-07, 2.283653e-07, 2.286829e-07, 2.301686e-07, 2.295591e-07, 
    2.305291e-07, 2.296577e-07, 2.298121e-07, 2.305606e-07, 2.297048e-07, 
    2.315761e-07, 2.303076e-07, 2.32663e-07, 2.313972e-07, 2.327422e-07, 
    2.324981e-07, 2.329023e-07, 2.332642e-07, 2.337194e-07, 2.345588e-07, 
    2.343645e-07, 2.350662e-07, 2.278817e-07, 2.283136e-07, 2.282756e-07, 
    2.287274e-07, 2.290615e-07, 2.297854e-07, 2.309456e-07, 2.305094e-07, 
    2.313101e-07, 2.314708e-07, 2.302543e-07, 2.310013e-07, 2.286026e-07, 
    2.289904e-07, 2.287595e-07, 2.279158e-07, 2.306099e-07, 2.292279e-07, 
    2.317789e-07, 2.31031e-07, 2.332126e-07, 2.32128e-07, 2.342575e-07, 
    2.351668e-07, 2.360221e-07, 2.370208e-07, 2.285493e-07, 2.282559e-07, 
    2.287812e-07, 2.295076e-07, 2.301814e-07, 2.310766e-07, 2.311682e-07, 
    2.313358e-07, 2.317699e-07, 2.321348e-07, 2.313888e-07, 2.322263e-07, 
    2.290803e-07, 2.307298e-07, 2.281449e-07, 2.289238e-07, 2.294648e-07, 
    2.292275e-07, 2.304596e-07, 2.307498e-07, 2.319285e-07, 2.313193e-07, 
    2.349424e-07, 2.333406e-07, 2.377808e-07, 2.365414e-07, 2.281533e-07, 
    2.285483e-07, 2.299219e-07, 2.292685e-07, 2.311364e-07, 2.315957e-07, 
    2.319691e-07, 2.324462e-07, 2.324977e-07, 2.327803e-07, 2.323172e-07, 
    2.32762e-07, 2.310785e-07, 2.318311e-07, 2.29765e-07, 2.302681e-07, 
    2.300367e-07, 2.297828e-07, 2.305663e-07, 2.314005e-07, 2.314184e-07, 
    2.316858e-07, 2.324389e-07, 2.311439e-07, 2.351489e-07, 2.326768e-07, 
    2.289788e-07, 2.297389e-07, 2.298475e-07, 2.295531e-07, 2.315497e-07, 
    2.308266e-07, 2.327734e-07, 2.322475e-07, 2.331091e-07, 2.32681e-07, 
    2.32618e-07, 2.32068e-07, 2.317255e-07, 2.308597e-07, 2.301549e-07, 
    2.295958e-07, 2.297258e-07, 2.3034e-07, 2.314516e-07, 2.325023e-07, 
    2.322722e-07, 2.330436e-07, 2.31001e-07, 2.318579e-07, 2.315267e-07, 
    2.3239e-07, 2.304978e-07, 2.321092e-07, 2.300857e-07, 2.302632e-07, 
    2.308122e-07, 2.319159e-07, 2.3216e-07, 2.324206e-07, 2.322598e-07, 
    2.314798e-07, 2.313519e-07, 2.307989e-07, 2.306461e-07, 2.302245e-07, 
    2.298754e-07, 2.301944e-07, 2.305293e-07, 2.314801e-07, 2.323364e-07, 
    2.332693e-07, 2.334976e-07, 2.345866e-07, 2.337001e-07, 2.351627e-07, 
    2.339193e-07, 2.36071e-07, 2.322025e-07, 2.338828e-07, 2.308372e-07, 
    2.311656e-07, 2.317594e-07, 2.331205e-07, 2.323859e-07, 2.33245e-07, 
    2.313469e-07, 2.303611e-07, 2.30106e-07, 2.296298e-07, 2.301169e-07, 
    2.300773e-07, 2.305432e-07, 2.303935e-07, 2.315116e-07, 2.309111e-07, 
    2.326164e-07, 2.332382e-07, 2.349927e-07, 2.360671e-07, 2.3716e-07, 
    2.376421e-07, 2.377888e-07, 2.378502e-07,
  2.166788e-07, 2.177054e-07, 2.175058e-07, 2.183338e-07, 2.178745e-07, 
    2.184166e-07, 2.168869e-07, 2.177461e-07, 2.171977e-07, 2.167712e-07, 
    2.199401e-07, 2.183707e-07, 2.215698e-07, 2.205693e-07, 2.230824e-07, 
    2.214141e-07, 2.234187e-07, 2.230342e-07, 2.241912e-07, 2.238598e-07, 
    2.253393e-07, 2.243441e-07, 2.261061e-07, 2.251017e-07, 2.252588e-07, 
    2.243113e-07, 2.186866e-07, 2.197448e-07, 2.186239e-07, 2.187748e-07, 
    2.18707e-07, 2.17884e-07, 2.174692e-07, 2.166003e-07, 2.167581e-07, 
    2.173962e-07, 2.188426e-07, 2.183517e-07, 2.195889e-07, 2.195609e-07, 
    2.20938e-07, 2.203172e-07, 2.226312e-07, 2.219736e-07, 2.238736e-07, 
    2.233958e-07, 2.238512e-07, 2.237131e-07, 2.23853e-07, 2.231522e-07, 
    2.234525e-07, 2.228359e-07, 2.204335e-07, 2.211396e-07, 2.190332e-07, 
    2.177663e-07, 2.169246e-07, 2.163273e-07, 2.164117e-07, 2.165727e-07, 
    2.173999e-07, 2.181776e-07, 2.187701e-07, 2.191665e-07, 2.195569e-07, 
    2.207388e-07, 2.213641e-07, 2.227642e-07, 2.225115e-07, 2.229395e-07, 
    2.233483e-07, 2.240346e-07, 2.239217e-07, 2.24224e-07, 2.229282e-07, 
    2.237894e-07, 2.223676e-07, 2.227565e-07, 2.196631e-07, 2.184841e-07, 
    2.179829e-07, 2.175442e-07, 2.164767e-07, 2.172139e-07, 2.169233e-07, 
    2.176146e-07, 2.180539e-07, 2.178366e-07, 2.191773e-07, 2.186561e-07, 
    2.214012e-07, 2.20219e-07, 2.233006e-07, 2.225634e-07, 2.234773e-07, 
    2.23011e-07, 2.2381e-07, 2.230909e-07, 2.243365e-07, 2.246077e-07, 
    2.244224e-07, 2.251343e-07, 2.23051e-07, 2.238512e-07, 2.178306e-07, 
    2.17866e-07, 2.180311e-07, 2.173054e-07, 2.17261e-07, 2.16596e-07, 
    2.171878e-07, 2.174397e-07, 2.180794e-07, 2.184577e-07, 2.188172e-07, 
    2.196078e-07, 2.204906e-07, 2.217247e-07, 2.226111e-07, 2.232053e-07, 
    2.22841e-07, 2.231626e-07, 2.228031e-07, 2.226345e-07, 2.245061e-07, 
    2.234553e-07, 2.250319e-07, 2.249446e-07, 2.242312e-07, 2.249545e-07, 
    2.178909e-07, 2.17687e-07, 2.16979e-07, 2.175331e-07, 2.165236e-07, 
    2.170887e-07, 2.174136e-07, 2.18667e-07, 2.189424e-07, 2.191977e-07, 
    2.197019e-07, 2.20349e-07, 2.214838e-07, 2.22471e-07, 2.233721e-07, 
    2.233061e-07, 2.233293e-07, 2.235306e-07, 2.23032e-07, 2.236124e-07, 
    2.237098e-07, 2.234551e-07, 2.24933e-07, 2.245108e-07, 2.249428e-07, 
    2.246679e-07, 2.177533e-07, 2.180963e-07, 2.17911e-07, 2.182595e-07, 
    2.18014e-07, 2.191059e-07, 2.194332e-07, 2.209647e-07, 2.203362e-07, 
    2.213364e-07, 2.204378e-07, 2.205971e-07, 2.21369e-07, 2.204864e-07, 
    2.224166e-07, 2.211081e-07, 2.235384e-07, 2.22232e-07, 2.236203e-07, 
    2.233682e-07, 2.237855e-07, 2.241593e-07, 2.246294e-07, 2.254969e-07, 
    2.25296e-07, 2.260213e-07, 2.186078e-07, 2.190527e-07, 2.190135e-07, 
    2.194791e-07, 2.198234e-07, 2.205695e-07, 2.21766e-07, 2.213161e-07, 
    2.22142e-07, 2.223078e-07, 2.21053e-07, 2.218235e-07, 2.193504e-07, 
    2.197501e-07, 2.195121e-07, 2.186429e-07, 2.214198e-07, 2.199948e-07, 
    2.226258e-07, 2.218541e-07, 2.24106e-07, 2.229862e-07, 2.251854e-07, 
    2.261254e-07, 2.270097e-07, 2.280431e-07, 2.192955e-07, 2.189932e-07, 
    2.195344e-07, 2.202832e-07, 2.209778e-07, 2.219012e-07, 2.219956e-07, 
    2.221686e-07, 2.226166e-07, 2.229932e-07, 2.222233e-07, 2.230876e-07, 
    2.198428e-07, 2.215435e-07, 2.188789e-07, 2.196814e-07, 2.202391e-07, 
    2.199944e-07, 2.212647e-07, 2.21564e-07, 2.227803e-07, 2.221516e-07, 
    2.258934e-07, 2.242382e-07, 2.288297e-07, 2.27547e-07, 2.188875e-07, 
    2.192944e-07, 2.207103e-07, 2.200367e-07, 2.219628e-07, 2.224368e-07, 
    2.228221e-07, 2.233146e-07, 2.233678e-07, 2.236596e-07, 2.231814e-07, 
    2.236407e-07, 2.219031e-07, 2.226797e-07, 2.205484e-07, 2.210672e-07, 
    2.208286e-07, 2.205668e-07, 2.213747e-07, 2.222354e-07, 2.222538e-07, 
    2.225297e-07, 2.233073e-07, 2.219706e-07, 2.26107e-07, 2.235529e-07, 
    2.197381e-07, 2.205216e-07, 2.206335e-07, 2.2033e-07, 2.223893e-07, 
    2.216432e-07, 2.236524e-07, 2.231095e-07, 2.239991e-07, 2.23557e-07, 
    2.23492e-07, 2.229242e-07, 2.225707e-07, 2.216775e-07, 2.209505e-07, 
    2.20374e-07, 2.205081e-07, 2.211413e-07, 2.222881e-07, 2.233726e-07, 
    2.23135e-07, 2.239315e-07, 2.218232e-07, 2.227073e-07, 2.223656e-07, 
    2.232566e-07, 2.213041e-07, 2.229668e-07, 2.208791e-07, 2.210622e-07, 
    2.216284e-07, 2.227673e-07, 2.230192e-07, 2.232882e-07, 2.231222e-07, 
    2.223171e-07, 2.221852e-07, 2.216147e-07, 2.214571e-07, 2.210223e-07, 
    2.206623e-07, 2.209912e-07, 2.213366e-07, 2.223175e-07, 2.232012e-07, 
    2.241646e-07, 2.244003e-07, 2.255257e-07, 2.246096e-07, 2.261212e-07, 
    2.248362e-07, 2.270605e-07, 2.230631e-07, 2.247983e-07, 2.216542e-07, 
    2.21993e-07, 2.226058e-07, 2.240109e-07, 2.232524e-07, 2.241395e-07, 
    2.221801e-07, 2.211632e-07, 2.209e-07, 2.204091e-07, 2.209113e-07, 
    2.208704e-07, 2.213509e-07, 2.211965e-07, 2.2235e-07, 2.217305e-07, 
    2.234904e-07, 2.241325e-07, 2.259453e-07, 2.270564e-07, 2.28187e-07, 
    2.286861e-07, 2.28838e-07, 2.289015e-07,
  2.081592e-07, 2.091281e-07, 2.089397e-07, 2.097215e-07, 2.092877e-07, 
    2.097998e-07, 2.083556e-07, 2.091666e-07, 2.086488e-07, 2.082464e-07, 
    2.112401e-07, 2.097564e-07, 2.127826e-07, 2.118352e-07, 2.142163e-07, 
    2.126352e-07, 2.145353e-07, 2.141706e-07, 2.152684e-07, 2.149538e-07, 
    2.163592e-07, 2.154136e-07, 2.170881e-07, 2.161333e-07, 2.162826e-07, 
    2.153825e-07, 2.100548e-07, 2.110553e-07, 2.099955e-07, 2.101382e-07, 
    2.100741e-07, 2.092967e-07, 2.089051e-07, 2.080852e-07, 2.08234e-07, 
    2.088362e-07, 2.102023e-07, 2.097384e-07, 2.109077e-07, 2.108813e-07, 
    2.121842e-07, 2.115966e-07, 2.137884e-07, 2.131651e-07, 2.149669e-07, 
    2.145136e-07, 2.149457e-07, 2.148146e-07, 2.149474e-07, 2.142825e-07, 
    2.145673e-07, 2.139824e-07, 2.117067e-07, 2.123751e-07, 2.103824e-07, 
    2.091857e-07, 2.083911e-07, 2.078277e-07, 2.079073e-07, 2.080592e-07, 
    2.088397e-07, 2.095739e-07, 2.101337e-07, 2.105083e-07, 2.108775e-07, 
    2.119957e-07, 2.125878e-07, 2.139145e-07, 2.136749e-07, 2.140807e-07, 
    2.144685e-07, 2.151198e-07, 2.150126e-07, 2.152996e-07, 2.1407e-07, 
    2.148871e-07, 2.135385e-07, 2.139072e-07, 2.109781e-07, 2.098635e-07, 
    2.093902e-07, 2.089759e-07, 2.079686e-07, 2.086641e-07, 2.083899e-07, 
    2.090424e-07, 2.094571e-07, 2.09252e-07, 2.105186e-07, 2.10026e-07, 
    2.126229e-07, 2.115037e-07, 2.144233e-07, 2.137241e-07, 2.145909e-07, 
    2.141485e-07, 2.149066e-07, 2.142243e-07, 2.154064e-07, 2.15664e-07, 
    2.15488e-07, 2.161642e-07, 2.141865e-07, 2.149457e-07, 2.092462e-07, 
    2.092797e-07, 2.094356e-07, 2.087505e-07, 2.087086e-07, 2.080811e-07, 
    2.086394e-07, 2.088773e-07, 2.094812e-07, 2.098385e-07, 2.101783e-07, 
    2.109256e-07, 2.117607e-07, 2.129293e-07, 2.137694e-07, 2.143328e-07, 
    2.139873e-07, 2.142923e-07, 2.139513e-07, 2.137915e-07, 2.155675e-07, 
    2.1457e-07, 2.160669e-07, 2.15984e-07, 2.153064e-07, 2.159934e-07, 
    2.093032e-07, 2.091107e-07, 2.084425e-07, 2.089653e-07, 2.080128e-07, 
    2.085459e-07, 2.088526e-07, 2.100364e-07, 2.102965e-07, 2.105379e-07, 
    2.110146e-07, 2.116267e-07, 2.127011e-07, 2.136366e-07, 2.14491e-07, 
    2.144284e-07, 2.144505e-07, 2.146414e-07, 2.141685e-07, 2.147191e-07, 
    2.148115e-07, 2.145699e-07, 2.159729e-07, 2.155719e-07, 2.159823e-07, 
    2.157212e-07, 2.091732e-07, 2.094972e-07, 2.093221e-07, 2.096514e-07, 
    2.094194e-07, 2.104511e-07, 2.107606e-07, 2.122095e-07, 2.116147e-07, 
    2.125615e-07, 2.117108e-07, 2.118615e-07, 2.125925e-07, 2.117567e-07, 
    2.13585e-07, 2.123453e-07, 2.146488e-07, 2.1341e-07, 2.147265e-07, 
    2.144873e-07, 2.148834e-07, 2.152382e-07, 2.156846e-07, 2.165089e-07, 
    2.163179e-07, 2.170075e-07, 2.099803e-07, 2.104008e-07, 2.103637e-07, 
    2.108039e-07, 2.111295e-07, 2.118354e-07, 2.129684e-07, 2.125422e-07, 
    2.133247e-07, 2.134818e-07, 2.122931e-07, 2.130229e-07, 2.106822e-07, 
    2.110602e-07, 2.108351e-07, 2.100135e-07, 2.126405e-07, 2.112917e-07, 
    2.137833e-07, 2.130518e-07, 2.151876e-07, 2.141251e-07, 2.162129e-07, 
    2.171065e-07, 2.179479e-07, 2.189321e-07, 2.106303e-07, 2.103445e-07, 
    2.108562e-07, 2.115645e-07, 2.122219e-07, 2.130965e-07, 2.131859e-07, 
    2.133498e-07, 2.137745e-07, 2.141316e-07, 2.134017e-07, 2.142212e-07, 
    2.11148e-07, 2.127576e-07, 2.102365e-07, 2.109953e-07, 2.115227e-07, 
    2.112913e-07, 2.124935e-07, 2.12777e-07, 2.139298e-07, 2.133337e-07, 
    2.168859e-07, 2.153132e-07, 2.196818e-07, 2.184595e-07, 2.102447e-07, 
    2.106293e-07, 2.119687e-07, 2.113312e-07, 2.131548e-07, 2.136041e-07, 
    2.139694e-07, 2.144365e-07, 2.144869e-07, 2.147638e-07, 2.143101e-07, 
    2.147459e-07, 2.130983e-07, 2.138343e-07, 2.118154e-07, 2.123066e-07, 
    2.120806e-07, 2.118328e-07, 2.125977e-07, 2.134132e-07, 2.134306e-07, 
    2.136922e-07, 2.144298e-07, 2.131622e-07, 2.170892e-07, 2.146628e-07, 
    2.110488e-07, 2.117902e-07, 2.11896e-07, 2.116088e-07, 2.13559e-07, 
    2.128521e-07, 2.147571e-07, 2.142419e-07, 2.15086e-07, 2.146665e-07, 
    2.146048e-07, 2.140662e-07, 2.13731e-07, 2.128845e-07, 2.121961e-07, 
    2.116504e-07, 2.117773e-07, 2.123768e-07, 2.134631e-07, 2.144915e-07, 
    2.142662e-07, 2.150219e-07, 2.130225e-07, 2.138606e-07, 2.135366e-07, 
    2.143814e-07, 2.125309e-07, 2.141068e-07, 2.121284e-07, 2.123018e-07, 
    2.12838e-07, 2.139175e-07, 2.141563e-07, 2.144115e-07, 2.14254e-07, 
    2.134907e-07, 2.133656e-07, 2.12825e-07, 2.126758e-07, 2.12264e-07, 
    2.119232e-07, 2.122346e-07, 2.125617e-07, 2.13491e-07, 2.14329e-07, 
    2.152432e-07, 2.15467e-07, 2.165364e-07, 2.156659e-07, 2.171027e-07, 
    2.158812e-07, 2.179963e-07, 2.141981e-07, 2.158452e-07, 2.128624e-07, 
    2.131834e-07, 2.137643e-07, 2.150974e-07, 2.143775e-07, 2.152194e-07, 
    2.133607e-07, 2.123975e-07, 2.121483e-07, 2.116836e-07, 2.121589e-07, 
    2.121202e-07, 2.125752e-07, 2.12429e-07, 2.135218e-07, 2.129347e-07, 
    2.146033e-07, 2.152127e-07, 2.169352e-07, 2.179923e-07, 2.190691e-07, 
    2.195448e-07, 2.196897e-07, 2.197502e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HTOP =
  0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 0.2411053, 
    0.2411053, 0.2411053 ;

 INT_SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAISHA =
  0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134, 0.001143134, 0.001143134, 
    0.001143134, 0.001143134, 0.001143134 ;

 LAISUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAKEICEFRAC =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAKEICETHICK =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAND_UPTAKE =
  6.358388e-08, 6.386347e-08, 6.380911e-08, 6.403462e-08, 6.390952e-08, 
    6.405718e-08, 6.364056e-08, 6.387457e-08, 6.372518e-08, 6.360905e-08, 
    6.447225e-08, 6.404468e-08, 6.491634e-08, 6.464366e-08, 6.532863e-08, 
    6.487392e-08, 6.542031e-08, 6.53155e-08, 6.563094e-08, 6.554057e-08, 
    6.594404e-08, 6.567264e-08, 6.615318e-08, 6.587923e-08, 6.592209e-08, 
    6.566369e-08, 6.413072e-08, 6.441902e-08, 6.411364e-08, 6.415475e-08, 
    6.41363e-08, 6.391211e-08, 6.379913e-08, 6.356251e-08, 6.360547e-08, 
    6.377926e-08, 6.417324e-08, 6.403949e-08, 6.437654e-08, 6.436893e-08, 
    6.474416e-08, 6.457498e-08, 6.520563e-08, 6.502638e-08, 6.554434e-08, 
    6.541408e-08, 6.553822e-08, 6.550058e-08, 6.553871e-08, 6.534768e-08, 
    6.542952e-08, 6.526142e-08, 6.460666e-08, 6.47991e-08, 6.422516e-08, 
    6.388007e-08, 6.365083e-08, 6.348817e-08, 6.351116e-08, 6.3555e-08, 
    6.378028e-08, 6.399208e-08, 6.415348e-08, 6.426145e-08, 6.436783e-08, 
    6.468986e-08, 6.486028e-08, 6.524188e-08, 6.5173e-08, 6.528968e-08, 
    6.540112e-08, 6.558825e-08, 6.555744e-08, 6.563989e-08, 6.528659e-08, 
    6.55214e-08, 6.513378e-08, 6.52398e-08, 6.439678e-08, 6.407557e-08, 
    6.393907e-08, 6.381956e-08, 6.352884e-08, 6.372961e-08, 6.365047e-08, 
    6.383875e-08, 6.395839e-08, 6.389921e-08, 6.426441e-08, 6.412242e-08, 
    6.487038e-08, 6.454822e-08, 6.538812e-08, 6.518714e-08, 6.54363e-08, 
    6.530916e-08, 6.5527e-08, 6.533094e-08, 6.567057e-08, 6.574452e-08, 
    6.569399e-08, 6.588811e-08, 6.532007e-08, 6.553822e-08, 6.389756e-08, 
    6.390721e-08, 6.395216e-08, 6.375454e-08, 6.374245e-08, 6.356133e-08, 
    6.372249e-08, 6.379111e-08, 6.396532e-08, 6.406837e-08, 6.416632e-08, 
    6.438169e-08, 6.462222e-08, 6.495855e-08, 6.520017e-08, 6.536213e-08, 
    6.526282e-08, 6.53505e-08, 6.525248e-08, 6.520654e-08, 6.571682e-08, 
    6.543029e-08, 6.586019e-08, 6.58364e-08, 6.564185e-08, 6.583908e-08, 
    6.391399e-08, 6.385844e-08, 6.366564e-08, 6.381653e-08, 6.354161e-08, 
    6.36955e-08, 6.378399e-08, 6.41254e-08, 6.420041e-08, 6.426996e-08, 
    6.440733e-08, 6.458363e-08, 6.489289e-08, 6.516198e-08, 6.54076e-08, 
    6.538961e-08, 6.539594e-08, 6.545082e-08, 6.531489e-08, 6.547314e-08, 
    6.54997e-08, 6.543026e-08, 6.583321e-08, 6.571809e-08, 6.58359e-08, 
    6.576094e-08, 6.38765e-08, 6.396994e-08, 6.391945e-08, 6.40144e-08, 
    6.394751e-08, 6.424496e-08, 6.433414e-08, 6.475143e-08, 6.458016e-08, 
    6.485271e-08, 6.460785e-08, 6.465124e-08, 6.486162e-08, 6.462108e-08, 
    6.514714e-08, 6.47905e-08, 6.545295e-08, 6.509682e-08, 6.547527e-08, 
    6.540655e-08, 6.552033e-08, 6.562224e-08, 6.575045e-08, 6.598701e-08, 
    6.593223e-08, 6.613006e-08, 6.410925e-08, 6.423046e-08, 6.421978e-08, 
    6.434662e-08, 6.444042e-08, 6.464373e-08, 6.496981e-08, 6.484719e-08, 
    6.507229e-08, 6.511748e-08, 6.477549e-08, 6.498548e-08, 6.431157e-08, 
    6.442045e-08, 6.435562e-08, 6.411882e-08, 6.487545e-08, 6.448715e-08, 
    6.520416e-08, 6.499381e-08, 6.560771e-08, 6.530242e-08, 6.590207e-08, 
    6.615844e-08, 6.639969e-08, 6.668164e-08, 6.42966e-08, 6.421424e-08, 
    6.43617e-08, 6.456572e-08, 6.4755e-08, 6.500665e-08, 6.503239e-08, 
    6.507953e-08, 6.520164e-08, 6.530431e-08, 6.509445e-08, 6.533005e-08, 
    6.444572e-08, 6.490915e-08, 6.418311e-08, 6.440175e-08, 6.455369e-08, 
    6.448703e-08, 6.483317e-08, 6.491475e-08, 6.524627e-08, 6.507489e-08, 
    6.609517e-08, 6.564377e-08, 6.689631e-08, 6.654629e-08, 6.418547e-08, 
    6.429631e-08, 6.468208e-08, 6.449854e-08, 6.502344e-08, 6.515264e-08, 
    6.525767e-08, 6.539194e-08, 6.540643e-08, 6.548598e-08, 6.535562e-08, 
    6.548083e-08, 6.500718e-08, 6.521884e-08, 6.463799e-08, 6.477936e-08, 
    6.471433e-08, 6.464298e-08, 6.486317e-08, 6.509775e-08, 6.510275e-08, 
    6.517797e-08, 6.538995e-08, 6.502557e-08, 6.615345e-08, 6.545692e-08, 
    6.441718e-08, 6.463069e-08, 6.466117e-08, 6.457847e-08, 6.513969e-08, 
    6.493634e-08, 6.548404e-08, 6.533602e-08, 6.557855e-08, 6.545803e-08, 
    6.54403e-08, 6.528551e-08, 6.518914e-08, 6.494567e-08, 6.474756e-08, 
    6.459047e-08, 6.4627e-08, 6.479956e-08, 6.51121e-08, 6.540775e-08, 
    6.534299e-08, 6.556012e-08, 6.498538e-08, 6.522639e-08, 6.513324e-08, 
    6.537611e-08, 6.484393e-08, 6.529714e-08, 6.472809e-08, 6.477798e-08, 
    6.493231e-08, 6.524274e-08, 6.53114e-08, 6.538474e-08, 6.533948e-08, 
    6.512003e-08, 6.508407e-08, 6.492856e-08, 6.488562e-08, 6.476711e-08, 
    6.466901e-08, 6.475865e-08, 6.485278e-08, 6.512012e-08, 6.536104e-08, 
    6.562369e-08, 6.568797e-08, 6.599488e-08, 6.574506e-08, 6.615733e-08, 
    6.580684e-08, 6.641355e-08, 6.532339e-08, 6.579651e-08, 6.493933e-08, 
    6.503167e-08, 6.519871e-08, 6.558179e-08, 6.537497e-08, 6.561685e-08, 
    6.508266e-08, 6.480552e-08, 6.47338e-08, 6.460002e-08, 6.473686e-08, 
    6.472573e-08, 6.485668e-08, 6.48146e-08, 6.512899e-08, 6.496011e-08, 
    6.543986e-08, 6.561493e-08, 6.610933e-08, 6.641241e-08, 6.672092e-08, 
    6.685712e-08, 6.689857e-08, 6.69159e-08 ;

 LAND_USE_FLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC =
  0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 0.1428187, 
    0.1428187, 0.1428187 ;

 LEAFC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC_LOSS =
  8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 8.453753e-10, 
    8.453753e-10, 8.453753e-10, 8.453753e-10 ;

 LEAFN =
  0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469, 0.003570469, 0.003570469, 
    0.003570469, 0.003570469, 0.003570469 ;

 LEAF_MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LFC2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LF_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITFALL =
  1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 1.322607e-09, 
    1.322607e-09, 1.322607e-09, 1.322607e-09 ;

 LITHR =
  9.028442e-13, 9.052879e-13, 9.048132e-13, 9.067824e-13, 9.056906e-13, 
    9.069795e-13, 9.033402e-13, 9.053846e-13, 9.040799e-13, 9.030648e-13, 
    9.105982e-13, 9.068703e-13, 9.144674e-13, 9.120941e-13, 9.180519e-13, 
    9.140977e-13, 9.188485e-13, 9.179387e-13, 9.20678e-13, 9.198936e-13, 
    9.233922e-13, 9.2104e-13, 9.252049e-13, 9.22831e-13, 9.232023e-13, 
    9.209622e-13, 9.076217e-13, 9.101342e-13, 9.074726e-13, 9.078311e-13, 
    9.076704e-13, 9.057128e-13, 9.047252e-13, 9.026579e-13, 9.030335e-13, 
    9.045521e-13, 9.079923e-13, 9.068256e-13, 9.097664e-13, 9.097e-13, 
    9.129694e-13, 9.114959e-13, 9.169837e-13, 9.154259e-13, 9.199265e-13, 
    9.187952e-13, 9.198731e-13, 9.195464e-13, 9.198775e-13, 9.182181e-13, 
    9.189291e-13, 9.174688e-13, 9.117717e-13, 9.134475e-13, 9.084456e-13, 
    9.054318e-13, 9.034297e-13, 9.020075e-13, 9.022086e-13, 9.025918e-13, 
    9.045609e-13, 9.064116e-13, 9.078206e-13, 9.087626e-13, 9.096905e-13, 
    9.124949e-13, 9.139795e-13, 9.172984e-13, 9.167003e-13, 9.177138e-13, 
    9.186827e-13, 9.203073e-13, 9.200401e-13, 9.207554e-13, 9.176876e-13, 
    9.197266e-13, 9.163595e-13, 9.172809e-13, 9.099401e-13, 9.071405e-13, 
    9.059473e-13, 9.049044e-13, 9.023632e-13, 9.041183e-13, 9.034265e-13, 
    9.050725e-13, 9.061174e-13, 9.056007e-13, 9.087884e-13, 9.075495e-13, 
    9.140674e-13, 9.112623e-13, 9.185697e-13, 9.168231e-13, 9.189882e-13, 
    9.178838e-13, 9.197755e-13, 9.180731e-13, 9.210217e-13, 9.21663e-13, 
    9.212248e-13, 9.229087e-13, 9.179786e-13, 9.198729e-13, 9.055861e-13, 
    9.056703e-13, 9.060631e-13, 9.043361e-13, 9.042305e-13, 9.026474e-13, 
    9.040563e-13, 9.046559e-13, 9.061781e-13, 9.070776e-13, 9.079325e-13, 
    9.098111e-13, 9.119069e-13, 9.14835e-13, 9.169363e-13, 9.183441e-13, 
    9.174812e-13, 9.18243e-13, 9.173913e-13, 9.169921e-13, 9.214226e-13, 
    9.189356e-13, 9.226666e-13, 9.224604e-13, 9.207722e-13, 9.224837e-13, 
    9.057296e-13, 9.052446e-13, 9.035593e-13, 9.048783e-13, 9.02475e-13, 
    9.038203e-13, 9.045932e-13, 9.075749e-13, 9.082301e-13, 9.088366e-13, 
    9.100349e-13, 9.115713e-13, 9.142639e-13, 9.16604e-13, 9.187392e-13, 
    9.185828e-13, 9.186378e-13, 9.191142e-13, 9.179335e-13, 9.19308e-13, 
    9.195383e-13, 9.189356e-13, 9.224327e-13, 9.214343e-13, 9.22456e-13, 
    9.218059e-13, 9.054023e-13, 9.062184e-13, 9.057774e-13, 9.066063e-13, 
    9.060222e-13, 9.086179e-13, 9.093956e-13, 9.130319e-13, 9.115409e-13, 
    9.13914e-13, 9.117823e-13, 9.1216e-13, 9.139903e-13, 9.118977e-13, 
    9.164746e-13, 9.133717e-13, 9.191327e-13, 9.160368e-13, 9.193266e-13, 
    9.187298e-13, 9.19718e-13, 9.206024e-13, 9.217149e-13, 9.237654e-13, 
    9.232908e-13, 9.250051e-13, 9.074346e-13, 9.084918e-13, 9.083992e-13, 
    9.095054e-13, 9.103231e-13, 9.120951e-13, 9.149334e-13, 9.138666e-13, 
    9.158252e-13, 9.162176e-13, 9.132426e-13, 9.150695e-13, 9.091994e-13, 
    9.101483e-13, 9.095837e-13, 9.075177e-13, 9.141118e-13, 9.107297e-13, 
    9.16971e-13, 9.151424e-13, 9.204762e-13, 9.178244e-13, 9.230294e-13, 
    9.252496e-13, 9.273394e-13, 9.297761e-13, 9.09069e-13, 9.083509e-13, 
    9.096371e-13, 9.114145e-13, 9.130638e-13, 9.152539e-13, 9.154781e-13, 
    9.15888e-13, 9.169495e-13, 9.178416e-13, 9.16017e-13, 9.180653e-13, 
    9.103673e-13, 9.144054e-13, 9.080788e-13, 9.099851e-13, 9.1131e-13, 
    9.107294e-13, 9.137448e-13, 9.144547e-13, 9.173367e-13, 9.158479e-13, 
    9.247014e-13, 9.207883e-13, 9.316315e-13, 9.286064e-13, 9.080998e-13, 
    9.090668e-13, 9.124286e-13, 9.108298e-13, 9.154002e-13, 9.165232e-13, 
    9.174365e-13, 9.186025e-13, 9.187289e-13, 9.194195e-13, 9.182876e-13, 
    9.193749e-13, 9.152585e-13, 9.170989e-13, 9.120451e-13, 9.13276e-13, 
    9.1271e-13, 9.120887e-13, 9.140057e-13, 9.160457e-13, 9.160901e-13, 
    9.167431e-13, 9.185824e-13, 9.154188e-13, 9.252044e-13, 9.191644e-13, 
    9.101208e-13, 9.119803e-13, 9.122468e-13, 9.115266e-13, 9.164106e-13, 
    9.146423e-13, 9.194028e-13, 9.181171e-13, 9.202234e-13, 9.19177e-13, 
    9.190229e-13, 9.176784e-13, 9.168406e-13, 9.147233e-13, 9.12999e-13, 
    9.116311e-13, 9.119493e-13, 9.134516e-13, 9.161706e-13, 9.187399e-13, 
    9.181771e-13, 9.200634e-13, 9.150691e-13, 9.171639e-13, 9.163541e-13, 
    9.184654e-13, 9.13838e-13, 9.177765e-13, 9.128299e-13, 9.132643e-13, 
    9.146073e-13, 9.173055e-13, 9.179033e-13, 9.1854e-13, 9.181473e-13, 
    9.162392e-13, 9.159274e-13, 9.145747e-13, 9.142008e-13, 9.131697e-13, 
    9.123154e-13, 9.130958e-13, 9.139149e-13, 9.162404e-13, 9.18334e-13, 
    9.206148e-13, 9.211729e-13, 9.238321e-13, 9.216665e-13, 9.252378e-13, 
    9.222001e-13, 9.274567e-13, 9.180057e-13, 9.221124e-13, 9.146686e-13, 
    9.154719e-13, 9.169229e-13, 9.202503e-13, 9.184554e-13, 9.205548e-13, 
    9.159151e-13, 9.135031e-13, 9.128796e-13, 9.117142e-13, 9.129063e-13, 
    9.128093e-13, 9.139494e-13, 9.135831e-13, 9.163176e-13, 9.148495e-13, 
    9.190188e-13, 9.205384e-13, 9.248251e-13, 9.274484e-13, 9.301169e-13, 
    9.312933e-13, 9.316515e-13, 9.318011e-13 ;

 LITR1C =
  3.186876e-05, 3.186863e-05, 3.186865e-05, 3.186855e-05, 3.186861e-05, 
    3.186855e-05, 3.186873e-05, 3.186863e-05, 3.186869e-05, 3.186875e-05, 
    3.186836e-05, 3.186855e-05, 3.186816e-05, 3.186828e-05, 3.186797e-05, 
    3.186817e-05, 3.186793e-05, 3.186798e-05, 3.186784e-05, 3.186788e-05, 
    3.186769e-05, 3.186782e-05, 3.18676e-05, 3.186772e-05, 3.18677e-05, 
    3.186782e-05, 3.186851e-05, 3.186838e-05, 3.186852e-05, 3.18685e-05, 
    3.186851e-05, 3.186861e-05, 3.186866e-05, 3.186877e-05, 3.186875e-05, 
    3.186867e-05, 3.186849e-05, 3.186855e-05, 3.18684e-05, 3.18684e-05, 
    3.186823e-05, 3.186831e-05, 3.186802e-05, 3.186811e-05, 3.186788e-05, 
    3.186793e-05, 3.186788e-05, 3.186789e-05, 3.186788e-05, 3.186796e-05, 
    3.186793e-05, 3.1868e-05, 3.186829e-05, 3.186821e-05, 3.186847e-05, 
    3.186862e-05, 3.186873e-05, 3.18688e-05, 3.186879e-05, 3.186877e-05, 
    3.186867e-05, 3.186857e-05, 3.18685e-05, 3.186845e-05, 3.18684e-05, 
    3.186826e-05, 3.186818e-05, 3.186801e-05, 3.186804e-05, 3.186799e-05, 
    3.186794e-05, 3.186785e-05, 3.186787e-05, 3.186783e-05, 3.186799e-05, 
    3.186788e-05, 3.186806e-05, 3.186801e-05, 3.186839e-05, 3.186853e-05, 
    3.18686e-05, 3.186865e-05, 3.186878e-05, 3.186869e-05, 3.186873e-05, 
    3.186864e-05, 3.186859e-05, 3.186861e-05, 3.186845e-05, 3.186851e-05, 
    3.186818e-05, 3.186832e-05, 3.186794e-05, 3.186804e-05, 3.186792e-05, 
    3.186798e-05, 3.186788e-05, 3.186797e-05, 3.186782e-05, 3.186778e-05, 
    3.186781e-05, 3.186772e-05, 3.186797e-05, 3.186788e-05, 3.186861e-05, 
    3.186861e-05, 3.186859e-05, 3.186868e-05, 3.186869e-05, 3.186877e-05, 
    3.186869e-05, 3.186867e-05, 3.186859e-05, 3.186854e-05, 3.186849e-05, 
    3.18684e-05, 3.186829e-05, 3.186814e-05, 3.186803e-05, 3.186796e-05, 
    3.1868e-05, 3.186796e-05, 3.186801e-05, 3.186802e-05, 3.18678e-05, 
    3.186793e-05, 3.186773e-05, 3.186774e-05, 3.186783e-05, 3.186774e-05, 
    3.186861e-05, 3.186863e-05, 3.186872e-05, 3.186865e-05, 3.186878e-05, 
    3.186871e-05, 3.186867e-05, 3.186851e-05, 3.186848e-05, 3.186845e-05, 
    3.186839e-05, 3.186831e-05, 3.186817e-05, 3.186805e-05, 3.186793e-05, 
    3.186794e-05, 3.186794e-05, 3.186792e-05, 3.186798e-05, 3.18679e-05, 
    3.186789e-05, 3.186793e-05, 3.186774e-05, 3.18678e-05, 3.186774e-05, 
    3.186778e-05, 3.186863e-05, 3.186858e-05, 3.186861e-05, 3.186856e-05, 
    3.186859e-05, 3.186846e-05, 3.186842e-05, 3.186823e-05, 3.186831e-05, 
    3.186819e-05, 3.186829e-05, 3.186828e-05, 3.186818e-05, 3.186829e-05, 
    3.186805e-05, 3.186821e-05, 3.186792e-05, 3.186808e-05, 3.18679e-05, 
    3.186794e-05, 3.186789e-05, 3.186784e-05, 3.186778e-05, 3.186768e-05, 
    3.18677e-05, 3.186761e-05, 3.186852e-05, 3.186847e-05, 3.186847e-05, 
    3.186841e-05, 3.186837e-05, 3.186828e-05, 3.186813e-05, 3.186819e-05, 
    3.186809e-05, 3.186806e-05, 3.186822e-05, 3.186813e-05, 3.186843e-05, 
    3.186838e-05, 3.186841e-05, 3.186852e-05, 3.186817e-05, 3.186835e-05, 
    3.186803e-05, 3.186812e-05, 3.186785e-05, 3.186798e-05, 3.186772e-05, 
    3.18676e-05, 3.186749e-05, 3.186737e-05, 3.186844e-05, 3.186847e-05, 
    3.186841e-05, 3.186831e-05, 3.186823e-05, 3.186812e-05, 3.18681e-05, 
    3.186808e-05, 3.186803e-05, 3.186798e-05, 3.186808e-05, 3.186797e-05, 
    3.186837e-05, 3.186816e-05, 3.186849e-05, 3.186839e-05, 3.186832e-05, 
    3.186835e-05, 3.186819e-05, 3.186816e-05, 3.186801e-05, 3.186809e-05, 
    3.186763e-05, 3.186783e-05, 3.186727e-05, 3.186742e-05, 3.186849e-05, 
    3.186844e-05, 3.186826e-05, 3.186835e-05, 3.186811e-05, 3.186805e-05, 
    3.1868e-05, 3.186794e-05, 3.186794e-05, 3.18679e-05, 3.186796e-05, 
    3.18679e-05, 3.186812e-05, 3.186802e-05, 3.186828e-05, 3.186822e-05, 
    3.186825e-05, 3.186828e-05, 3.186818e-05, 3.186808e-05, 3.186807e-05, 
    3.186804e-05, 3.186794e-05, 3.186811e-05, 3.18676e-05, 3.186791e-05, 
    3.186838e-05, 3.186828e-05, 3.186827e-05, 3.186831e-05, 3.186806e-05, 
    3.186815e-05, 3.18679e-05, 3.186797e-05, 3.186786e-05, 3.186791e-05, 
    3.186792e-05, 3.186799e-05, 3.186803e-05, 3.186814e-05, 3.186823e-05, 
    3.18683e-05, 3.186829e-05, 3.186821e-05, 3.186807e-05, 3.186793e-05, 
    3.186796e-05, 3.186787e-05, 3.186813e-05, 3.186802e-05, 3.186806e-05, 
    3.186795e-05, 3.186819e-05, 3.186798e-05, 3.186824e-05, 3.186822e-05, 
    3.186815e-05, 3.186801e-05, 3.186798e-05, 3.186794e-05, 3.186797e-05, 
    3.186806e-05, 3.186808e-05, 3.186815e-05, 3.186817e-05, 3.186823e-05, 
    3.186827e-05, 3.186823e-05, 3.186819e-05, 3.186806e-05, 3.186796e-05, 
    3.186784e-05, 3.186781e-05, 3.186767e-05, 3.186778e-05, 3.18676e-05, 
    3.186776e-05, 3.186749e-05, 3.186797e-05, 3.186776e-05, 3.186815e-05, 
    3.18681e-05, 3.186803e-05, 3.186786e-05, 3.186795e-05, 3.186784e-05, 
    3.186808e-05, 3.186821e-05, 3.186824e-05, 3.18683e-05, 3.186824e-05, 
    3.186824e-05, 3.186818e-05, 3.18682e-05, 3.186806e-05, 3.186814e-05, 
    3.186792e-05, 3.186784e-05, 3.186762e-05, 3.186749e-05, 3.186735e-05, 
    3.186729e-05, 3.186727e-05, 3.186726e-05 ;

 LITR1C_TO_SOIL1C =
  6.013331e-13, 6.029604e-13, 6.026443e-13, 6.039556e-13, 6.032286e-13, 
    6.040869e-13, 6.016634e-13, 6.030248e-13, 6.02156e-13, 6.0148e-13, 
    6.064967e-13, 6.040142e-13, 6.090732e-13, 6.074928e-13, 6.114602e-13, 
    6.088271e-13, 6.119907e-13, 6.113848e-13, 6.13209e-13, 6.126867e-13, 
    6.150163e-13, 6.1345e-13, 6.162235e-13, 6.146427e-13, 6.148899e-13, 
    6.133982e-13, 6.045146e-13, 6.061876e-13, 6.044153e-13, 6.04654e-13, 
    6.04547e-13, 6.032434e-13, 6.025857e-13, 6.01209e-13, 6.014591e-13, 
    6.024704e-13, 6.047614e-13, 6.039844e-13, 6.059428e-13, 6.058986e-13, 
    6.080756e-13, 6.070945e-13, 6.107489e-13, 6.097115e-13, 6.127085e-13, 
    6.119551e-13, 6.12673e-13, 6.124555e-13, 6.126758e-13, 6.115709e-13, 
    6.120444e-13, 6.110719e-13, 6.072782e-13, 6.08394e-13, 6.050633e-13, 
    6.030562e-13, 6.01723e-13, 6.007759e-13, 6.009099e-13, 6.011651e-13, 
    6.024763e-13, 6.037087e-13, 6.04647e-13, 6.052743e-13, 6.058922e-13, 
    6.077597e-13, 6.087483e-13, 6.109584e-13, 6.105602e-13, 6.112351e-13, 
    6.118802e-13, 6.129621e-13, 6.127841e-13, 6.132605e-13, 6.112176e-13, 
    6.125755e-13, 6.103332e-13, 6.109467e-13, 6.060584e-13, 6.041941e-13, 
    6.033995e-13, 6.027051e-13, 6.010128e-13, 6.021816e-13, 6.017209e-13, 
    6.02817e-13, 6.035128e-13, 6.031687e-13, 6.052915e-13, 6.044665e-13, 
    6.088069e-13, 6.069389e-13, 6.11805e-13, 6.10642e-13, 6.120837e-13, 
    6.113483e-13, 6.12608e-13, 6.114743e-13, 6.134378e-13, 6.138649e-13, 
    6.13573e-13, 6.146944e-13, 6.114114e-13, 6.126728e-13, 6.03159e-13, 
    6.032151e-13, 6.034767e-13, 6.023266e-13, 6.022563e-13, 6.012021e-13, 
    6.021403e-13, 6.025396e-13, 6.035532e-13, 6.041522e-13, 6.047215e-13, 
    6.059725e-13, 6.073682e-13, 6.093181e-13, 6.107174e-13, 6.116548e-13, 
    6.110801e-13, 6.115874e-13, 6.110202e-13, 6.107544e-13, 6.137048e-13, 
    6.120487e-13, 6.145332e-13, 6.143958e-13, 6.132717e-13, 6.144114e-13, 
    6.032545e-13, 6.029316e-13, 6.018093e-13, 6.026877e-13, 6.010873e-13, 
    6.019831e-13, 6.024978e-13, 6.044834e-13, 6.049197e-13, 6.053236e-13, 
    6.061215e-13, 6.071447e-13, 6.089377e-13, 6.104961e-13, 6.119178e-13, 
    6.118137e-13, 6.118504e-13, 6.121676e-13, 6.113814e-13, 6.122967e-13, 
    6.1245e-13, 6.120487e-13, 6.143775e-13, 6.137125e-13, 6.143929e-13, 
    6.139601e-13, 6.030366e-13, 6.0358e-13, 6.032864e-13, 6.038384e-13, 
    6.034494e-13, 6.05178e-13, 6.056958e-13, 6.081173e-13, 6.071244e-13, 
    6.087048e-13, 6.072852e-13, 6.075367e-13, 6.087555e-13, 6.07362e-13, 
    6.104098e-13, 6.083436e-13, 6.1218e-13, 6.101183e-13, 6.12309e-13, 
    6.119117e-13, 6.125697e-13, 6.131586e-13, 6.138994e-13, 6.152649e-13, 
    6.149489e-13, 6.160904e-13, 6.043899e-13, 6.050939e-13, 6.050323e-13, 
    6.05769e-13, 6.063134e-13, 6.074934e-13, 6.093835e-13, 6.086732e-13, 
    6.099775e-13, 6.102387e-13, 6.082576e-13, 6.094742e-13, 6.055651e-13, 
    6.061971e-13, 6.058211e-13, 6.044453e-13, 6.088364e-13, 6.065842e-13, 
    6.107404e-13, 6.095227e-13, 6.130746e-13, 6.113087e-13, 6.147748e-13, 
    6.162532e-13, 6.176448e-13, 6.192675e-13, 6.054784e-13, 6.050001e-13, 
    6.058566e-13, 6.070402e-13, 6.081385e-13, 6.09597e-13, 6.097463e-13, 
    6.100192e-13, 6.10726e-13, 6.113202e-13, 6.101052e-13, 6.114692e-13, 
    6.063429e-13, 6.090319e-13, 6.04819e-13, 6.060884e-13, 6.069706e-13, 
    6.06584e-13, 6.08592e-13, 6.090648e-13, 6.109839e-13, 6.099925e-13, 
    6.158881e-13, 6.132824e-13, 6.20503e-13, 6.184886e-13, 6.048329e-13, 
    6.054769e-13, 6.077155e-13, 6.066509e-13, 6.096944e-13, 6.104422e-13, 
    6.110504e-13, 6.118269e-13, 6.11911e-13, 6.123709e-13, 6.116171e-13, 
    6.123412e-13, 6.096e-13, 6.108255e-13, 6.074602e-13, 6.082799e-13, 
    6.079029e-13, 6.074892e-13, 6.087658e-13, 6.101243e-13, 6.101538e-13, 
    6.105887e-13, 6.118134e-13, 6.097068e-13, 6.162231e-13, 6.12201e-13, 
    6.061787e-13, 6.074171e-13, 6.075945e-13, 6.071149e-13, 6.103672e-13, 
    6.091897e-13, 6.123597e-13, 6.115037e-13, 6.129062e-13, 6.122094e-13, 
    6.121068e-13, 6.112114e-13, 6.106536e-13, 6.092436e-13, 6.080954e-13, 
    6.071845e-13, 6.073964e-13, 6.083968e-13, 6.102074e-13, 6.119183e-13, 
    6.115435e-13, 6.127997e-13, 6.09474e-13, 6.108689e-13, 6.103296e-13, 
    6.117355e-13, 6.086541e-13, 6.112768e-13, 6.079827e-13, 6.08272e-13, 
    6.091663e-13, 6.109631e-13, 6.113612e-13, 6.117853e-13, 6.115237e-13, 
    6.102531e-13, 6.100454e-13, 6.091447e-13, 6.088957e-13, 6.082091e-13, 
    6.076401e-13, 6.081598e-13, 6.087053e-13, 6.102539e-13, 6.11648e-13, 
    6.131669e-13, 6.135385e-13, 6.153093e-13, 6.138672e-13, 6.162454e-13, 
    6.142226e-13, 6.177229e-13, 6.114295e-13, 6.141642e-13, 6.092072e-13, 
    6.097422e-13, 6.107084e-13, 6.129242e-13, 6.117289e-13, 6.131269e-13, 
    6.100373e-13, 6.084311e-13, 6.080159e-13, 6.072398e-13, 6.080336e-13, 
    6.079691e-13, 6.087282e-13, 6.084843e-13, 6.103053e-13, 6.093276e-13, 
    6.121041e-13, 6.13116e-13, 6.159706e-13, 6.177175e-13, 6.194944e-13, 
    6.202779e-13, 6.205163e-13, 6.206159e-13 ;

 LITR1C_vr =
  0.001819739, 0.001819732, 0.001819733, 0.001819727, 0.001819731, 
    0.001819727, 0.001819737, 0.001819731, 0.001819735, 0.001819738, 
    0.001819716, 0.001819727, 0.001819705, 0.001819712, 0.001819694, 
    0.001819706, 0.001819692, 0.001819694, 0.001819686, 0.001819689, 
    0.001819678, 0.001819685, 0.001819673, 0.00181968, 0.001819679, 
    0.001819685, 0.001819725, 0.001819717, 0.001819725, 0.001819724, 
    0.001819725, 0.001819731, 0.001819733, 0.001819739, 0.001819738, 
    0.001819734, 0.001819724, 0.001819727, 0.001819719, 0.001819719, 
    0.001819709, 0.001819713, 0.001819697, 0.001819702, 0.001819689, 
    0.001819692, 0.001819689, 0.00181969, 0.001819689, 0.001819694, 
    0.001819692, 0.001819696, 0.001819713, 0.001819708, 0.001819722, 
    0.001819731, 0.001819737, 0.001819741, 0.001819741, 0.00181974, 
    0.001819734, 0.001819728, 0.001819724, 0.001819722, 0.001819719, 
    0.00181971, 0.001819706, 0.001819696, 0.001819698, 0.001819695, 
    0.001819692, 0.001819687, 0.001819688, 0.001819686, 0.001819695, 
    0.001819689, 0.001819699, 0.001819696, 0.001819718, 0.001819726, 
    0.00181973, 0.001819733, 0.00181974, 0.001819735, 0.001819737, 
    0.001819732, 0.001819729, 0.001819731, 0.001819721, 0.001819725, 
    0.001819706, 0.001819714, 0.001819693, 0.001819698, 0.001819691, 
    0.001819695, 0.001819689, 0.001819694, 0.001819685, 0.001819683, 
    0.001819685, 0.00181968, 0.001819694, 0.001819689, 0.001819731, 
    0.001819731, 0.001819729, 0.001819735, 0.001819735, 0.00181974, 
    0.001819735, 0.001819734, 0.001819729, 0.001819726, 0.001819724, 
    0.001819718, 0.001819712, 0.001819704, 0.001819697, 0.001819693, 
    0.001819696, 0.001819693, 0.001819696, 0.001819697, 0.001819684, 
    0.001819692, 0.00181968, 0.001819681, 0.001819686, 0.001819681, 
    0.001819731, 0.001819732, 0.001819737, 0.001819733, 0.00181974, 
    0.001819736, 0.001819734, 0.001819725, 0.001819723, 0.001819721, 
    0.001819718, 0.001819713, 0.001819705, 0.001819698, 0.001819692, 
    0.001819693, 0.001819692, 0.001819691, 0.001819694, 0.00181969, 
    0.00181969, 0.001819692, 0.001819681, 0.001819684, 0.001819681, 
    0.001819683, 0.001819731, 0.001819729, 0.00181973, 0.001819728, 
    0.00181973, 0.001819722, 0.00181972, 0.001819709, 0.001819713, 
    0.001819706, 0.001819713, 0.001819712, 0.001819706, 0.001819712, 
    0.001819699, 0.001819708, 0.001819691, 0.0018197, 0.00181969, 
    0.001819692, 0.001819689, 0.001819687, 0.001819683, 0.001819677, 
    0.001819679, 0.001819674, 0.001819725, 0.001819722, 0.001819723, 
    0.001819719, 0.001819717, 0.001819712, 0.001819703, 0.001819706, 
    0.001819701, 0.0018197, 0.001819708, 0.001819703, 0.00181972, 
    0.001819717, 0.001819719, 0.001819725, 0.001819706, 0.001819716, 
    0.001819697, 0.001819703, 0.001819687, 0.001819695, 0.001819679, 
    0.001819673, 0.001819667, 0.001819659, 0.001819721, 0.001819723, 
    0.001819719, 0.001819714, 0.001819709, 0.001819702, 0.001819702, 
    0.0018197, 0.001819697, 0.001819695, 0.0018197, 0.001819694, 0.001819717, 
    0.001819705, 0.001819724, 0.001819718, 0.001819714, 0.001819716, 
    0.001819707, 0.001819705, 0.001819696, 0.001819701, 0.001819675, 
    0.001819686, 0.001819654, 0.001819663, 0.001819723, 0.001819721, 
    0.001819711, 0.001819715, 0.001819702, 0.001819699, 0.001819696, 
    0.001819692, 0.001819692, 0.00181969, 0.001819693, 0.00181969, 
    0.001819702, 0.001819697, 0.001819712, 0.001819708, 0.00181971, 
    0.001819712, 0.001819706, 0.0018197, 0.0018197, 0.001819698, 0.001819693, 
    0.001819702, 0.001819673, 0.001819691, 0.001819717, 0.001819712, 
    0.001819711, 0.001819713, 0.001819699, 0.001819704, 0.00181969, 
    0.001819694, 0.001819688, 0.001819691, 0.001819691, 0.001819695, 
    0.001819698, 0.001819704, 0.001819709, 0.001819713, 0.001819712, 
    0.001819708, 0.0018197, 0.001819692, 0.001819694, 0.001819688, 
    0.001819703, 0.001819697, 0.001819699, 0.001819693, 0.001819707, 
    0.001819695, 0.00181971, 0.001819708, 0.001819704, 0.001819696, 
    0.001819695, 0.001819693, 0.001819694, 0.001819699, 0.0018197, 
    0.001819704, 0.001819705, 0.001819709, 0.001819711, 0.001819709, 
    0.001819706, 0.001819699, 0.001819693, 0.001819686, 0.001819685, 
    0.001819677, 0.001819683, 0.001819673, 0.001819682, 0.001819666, 
    0.001819694, 0.001819682, 0.001819704, 0.001819702, 0.001819697, 
    0.001819688, 0.001819693, 0.001819687, 0.0018197, 0.001819707, 
    0.001819709, 0.001819713, 0.001819709, 0.00181971, 0.001819706, 
    0.001819707, 0.001819699, 0.001819703, 0.001819691, 0.001819687, 
    0.001819674, 0.001819666, 0.001819658, 0.001819655, 0.001819654, 
    0.001819654,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N =
  1.011397e-06, 1.011393e-06, 1.011394e-06, 1.01139e-06, 1.011392e-06, 
    1.01139e-06, 1.011396e-06, 1.011393e-06, 1.011395e-06, 1.011396e-06, 
    1.011384e-06, 1.01139e-06, 1.011378e-06, 1.011382e-06, 1.011372e-06, 
    1.011378e-06, 1.011371e-06, 1.011372e-06, 1.011368e-06, 1.011369e-06, 
    1.011363e-06, 1.011367e-06, 1.01136e-06, 1.011364e-06, 1.011363e-06, 
    1.011367e-06, 1.011389e-06, 1.011385e-06, 1.011389e-06, 1.011389e-06, 
    1.011389e-06, 1.011392e-06, 1.011394e-06, 1.011397e-06, 1.011396e-06, 
    1.011394e-06, 1.011388e-06, 1.01139e-06, 1.011385e-06, 1.011386e-06, 
    1.01138e-06, 1.011383e-06, 1.011374e-06, 1.011376e-06, 1.011369e-06, 
    1.011371e-06, 1.011369e-06, 1.011369e-06, 1.011369e-06, 1.011372e-06, 
    1.01137e-06, 1.011373e-06, 1.011382e-06, 1.011379e-06, 1.011388e-06, 
    1.011393e-06, 1.011396e-06, 1.011398e-06, 1.011398e-06, 1.011397e-06, 
    1.011394e-06, 1.011391e-06, 1.011389e-06, 1.011387e-06, 1.011386e-06, 
    1.011381e-06, 1.011378e-06, 1.011373e-06, 1.011374e-06, 1.011372e-06, 
    1.011371e-06, 1.011368e-06, 1.011369e-06, 1.011367e-06, 1.011372e-06, 
    1.011369e-06, 1.011375e-06, 1.011373e-06, 1.011385e-06, 1.01139e-06, 
    1.011392e-06, 1.011393e-06, 1.011398e-06, 1.011395e-06, 1.011396e-06, 
    1.011393e-06, 1.011391e-06, 1.011392e-06, 1.011387e-06, 1.011389e-06, 
    1.011378e-06, 1.011383e-06, 1.011371e-06, 1.011374e-06, 1.01137e-06, 
    1.011372e-06, 1.011369e-06, 1.011372e-06, 1.011367e-06, 1.011366e-06, 
    1.011367e-06, 1.011364e-06, 1.011372e-06, 1.011369e-06, 1.011392e-06, 
    1.011392e-06, 1.011392e-06, 1.011394e-06, 1.011394e-06, 1.011397e-06, 
    1.011395e-06, 1.011394e-06, 1.011391e-06, 1.01139e-06, 1.011388e-06, 
    1.011385e-06, 1.011382e-06, 1.011377e-06, 1.011374e-06, 1.011371e-06, 
    1.011373e-06, 1.011372e-06, 1.011373e-06, 1.011374e-06, 1.011366e-06, 
    1.01137e-06, 1.011364e-06, 1.011365e-06, 1.011367e-06, 1.011365e-06, 
    1.011392e-06, 1.011393e-06, 1.011396e-06, 1.011393e-06, 1.011397e-06, 
    1.011395e-06, 1.011394e-06, 1.011389e-06, 1.011388e-06, 1.011387e-06, 
    1.011385e-06, 1.011382e-06, 1.011378e-06, 1.011374e-06, 1.011371e-06, 
    1.011371e-06, 1.011371e-06, 1.01137e-06, 1.011372e-06, 1.01137e-06, 
    1.011369e-06, 1.01137e-06, 1.011365e-06, 1.011366e-06, 1.011365e-06, 
    1.011366e-06, 1.011393e-06, 1.011391e-06, 1.011392e-06, 1.011391e-06, 
    1.011392e-06, 1.011387e-06, 1.011386e-06, 1.01138e-06, 1.011383e-06, 
    1.011379e-06, 1.011382e-06, 1.011382e-06, 1.011378e-06, 1.011382e-06, 
    1.011374e-06, 1.011379e-06, 1.01137e-06, 1.011375e-06, 1.01137e-06, 
    1.011371e-06, 1.011369e-06, 1.011368e-06, 1.011366e-06, 1.011362e-06, 
    1.011363e-06, 1.01136e-06, 1.011389e-06, 1.011388e-06, 1.011388e-06, 
    1.011386e-06, 1.011384e-06, 1.011382e-06, 1.011377e-06, 1.011379e-06, 
    1.011376e-06, 1.011375e-06, 1.01138e-06, 1.011377e-06, 1.011386e-06, 
    1.011385e-06, 1.011386e-06, 1.011389e-06, 1.011378e-06, 1.011384e-06, 
    1.011374e-06, 1.011377e-06, 1.011368e-06, 1.011372e-06, 1.011364e-06, 
    1.01136e-06, 1.011357e-06, 1.011353e-06, 1.011387e-06, 1.011388e-06, 
    1.011386e-06, 1.011383e-06, 1.01138e-06, 1.011376e-06, 1.011376e-06, 
    1.011375e-06, 1.011374e-06, 1.011372e-06, 1.011375e-06, 1.011372e-06, 
    1.011384e-06, 1.011378e-06, 1.011388e-06, 1.011385e-06, 1.011383e-06, 
    1.011384e-06, 1.011379e-06, 1.011378e-06, 1.011373e-06, 1.011375e-06, 
    1.011361e-06, 1.011367e-06, 1.01135e-06, 1.011354e-06, 1.011388e-06, 
    1.011387e-06, 1.011381e-06, 1.011384e-06, 1.011376e-06, 1.011374e-06, 
    1.011373e-06, 1.011371e-06, 1.011371e-06, 1.01137e-06, 1.011371e-06, 
    1.01137e-06, 1.011376e-06, 1.011373e-06, 1.011382e-06, 1.01138e-06, 
    1.011381e-06, 1.011382e-06, 1.011378e-06, 1.011375e-06, 1.011375e-06, 
    1.011374e-06, 1.011371e-06, 1.011376e-06, 1.01136e-06, 1.01137e-06, 
    1.011385e-06, 1.011382e-06, 1.011381e-06, 1.011383e-06, 1.011374e-06, 
    1.011377e-06, 1.01137e-06, 1.011372e-06, 1.011368e-06, 1.01137e-06, 
    1.01137e-06, 1.011372e-06, 1.011374e-06, 1.011377e-06, 1.01138e-06, 
    1.011382e-06, 1.011382e-06, 1.011379e-06, 1.011375e-06, 1.011371e-06, 
    1.011372e-06, 1.011369e-06, 1.011377e-06, 1.011373e-06, 1.011375e-06, 
    1.011371e-06, 1.011379e-06, 1.011372e-06, 1.01138e-06, 1.01138e-06, 
    1.011377e-06, 1.011373e-06, 1.011372e-06, 1.011371e-06, 1.011372e-06, 
    1.011375e-06, 1.011375e-06, 1.011378e-06, 1.011378e-06, 1.01138e-06, 
    1.011381e-06, 1.01138e-06, 1.011379e-06, 1.011375e-06, 1.011371e-06, 
    1.011368e-06, 1.011367e-06, 1.011362e-06, 1.011366e-06, 1.01136e-06, 
    1.011365e-06, 1.011356e-06, 1.011372e-06, 1.011365e-06, 1.011377e-06, 
    1.011376e-06, 1.011374e-06, 1.011368e-06, 1.011371e-06, 1.011368e-06, 
    1.011375e-06, 1.011379e-06, 1.01138e-06, 1.011382e-06, 1.01138e-06, 
    1.01138e-06, 1.011379e-06, 1.011379e-06, 1.011375e-06, 1.011377e-06, 
    1.01137e-06, 1.011368e-06, 1.011361e-06, 1.011356e-06, 1.011352e-06, 
    1.01135e-06, 1.01135e-06, 1.011349e-06 ;

 LITR1N_TNDNCY_VERT_TRANS =
  2.745014e-25, -4.901811e-26, -2.352869e-25, 2.352869e-25, -3.725376e-25, 
    1.764652e-25, -4.803775e-25, -6.078246e-25, 5.588064e-25, 7.352717e-25, 
    1.078398e-25, -5.686101e-25, -5.490028e-25, 2.058761e-25, 3.62734e-25, 
    -9.215405e-25, -1.56858e-25, -8.82326e-26, -1.470543e-25, -6.176282e-25, 
    -4.215557e-25, -1.274471e-25, 3.921449e-25, 1.176435e-25, 3.62734e-25, 
    6.764499e-25, 4.41163e-25, -1.666616e-25, -3.431268e-25, 3.333231e-25, 
    -1.960724e-26, -3.529304e-25, -3.235195e-25, 9.803622e-27, 1.019577e-24, 
    1.470543e-25, -3.921449e-25, 1.666616e-25, -1.176435e-25, 5.391992e-25, 
    1.372507e-25, 1.205845e-24, -1.56858e-25, -7.646825e-25, -4.41163e-25, 
    3.235195e-25, 1.088202e-24, 7.842898e-26, -1.862688e-25, 1.274471e-25, 
    9.803622e-27, -8.333079e-25, 2.254833e-25, -2.646978e-25, 9.901658e-25, 
    1.960724e-25, -3.235195e-25, 6.274318e-25, 3.235195e-25, -2.058761e-25, 
    2.941087e-25, -2.646978e-25, 5.391992e-25, 2.254833e-25, -2.058761e-25, 
    4.509666e-25, -4.215557e-25, 1.764652e-25, 7.450753e-25, -2.058761e-25, 
    -4.803775e-25, 3.235195e-25, -9.803622e-26, -1.372507e-25, 4.999847e-25, 
    5.19592e-25, 3.62734e-25, 3.823413e-25, -2.254833e-25, 5.588064e-25, 
    1.666616e-25, 2.843051e-25, -2.450906e-25, -2.941087e-26, -7.058608e-25, 
    2.941087e-25, 2.156797e-25, -1.470543e-25, 5.19592e-25, -8.235043e-25, 
    2.156797e-25, 6.078246e-25, -1.176435e-25, 7.646825e-25, -2.843051e-25, 
    3.62734e-25, 1.176435e-25, 3.431268e-25, 3.333231e-25, 3.235195e-25, 
    2.941087e-26, -2.058761e-25, -6.47039e-25, -8.82326e-26, 1.764652e-25, 
    7.842898e-26, 9.803622e-26, -4.41163e-25, 4.117521e-25, -2.450906e-25, 
    -2.745014e-25, -1.764652e-25, 3.039123e-25, -1.960724e-25, -3.725376e-25, 
    -5.097883e-25, -5.588064e-25, -5.882173e-26, 1.274471e-25, 4.019485e-25, 
    -2.352869e-25, 4.509666e-25, -5.882173e-25, -5.588064e-25, 6.960572e-25, 
    4.705739e-25, 3.333231e-25, 3.039123e-25, 2.352869e-25, -2.450906e-25, 
    -8.137007e-25, -4.705739e-25, 1.215649e-24, -3.62734e-25, 7.25468e-25, 
    2.745014e-25, 5.784137e-25, 1.274471e-25, -3.333231e-25, 1.470543e-25, 
    4.607703e-25, -3.921449e-25, -3.529304e-25, -2.450906e-25, 2.941087e-26, 
    -1.470543e-25, 5.98021e-25, 2.156797e-25, -3.039123e-25, 2.941087e-25, 
    9.901658e-25, -3.235195e-25, -2.352869e-25, -5.490028e-25, -3.039123e-25, 
    -7.450753e-25, 1.372507e-25, 4.019485e-25, -2.745014e-25, -6.862535e-26, 
    -1.176435e-25, 1.960724e-26, -7.940934e-25, -3.62734e-25, 8.82326e-25, 
    9.803622e-26, -6.372354e-25, 3.921449e-26, 3.725376e-25, -1.470543e-25, 
    4.901811e-26, 7.156644e-25, 1.372507e-25, -2.450906e-25, 2.450906e-25, 0, 
    1.764652e-25, -3.921449e-25, 1.215649e-24, -2.941087e-26, -7.058608e-25, 
    -1.764652e-25, 3.529304e-25, 4.215557e-25, 7.842898e-26, 7.058608e-25, 
    8.627187e-25, 4.509666e-25, 4.313593e-25, 1.372507e-25, -3.62734e-25, 
    2.548942e-25, -5.686101e-25, 4.117521e-25, -4.803775e-25, -3.529304e-25, 
    -7.744861e-25, -6.078246e-25, 1.862688e-25, 9.313441e-25, -2.058761e-25, 
    -1.666616e-25, 6.764499e-25, 6.078246e-25, -5.882173e-26, 2.058761e-25, 
    1.960724e-25, -7.156644e-25, -1.862688e-25, 3.62734e-25, 7.058608e-25, 
    2.646978e-25, -7.450753e-25, -5.784137e-25, -1.470543e-25, -1.960724e-26, 
    -2.745014e-25, -8.137007e-25, 3.235195e-25, 7.25468e-25, -7.842898e-26, 
    -1.960724e-25, 5.882173e-26, 4.509666e-25, 1.862688e-25, 2.646978e-25, 
    -6.176282e-25, 9.803622e-27, 4.117521e-25, 6.862535e-26, 8.529151e-25, 
    -2.058761e-25, -1.56858e-25, -7.744861e-25, -1.862688e-25, 2.450906e-25, 
    -7.744861e-25, -7.940934e-25, -4.705739e-25, -8.431115e-25, 
    -2.450906e-25, 1.862688e-25, 2.058761e-25, 4.803775e-25, -5.293956e-25, 
    -1.274471e-25, 2.058761e-25, -5.490028e-25, -1.960724e-25, -5.882173e-25, 
    -5.588064e-25, 4.901811e-25, 4.803775e-25, -7.058608e-25, 9.803622e-27, 
    -5.882173e-26, 1.470543e-25, -6.122413e-41, -3.431268e-25, -1.470543e-25, 
    0, -4.313593e-25, 1.274471e-25, -1.862688e-25, -2.254833e-25, 
    -2.843051e-25, -7.842898e-25, 1.274471e-25, -5.784137e-25, -6.274318e-25, 
    -2.941087e-26, 9.803622e-27, -8.137007e-25, -2.156797e-25, 7.744861e-25, 
    -3.431268e-25, -2.646978e-25, -1.372507e-25, -4.215557e-25, 
    -6.960572e-25, 4.313593e-25, 2.352869e-25, -1.764652e-25, -2.254833e-25, 
    3.235195e-25, 1.764652e-25, 3.921449e-26, -2.254833e-25, 1.372507e-25, 
    6.47039e-25, -6.47039e-25, 1.862688e-25, 1.274471e-25, 5.686101e-25, 
    4.999847e-25, -5.686101e-25, -5.097883e-25, 3.039123e-25, -6.176282e-25, 
    4.607703e-25, 7.842898e-26, -4.901811e-26, 2.548942e-25, -3.333231e-25, 
    6.862535e-26, 1.176435e-25, 4.607703e-25, 7.646825e-25, 1.56858e-25, 
    -3.333231e-25, -2.941087e-26, 7.058608e-25, 8.82326e-26, 5.588064e-25, 
    3.823413e-25, 5.882173e-26, 3.039123e-25, 1.196042e-24, -5.588064e-25, 
    6.47039e-25, -2.058761e-25, -6.960572e-25, -7.352717e-25, 6.862535e-26, 
    2.254833e-25, -7.646825e-25, 3.823413e-25, 4.215557e-25, -3.529304e-25, 
    -1.862688e-25, -3.725376e-25, 1.176435e-25, 9.803622e-27, -1.666616e-25, 
    3.725376e-25, 8.921296e-25, 9.803622e-26, -4.901811e-26,
  9.819577e-32, 9.819537e-32, 9.819544e-32, 9.819512e-32, 9.81953e-32, 
    9.819509e-32, 9.819568e-32, 9.819535e-32, 9.819557e-32, 9.819573e-32, 
    9.819449e-32, 9.81951e-32, 9.819385e-32, 9.819424e-32, 9.819326e-32, 
    9.819392e-32, 9.819313e-32, 9.819328e-32, 9.819283e-32, 9.819296e-32, 
    9.819238e-32, 9.819277e-32, 9.819208e-32, 9.819248e-32, 9.819241e-32, 
    9.819278e-32, 9.819498e-32, 9.819457e-32, 9.8195e-32, 9.819494e-32, 
    9.819497e-32, 9.81953e-32, 9.819546e-32, 9.81958e-32, 9.819574e-32, 
    9.819548e-32, 9.819492e-32, 9.819511e-32, 9.819463e-32, 9.819464e-32, 
    9.81941e-32, 9.819434e-32, 9.819344e-32, 9.819369e-32, 9.819295e-32, 
    9.819314e-32, 9.819296e-32, 9.819302e-32, 9.819296e-32, 9.819323e-32, 
    9.819312e-32, 9.819336e-32, 9.81943e-32, 9.819402e-32, 9.819484e-32, 
    9.819534e-32, 9.819567e-32, 9.819591e-32, 9.819587e-32, 9.819581e-32, 
    9.819548e-32, 9.819518e-32, 9.819495e-32, 9.819479e-32, 9.819464e-32, 
    9.819418e-32, 9.819393e-32, 9.819339e-32, 9.819349e-32, 9.819332e-32, 
    9.819316e-32, 9.819289e-32, 9.819293e-32, 9.819282e-32, 9.819332e-32, 
    9.819299e-32, 9.819354e-32, 9.819339e-32, 9.81946e-32, 9.819506e-32, 
    9.819526e-32, 9.819543e-32, 9.819585e-32, 9.819556e-32, 9.819567e-32, 
    9.81954e-32, 9.819523e-32, 9.819531e-32, 9.819479e-32, 9.819499e-32, 
    9.819392e-32, 9.819438e-32, 9.819317e-32, 9.819346e-32, 9.819311e-32, 
    9.819329e-32, 9.819298e-32, 9.819326e-32, 9.819278e-32, 9.819267e-32, 
    9.819274e-32, 9.819246e-32, 9.819327e-32, 9.819296e-32, 9.819531e-32, 
    9.81953e-32, 9.819524e-32, 9.819552e-32, 9.819554e-32, 9.81958e-32, 
    9.819557e-32, 9.819547e-32, 9.819522e-32, 9.819507e-32, 9.819493e-32, 
    9.819462e-32, 9.819427e-32, 9.819379e-32, 9.819345e-32, 9.819322e-32, 
    9.819336e-32, 9.819323e-32, 9.819337e-32, 9.819344e-32, 9.81927e-32, 
    9.819312e-32, 9.81925e-32, 9.819253e-32, 9.819282e-32, 9.819253e-32, 
    9.819529e-32, 9.819537e-32, 9.819565e-32, 9.819543e-32, 9.819583e-32, 
    9.819561e-32, 9.819548e-32, 9.819499e-32, 9.819488e-32, 9.819478e-32, 
    9.819459e-32, 9.819433e-32, 9.819389e-32, 9.81935e-32, 9.819315e-32, 
    9.819317e-32, 9.819316e-32, 9.819309e-32, 9.819328e-32, 9.819306e-32, 
    9.819302e-32, 9.819312e-32, 9.819254e-32, 9.81927e-32, 9.819253e-32, 
    9.819265e-32, 9.819534e-32, 9.819521e-32, 9.819528e-32, 9.819515e-32, 
    9.819524e-32, 9.819481e-32, 9.819469e-32, 9.819409e-32, 9.819433e-32, 
    9.819394e-32, 9.81943e-32, 9.819423e-32, 9.819393e-32, 9.819427e-32, 
    9.819352e-32, 9.819403e-32, 9.819309e-32, 9.819359e-32, 9.819305e-32, 
    9.819315e-32, 9.819299e-32, 9.819284e-32, 9.819266e-32, 9.819232e-32, 
    9.81924e-32, 9.819212e-32, 9.819501e-32, 9.819484e-32, 9.819485e-32, 
    9.819467e-32, 9.819453e-32, 9.819424e-32, 9.819377e-32, 9.819395e-32, 
    9.819363e-32, 9.819356e-32, 9.819406e-32, 9.819375e-32, 9.819472e-32, 
    9.819456e-32, 9.819466e-32, 9.8195e-32, 9.819391e-32, 9.819447e-32, 
    9.819344e-32, 9.819374e-32, 9.819286e-32, 9.81933e-32, 9.819244e-32, 
    9.819208e-32, 9.819174e-32, 9.819133e-32, 9.819474e-32, 9.819486e-32, 
    9.819465e-32, 9.819436e-32, 9.819409e-32, 9.819372e-32, 9.819369e-32, 
    9.819362e-32, 9.819345e-32, 9.81933e-32, 9.81936e-32, 9.819326e-32, 
    9.819453e-32, 9.819386e-32, 9.81949e-32, 9.819459e-32, 9.819437e-32, 
    9.819447e-32, 9.819397e-32, 9.819386e-32, 9.819338e-32, 9.819363e-32, 
    9.819216e-32, 9.819281e-32, 9.819102e-32, 9.819152e-32, 9.81949e-32, 
    9.819474e-32, 9.819419e-32, 9.819445e-32, 9.81937e-32, 9.819352e-32, 
    9.819336e-32, 9.819317e-32, 9.819315e-32, 9.819303e-32, 9.819322e-32, 
    9.819305e-32, 9.819372e-32, 9.819342e-32, 9.819425e-32, 9.819405e-32, 
    9.819414e-32, 9.819424e-32, 9.819393e-32, 9.819359e-32, 9.819359e-32, 
    9.819347e-32, 9.819317e-32, 9.81937e-32, 9.819208e-32, 9.819308e-32, 
    9.819457e-32, 9.819426e-32, 9.819422e-32, 9.819434e-32, 9.819353e-32, 
    9.819382e-32, 9.819304e-32, 9.819325e-32, 9.81929e-32, 9.819308e-32, 
    9.81931e-32, 9.819332e-32, 9.819346e-32, 9.819381e-32, 9.819409e-32, 
    9.819432e-32, 9.819427e-32, 9.819402e-32, 9.819357e-32, 9.819315e-32, 
    9.819324e-32, 9.819293e-32, 9.819375e-32, 9.819341e-32, 9.819354e-32, 
    9.819319e-32, 9.819396e-32, 9.81933e-32, 9.819412e-32, 9.819405e-32, 
    9.819383e-32, 9.819339e-32, 9.819329e-32, 9.819318e-32, 9.819325e-32, 
    9.819356e-32, 9.819361e-32, 9.819383e-32, 9.81939e-32, 9.819407e-32, 
    9.819421e-32, 9.819408e-32, 9.819394e-32, 9.819356e-32, 9.819322e-32, 
    9.819284e-32, 9.819275e-32, 9.819231e-32, 9.819266e-32, 9.819208e-32, 
    9.819258e-32, 9.819171e-32, 9.819327e-32, 9.819259e-32, 9.819382e-32, 
    9.819369e-32, 9.819345e-32, 9.81929e-32, 9.81932e-32, 9.819285e-32, 
    9.819362e-32, 9.819401e-32, 9.819412e-32, 9.81943e-32, 9.819411e-32, 
    9.819413e-32, 9.819394e-32, 9.8194e-32, 9.819355e-32, 9.819379e-32, 
    9.81931e-32, 9.819285e-32, 9.819215e-32, 9.819171e-32, 9.819128e-32, 
    9.819108e-32, 9.819102e-32, 9.8191e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N_TO_SOIL1N =
  4.240894e-14, 4.252371e-14, 4.250141e-14, 4.25939e-14, 4.254262e-14, 
    4.260315e-14, 4.243223e-14, 4.252825e-14, 4.246697e-14, 4.24193e-14, 
    4.27731e-14, 4.259802e-14, 4.295481e-14, 4.284335e-14, 4.312315e-14, 
    4.293745e-14, 4.316056e-14, 4.311783e-14, 4.324648e-14, 4.320965e-14, 
    4.337395e-14, 4.326348e-14, 4.345908e-14, 4.33476e-14, 4.336503e-14, 
    4.325983e-14, 4.263331e-14, 4.27513e-14, 4.262631e-14, 4.264315e-14, 
    4.26356e-14, 4.254366e-14, 4.249728e-14, 4.240019e-14, 4.241783e-14, 
    4.248915e-14, 4.265072e-14, 4.259592e-14, 4.273404e-14, 4.273092e-14, 
    4.288445e-14, 4.281526e-14, 4.307299e-14, 4.299982e-14, 4.321119e-14, 
    4.315806e-14, 4.320868e-14, 4.319334e-14, 4.320888e-14, 4.313096e-14, 
    4.316435e-14, 4.309577e-14, 4.282821e-14, 4.290691e-14, 4.267201e-14, 
    4.253046e-14, 4.243644e-14, 4.236965e-14, 4.237909e-14, 4.239709e-14, 
    4.248957e-14, 4.257648e-14, 4.264265e-14, 4.268689e-14, 4.273047e-14, 
    4.286217e-14, 4.29319e-14, 4.308776e-14, 4.305968e-14, 4.310728e-14, 
    4.315277e-14, 4.322907e-14, 4.321652e-14, 4.325012e-14, 4.310604e-14, 
    4.32018e-14, 4.304367e-14, 4.308694e-14, 4.274219e-14, 4.261071e-14, 
    4.255467e-14, 4.25057e-14, 4.238635e-14, 4.246878e-14, 4.243629e-14, 
    4.251359e-14, 4.256266e-14, 4.25384e-14, 4.26881e-14, 4.262992e-14, 
    4.293603e-14, 4.280428e-14, 4.314747e-14, 4.306545e-14, 4.316712e-14, 
    4.311526e-14, 4.32041e-14, 4.312414e-14, 4.326263e-14, 4.329274e-14, 
    4.327216e-14, 4.335124e-14, 4.311971e-14, 4.320867e-14, 4.253771e-14, 
    4.254167e-14, 4.256012e-14, 4.2479e-14, 4.247405e-14, 4.23997e-14, 
    4.246587e-14, 4.249402e-14, 4.256551e-14, 4.260776e-14, 4.264791e-14, 
    4.273613e-14, 4.283456e-14, 4.297208e-14, 4.307076e-14, 4.313687e-14, 
    4.309635e-14, 4.313212e-14, 4.309212e-14, 4.307338e-14, 4.328145e-14, 
    4.316465e-14, 4.333987e-14, 4.333019e-14, 4.325091e-14, 4.333128e-14, 
    4.254445e-14, 4.252167e-14, 4.244253e-14, 4.250447e-14, 4.23916e-14, 
    4.245478e-14, 4.249108e-14, 4.263111e-14, 4.266188e-14, 4.269037e-14, 
    4.274664e-14, 4.28188e-14, 4.294525e-14, 4.305516e-14, 4.315542e-14, 
    4.314809e-14, 4.315067e-14, 4.317304e-14, 4.311759e-14, 4.318214e-14, 
    4.319296e-14, 4.316465e-14, 4.332889e-14, 4.3282e-14, 4.332998e-14, 
    4.329946e-14, 4.252908e-14, 4.25674e-14, 4.25467e-14, 4.258562e-14, 
    4.255819e-14, 4.26801e-14, 4.271662e-14, 4.288739e-14, 4.281737e-14, 
    4.292882e-14, 4.282871e-14, 4.284645e-14, 4.29324e-14, 4.283413e-14, 
    4.304907e-14, 4.290335e-14, 4.317391e-14, 4.302851e-14, 4.318301e-14, 
    4.315499e-14, 4.32014e-14, 4.324293e-14, 4.329518e-14, 4.339148e-14, 
    4.336919e-14, 4.34497e-14, 4.262452e-14, 4.267417e-14, 4.266982e-14, 
    4.272178e-14, 4.276018e-14, 4.284339e-14, 4.29767e-14, 4.292659e-14, 
    4.301858e-14, 4.303701e-14, 4.289729e-14, 4.298309e-14, 4.27074e-14, 
    4.275197e-14, 4.272545e-14, 4.262842e-14, 4.293811e-14, 4.277928e-14, 
    4.307239e-14, 4.298651e-14, 4.3237e-14, 4.311247e-14, 4.335691e-14, 
    4.346118e-14, 4.355932e-14, 4.367376e-14, 4.270128e-14, 4.266756e-14, 
    4.272796e-14, 4.281143e-14, 4.288889e-14, 4.299175e-14, 4.300228e-14, 
    4.302153e-14, 4.307137e-14, 4.311328e-14, 4.302759e-14, 4.312378e-14, 
    4.276226e-14, 4.29519e-14, 4.265478e-14, 4.27443e-14, 4.280653e-14, 
    4.277926e-14, 4.292087e-14, 4.295421e-14, 4.308956e-14, 4.301964e-14, 
    4.343543e-14, 4.325166e-14, 4.376089e-14, 4.361883e-14, 4.265576e-14, 
    4.270118e-14, 4.285906e-14, 4.278397e-14, 4.299862e-14, 4.305136e-14, 
    4.309425e-14, 4.314901e-14, 4.315494e-14, 4.318738e-14, 4.313422e-14, 
    4.318529e-14, 4.299196e-14, 4.307839e-14, 4.284105e-14, 4.289886e-14, 
    4.287227e-14, 4.284309e-14, 4.293313e-14, 4.302893e-14, 4.303102e-14, 
    4.306169e-14, 4.314807e-14, 4.299949e-14, 4.345905e-14, 4.317539e-14, 
    4.275068e-14, 4.283801e-14, 4.285052e-14, 4.28167e-14, 4.304607e-14, 
    4.296303e-14, 4.318659e-14, 4.312622e-14, 4.322513e-14, 4.317599e-14, 
    4.316875e-14, 4.31056e-14, 4.306626e-14, 4.296683e-14, 4.288585e-14, 
    4.282161e-14, 4.283655e-14, 4.290711e-14, 4.30348e-14, 4.315546e-14, 
    4.312903e-14, 4.321762e-14, 4.298307e-14, 4.308145e-14, 4.304342e-14, 
    4.314257e-14, 4.292525e-14, 4.311022e-14, 4.287791e-14, 4.289831e-14, 
    4.296138e-14, 4.30881e-14, 4.311617e-14, 4.314608e-14, 4.312763e-14, 
    4.303802e-14, 4.302337e-14, 4.295985e-14, 4.294229e-14, 4.289387e-14, 
    4.285374e-14, 4.289039e-14, 4.292886e-14, 4.303808e-14, 4.31364e-14, 
    4.324351e-14, 4.326972e-14, 4.339461e-14, 4.32929e-14, 4.346062e-14, 
    4.331797e-14, 4.356483e-14, 4.312098e-14, 4.331385e-14, 4.296426e-14, 
    4.300199e-14, 4.307013e-14, 4.32264e-14, 4.31421e-14, 4.324069e-14, 
    4.30228e-14, 4.290952e-14, 4.288024e-14, 4.282551e-14, 4.288149e-14, 
    4.287694e-14, 4.293048e-14, 4.291328e-14, 4.30417e-14, 4.297275e-14, 
    4.316856e-14, 4.323992e-14, 4.344125e-14, 4.356445e-14, 4.368976e-14, 
    4.374502e-14, 4.376183e-14, 4.376886e-14 ;

 LITR1N_vr =
  5.77518e-05, 5.775157e-05, 5.775161e-05, 5.775143e-05, 5.775153e-05, 
    5.775141e-05, 5.775175e-05, 5.775156e-05, 5.775168e-05, 5.775178e-05, 
    5.775107e-05, 5.775142e-05, 5.775071e-05, 5.775093e-05, 5.775038e-05, 
    5.775075e-05, 5.77503e-05, 5.775039e-05, 5.775013e-05, 5.77502e-05, 
    5.774988e-05, 5.77501e-05, 5.774971e-05, 5.774993e-05, 5.774989e-05, 
    5.775011e-05, 5.775135e-05, 5.775112e-05, 5.775137e-05, 5.775133e-05, 
    5.775135e-05, 5.775153e-05, 5.775163e-05, 5.775182e-05, 5.775178e-05, 
    5.775164e-05, 5.775132e-05, 5.775143e-05, 5.775115e-05, 5.775116e-05, 
    5.775085e-05, 5.775099e-05, 5.775048e-05, 5.775062e-05, 5.77502e-05, 
    5.775031e-05, 5.775021e-05, 5.775024e-05, 5.775021e-05, 5.775036e-05, 
    5.775029e-05, 5.775043e-05, 5.775096e-05, 5.775081e-05, 5.775128e-05, 
    5.775156e-05, 5.775175e-05, 5.775188e-05, 5.775186e-05, 5.775183e-05, 
    5.775164e-05, 5.775147e-05, 5.775133e-05, 5.775125e-05, 5.775116e-05, 
    5.77509e-05, 5.775076e-05, 5.775045e-05, 5.77505e-05, 5.775041e-05, 
    5.775032e-05, 5.775017e-05, 5.775019e-05, 5.775012e-05, 5.775041e-05, 
    5.775022e-05, 5.775053e-05, 5.775045e-05, 5.775113e-05, 5.77514e-05, 
    5.775151e-05, 5.775161e-05, 5.775185e-05, 5.775168e-05, 5.775175e-05, 
    5.775159e-05, 5.775149e-05, 5.775154e-05, 5.775124e-05, 5.775136e-05, 
    5.775075e-05, 5.775101e-05, 5.775033e-05, 5.775049e-05, 5.775029e-05, 
    5.775039e-05, 5.775021e-05, 5.775037e-05, 5.77501e-05, 5.775004e-05, 
    5.775008e-05, 5.774992e-05, 5.775039e-05, 5.775021e-05, 5.775155e-05, 
    5.775153e-05, 5.77515e-05, 5.775166e-05, 5.775167e-05, 5.775182e-05, 
    5.775169e-05, 5.775163e-05, 5.775149e-05, 5.77514e-05, 5.775132e-05, 
    5.775115e-05, 5.775095e-05, 5.775068e-05, 5.775048e-05, 5.775035e-05, 
    5.775043e-05, 5.775036e-05, 5.775044e-05, 5.775048e-05, 5.775006e-05, 
    5.775029e-05, 5.774994e-05, 5.774996e-05, 5.775012e-05, 5.774996e-05, 
    5.775153e-05, 5.775157e-05, 5.775173e-05, 5.775161e-05, 5.775184e-05, 
    5.775171e-05, 5.775164e-05, 5.775136e-05, 5.775129e-05, 5.775124e-05, 
    5.775113e-05, 5.775098e-05, 5.775073e-05, 5.775051e-05, 5.775031e-05, 
    5.775033e-05, 5.775032e-05, 5.775028e-05, 5.775039e-05, 5.775026e-05, 
    5.775024e-05, 5.775029e-05, 5.774997e-05, 5.775006e-05, 5.774996e-05, 
    5.775003e-05, 5.775156e-05, 5.775148e-05, 5.775153e-05, 5.775145e-05, 
    5.77515e-05, 5.775126e-05, 5.775119e-05, 5.775085e-05, 5.775099e-05, 
    5.775076e-05, 5.775096e-05, 5.775093e-05, 5.775076e-05, 5.775095e-05, 
    5.775052e-05, 5.775081e-05, 5.775028e-05, 5.775056e-05, 5.775026e-05, 
    5.775031e-05, 5.775022e-05, 5.775014e-05, 5.775003e-05, 5.774984e-05, 
    5.774989e-05, 5.774973e-05, 5.775137e-05, 5.775127e-05, 5.775128e-05, 
    5.775118e-05, 5.77511e-05, 5.775093e-05, 5.775067e-05, 5.775077e-05, 
    5.775059e-05, 5.775055e-05, 5.775083e-05, 5.775065e-05, 5.775121e-05, 
    5.775112e-05, 5.775117e-05, 5.775136e-05, 5.775075e-05, 5.775106e-05, 
    5.775048e-05, 5.775065e-05, 5.775015e-05, 5.77504e-05, 5.774991e-05, 
    5.77497e-05, 5.774951e-05, 5.774928e-05, 5.775122e-05, 5.775128e-05, 
    5.775116e-05, 5.7751e-05, 5.775084e-05, 5.775064e-05, 5.775062e-05, 
    5.775058e-05, 5.775048e-05, 5.77504e-05, 5.775057e-05, 5.775037e-05, 
    5.775109e-05, 5.775072e-05, 5.775131e-05, 5.775113e-05, 5.775101e-05, 
    5.775106e-05, 5.775078e-05, 5.775071e-05, 5.775044e-05, 5.775058e-05, 
    5.774975e-05, 5.775012e-05, 5.77491e-05, 5.774939e-05, 5.775131e-05, 
    5.775122e-05, 5.77509e-05, 5.775105e-05, 5.775063e-05, 5.775052e-05, 
    5.775043e-05, 5.775032e-05, 5.775031e-05, 5.775025e-05, 5.775036e-05, 
    5.775025e-05, 5.775064e-05, 5.775047e-05, 5.775094e-05, 5.775083e-05, 
    5.775088e-05, 5.775093e-05, 5.775076e-05, 5.775056e-05, 5.775056e-05, 
    5.77505e-05, 5.775033e-05, 5.775062e-05, 5.77497e-05, 5.775027e-05, 
    5.775112e-05, 5.775095e-05, 5.775092e-05, 5.775099e-05, 5.775053e-05, 
    5.775069e-05, 5.775025e-05, 5.775037e-05, 5.775017e-05, 5.775027e-05, 
    5.775029e-05, 5.775041e-05, 5.775049e-05, 5.775069e-05, 5.775085e-05, 
    5.775098e-05, 5.775095e-05, 5.775081e-05, 5.775055e-05, 5.775031e-05, 
    5.775036e-05, 5.775019e-05, 5.775065e-05, 5.775046e-05, 5.775053e-05, 
    5.775034e-05, 5.775077e-05, 5.77504e-05, 5.775087e-05, 5.775083e-05, 
    5.77507e-05, 5.775045e-05, 5.775039e-05, 5.775033e-05, 5.775037e-05, 
    5.775055e-05, 5.775057e-05, 5.77507e-05, 5.775074e-05, 5.775083e-05, 
    5.775091e-05, 5.775084e-05, 5.775076e-05, 5.775055e-05, 5.775035e-05, 
    5.775014e-05, 5.775008e-05, 5.774984e-05, 5.775004e-05, 5.77497e-05, 
    5.774999e-05, 5.77495e-05, 5.775038e-05, 5.775e-05, 5.775069e-05, 
    5.775062e-05, 5.775048e-05, 5.775017e-05, 5.775034e-05, 5.775014e-05, 
    5.775058e-05, 5.77508e-05, 5.775086e-05, 5.775097e-05, 5.775086e-05, 
    5.775087e-05, 5.775076e-05, 5.77508e-05, 5.775054e-05, 5.775068e-05, 
    5.775029e-05, 5.775015e-05, 5.774974e-05, 5.77495e-05, 5.774925e-05, 
    5.774914e-05, 5.77491e-05, 5.774909e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1_HR =
  7.349627e-13, 7.369517e-13, 7.365653e-13, 7.38168e-13, 7.372793e-13, 
    7.383284e-13, 7.353664e-13, 7.370303e-13, 7.359684e-13, 7.351423e-13, 
    7.412737e-13, 7.382395e-13, 7.444228e-13, 7.424911e-13, 7.473402e-13, 
    7.441219e-13, 7.479886e-13, 7.472481e-13, 7.494776e-13, 7.488393e-13, 
    7.516866e-13, 7.497722e-13, 7.53162e-13, 7.5123e-13, 7.515321e-13, 
    7.497089e-13, 7.388511e-13, 7.40896e-13, 7.387298e-13, 7.390216e-13, 
    7.388908e-13, 7.372975e-13, 7.364937e-13, 7.34811e-13, 7.351168e-13, 
    7.363528e-13, 7.391528e-13, 7.382032e-13, 7.405967e-13, 7.405427e-13, 
    7.432035e-13, 7.420043e-13, 7.464709e-13, 7.452029e-13, 7.488659e-13, 
    7.479452e-13, 7.488226e-13, 7.485567e-13, 7.48826e-13, 7.474755e-13, 
    7.480542e-13, 7.468657e-13, 7.422289e-13, 7.435927e-13, 7.395217e-13, 
    7.370687e-13, 7.354393e-13, 7.342817e-13, 7.344454e-13, 7.347573e-13, 
    7.3636e-13, 7.378662e-13, 7.390131e-13, 7.397798e-13, 7.40535e-13, 
    7.428174e-13, 7.440257e-13, 7.46727e-13, 7.462402e-13, 7.470651e-13, 
    7.478536e-13, 7.491759e-13, 7.489584e-13, 7.495406e-13, 7.470438e-13, 
    7.487033e-13, 7.459628e-13, 7.467127e-13, 7.40738e-13, 7.384595e-13, 
    7.374884e-13, 7.366395e-13, 7.345712e-13, 7.359996e-13, 7.354366e-13, 
    7.367763e-13, 7.376267e-13, 7.372062e-13, 7.398007e-13, 7.387924e-13, 
    7.440973e-13, 7.418142e-13, 7.477617e-13, 7.463402e-13, 7.481023e-13, 
    7.472034e-13, 7.487431e-13, 7.473575e-13, 7.497574e-13, 7.502793e-13, 
    7.499226e-13, 7.512932e-13, 7.472805e-13, 7.488223e-13, 7.371944e-13, 
    7.37263e-13, 7.375826e-13, 7.361769e-13, 7.36091e-13, 7.348026e-13, 
    7.359493e-13, 7.364372e-13, 7.376762e-13, 7.384082e-13, 7.39104e-13, 
    7.406331e-13, 7.423389e-13, 7.447221e-13, 7.464323e-13, 7.475781e-13, 
    7.468757e-13, 7.474958e-13, 7.468025e-13, 7.464776e-13, 7.500836e-13, 
    7.480595e-13, 7.510961e-13, 7.509283e-13, 7.495543e-13, 7.509472e-13, 
    7.373111e-13, 7.369164e-13, 7.355448e-13, 7.366183e-13, 7.346622e-13, 
    7.357571e-13, 7.363862e-13, 7.38813e-13, 7.393463e-13, 7.3984e-13, 
    7.408152e-13, 7.420657e-13, 7.442572e-13, 7.461619e-13, 7.478996e-13, 
    7.477723e-13, 7.478171e-13, 7.482048e-13, 7.472439e-13, 7.483626e-13, 
    7.4855e-13, 7.480595e-13, 7.509058e-13, 7.500931e-13, 7.509247e-13, 
    7.503957e-13, 7.370448e-13, 7.377089e-13, 7.3735e-13, 7.380247e-13, 
    7.375492e-13, 7.39662e-13, 7.402949e-13, 7.432545e-13, 7.42041e-13, 
    7.439725e-13, 7.422374e-13, 7.425449e-13, 7.440345e-13, 7.423314e-13, 
    7.460564e-13, 7.435311e-13, 7.4822e-13, 7.457002e-13, 7.483777e-13, 
    7.47892e-13, 7.486962e-13, 7.49416e-13, 7.503215e-13, 7.519904e-13, 
    7.516042e-13, 7.529994e-13, 7.386988e-13, 7.395592e-13, 7.394839e-13, 
    7.403843e-13, 7.410498e-13, 7.42492e-13, 7.448021e-13, 7.439338e-13, 
    7.45528e-13, 7.458473e-13, 7.434259e-13, 7.449129e-13, 7.401352e-13, 
    7.409075e-13, 7.40448e-13, 7.387664e-13, 7.441334e-13, 7.413808e-13, 
    7.464605e-13, 7.449722e-13, 7.493134e-13, 7.471551e-13, 7.513914e-13, 
    7.531983e-13, 7.548992e-13, 7.568825e-13, 7.400291e-13, 7.394446e-13, 
    7.404914e-13, 7.419381e-13, 7.432804e-13, 7.45063e-13, 7.452454e-13, 
    7.455791e-13, 7.464429e-13, 7.471691e-13, 7.456841e-13, 7.473512e-13, 
    7.410857e-13, 7.443723e-13, 7.392232e-13, 7.407747e-13, 7.41853e-13, 
    7.413805e-13, 7.438347e-13, 7.444125e-13, 7.467581e-13, 7.455464e-13, 
    7.527522e-13, 7.495674e-13, 7.583925e-13, 7.559305e-13, 7.392402e-13, 
    7.400273e-13, 7.427634e-13, 7.414621e-13, 7.451821e-13, 7.460961e-13, 
    7.468393e-13, 7.477884e-13, 7.478912e-13, 7.484533e-13, 7.47532e-13, 
    7.484171e-13, 7.450667e-13, 7.465645e-13, 7.424513e-13, 7.434532e-13, 
    7.429925e-13, 7.424867e-13, 7.440471e-13, 7.457074e-13, 7.457435e-13, 
    7.462751e-13, 7.47772e-13, 7.451971e-13, 7.531616e-13, 7.482456e-13, 
    7.408851e-13, 7.423987e-13, 7.426155e-13, 7.420293e-13, 7.460044e-13, 
    7.445652e-13, 7.484397e-13, 7.473934e-13, 7.491076e-13, 7.482559e-13, 
    7.481306e-13, 7.470362e-13, 7.463544e-13, 7.446311e-13, 7.432277e-13, 
    7.421144e-13, 7.423734e-13, 7.435961e-13, 7.458091e-13, 7.479002e-13, 
    7.474421e-13, 7.489774e-13, 7.449126e-13, 7.466176e-13, 7.459584e-13, 
    7.476767e-13, 7.439106e-13, 7.471161e-13, 7.430901e-13, 7.434436e-13, 
    7.445366e-13, 7.467327e-13, 7.472193e-13, 7.477375e-13, 7.474179e-13, 
    7.458649e-13, 7.456111e-13, 7.445102e-13, 7.442059e-13, 7.433666e-13, 
    7.426713e-13, 7.433065e-13, 7.439731e-13, 7.458659e-13, 7.475699e-13, 
    7.494262e-13, 7.498804e-13, 7.520447e-13, 7.502821e-13, 7.531888e-13, 
    7.507165e-13, 7.549947e-13, 7.473027e-13, 7.506451e-13, 7.445866e-13, 
    7.452404e-13, 7.464214e-13, 7.491295e-13, 7.476686e-13, 7.493773e-13, 
    7.456012e-13, 7.43638e-13, 7.431305e-13, 7.42182e-13, 7.431522e-13, 
    7.430733e-13, 7.440012e-13, 7.437031e-13, 7.459287e-13, 7.447338e-13, 
    7.481272e-13, 7.493639e-13, 7.52853e-13, 7.54988e-13, 7.571598e-13, 
    7.581174e-13, 7.584088e-13, 7.585306e-13 ;

 LITR2C =
  2.015623e-05, 2.015621e-05, 2.015622e-05, 2.01562e-05, 2.015621e-05, 
    2.01562e-05, 2.015623e-05, 2.015621e-05, 2.015622e-05, 2.015623e-05, 
    2.015617e-05, 2.01562e-05, 2.015613e-05, 2.015615e-05, 2.01561e-05, 
    2.015614e-05, 2.015609e-05, 2.01561e-05, 2.015608e-05, 2.015609e-05, 
    2.015606e-05, 2.015608e-05, 2.015604e-05, 2.015606e-05, 2.015606e-05, 
    2.015608e-05, 2.015619e-05, 2.015617e-05, 2.015619e-05, 2.015619e-05, 
    2.015619e-05, 2.015621e-05, 2.015622e-05, 2.015623e-05, 2.015623e-05, 
    2.015622e-05, 2.015619e-05, 2.01562e-05, 2.015617e-05, 2.015617e-05, 
    2.015615e-05, 2.015616e-05, 2.015611e-05, 2.015612e-05, 2.015609e-05, 
    2.015609e-05, 2.015609e-05, 2.015609e-05, 2.015609e-05, 2.01561e-05, 
    2.015609e-05, 2.015611e-05, 2.015616e-05, 2.015614e-05, 2.015619e-05, 
    2.015621e-05, 2.015623e-05, 2.015624e-05, 2.015624e-05, 2.015623e-05, 
    2.015622e-05, 2.01562e-05, 2.015619e-05, 2.015618e-05, 2.015617e-05, 
    2.015615e-05, 2.015614e-05, 2.015611e-05, 2.015611e-05, 2.015611e-05, 
    2.01561e-05, 2.015608e-05, 2.015608e-05, 2.015608e-05, 2.015611e-05, 
    2.015609e-05, 2.015612e-05, 2.015611e-05, 2.015617e-05, 2.01562e-05, 
    2.015621e-05, 2.015621e-05, 2.015624e-05, 2.015622e-05, 2.015623e-05, 
    2.015621e-05, 2.015621e-05, 2.015621e-05, 2.015618e-05, 2.015619e-05, 
    2.015614e-05, 2.015616e-05, 2.01561e-05, 2.015611e-05, 2.015609e-05, 
    2.01561e-05, 2.015609e-05, 2.01561e-05, 2.015608e-05, 2.015607e-05, 
    2.015607e-05, 2.015606e-05, 2.01561e-05, 2.015609e-05, 2.015621e-05, 
    2.015621e-05, 2.015621e-05, 2.015622e-05, 2.015622e-05, 2.015623e-05, 
    2.015622e-05, 2.015622e-05, 2.01562e-05, 2.01562e-05, 2.015619e-05, 
    2.015617e-05, 2.015615e-05, 2.015613e-05, 2.015611e-05, 2.01561e-05, 
    2.015611e-05, 2.01561e-05, 2.015611e-05, 2.015611e-05, 2.015607e-05, 
    2.015609e-05, 2.015606e-05, 2.015606e-05, 2.015608e-05, 2.015606e-05, 
    2.015621e-05, 2.015621e-05, 2.015623e-05, 2.015622e-05, 2.015624e-05, 
    2.015623e-05, 2.015622e-05, 2.015619e-05, 2.015619e-05, 2.015618e-05, 
    2.015617e-05, 2.015616e-05, 2.015613e-05, 2.015611e-05, 2.01561e-05, 
    2.01561e-05, 2.01561e-05, 2.015609e-05, 2.01561e-05, 2.015609e-05, 
    2.015609e-05, 2.015609e-05, 2.015606e-05, 2.015607e-05, 2.015606e-05, 
    2.015607e-05, 2.015621e-05, 2.01562e-05, 2.015621e-05, 2.01562e-05, 
    2.015621e-05, 2.015618e-05, 2.015618e-05, 2.015615e-05, 2.015616e-05, 
    2.015614e-05, 2.015616e-05, 2.015615e-05, 2.015614e-05, 2.015615e-05, 
    2.015611e-05, 2.015614e-05, 2.015609e-05, 2.015612e-05, 2.015609e-05, 
    2.01561e-05, 2.015609e-05, 2.015608e-05, 2.015607e-05, 2.015605e-05, 
    2.015606e-05, 2.015604e-05, 2.015619e-05, 2.015618e-05, 2.015619e-05, 
    2.015618e-05, 2.015617e-05, 2.015615e-05, 2.015613e-05, 2.015614e-05, 
    2.015612e-05, 2.015612e-05, 2.015614e-05, 2.015613e-05, 2.015618e-05, 
    2.015617e-05, 2.015617e-05, 2.015619e-05, 2.015614e-05, 2.015617e-05, 
    2.015611e-05, 2.015613e-05, 2.015608e-05, 2.01561e-05, 2.015606e-05, 
    2.015604e-05, 2.015602e-05, 2.0156e-05, 2.015618e-05, 2.015619e-05, 
    2.015617e-05, 2.015616e-05, 2.015615e-05, 2.015613e-05, 2.015612e-05, 
    2.015612e-05, 2.015611e-05, 2.01561e-05, 2.015612e-05, 2.01561e-05, 
    2.015617e-05, 2.015613e-05, 2.015619e-05, 2.015617e-05, 2.015616e-05, 
    2.015617e-05, 2.015614e-05, 2.015613e-05, 2.015611e-05, 2.015612e-05, 
    2.015604e-05, 2.015608e-05, 2.015598e-05, 2.015601e-05, 2.015619e-05, 
    2.015618e-05, 2.015615e-05, 2.015616e-05, 2.015613e-05, 2.015611e-05, 
    2.015611e-05, 2.01561e-05, 2.01561e-05, 2.015609e-05, 2.01561e-05, 
    2.015609e-05, 2.015613e-05, 2.015611e-05, 2.015615e-05, 2.015614e-05, 
    2.015615e-05, 2.015615e-05, 2.015614e-05, 2.015612e-05, 2.015612e-05, 
    2.015611e-05, 2.01561e-05, 2.015612e-05, 2.015604e-05, 2.015609e-05, 
    2.015617e-05, 2.015615e-05, 2.015615e-05, 2.015616e-05, 2.015612e-05, 
    2.015613e-05, 2.015609e-05, 2.01561e-05, 2.015608e-05, 2.015609e-05, 
    2.015609e-05, 2.015611e-05, 2.015611e-05, 2.015613e-05, 2.015615e-05, 
    2.015616e-05, 2.015615e-05, 2.015614e-05, 2.015612e-05, 2.01561e-05, 
    2.01561e-05, 2.015608e-05, 2.015613e-05, 2.015611e-05, 2.015612e-05, 
    2.01561e-05, 2.015614e-05, 2.01561e-05, 2.015615e-05, 2.015614e-05, 
    2.015613e-05, 2.015611e-05, 2.01561e-05, 2.01561e-05, 2.01561e-05, 
    2.015612e-05, 2.015612e-05, 2.015613e-05, 2.015613e-05, 2.015614e-05, 
    2.015615e-05, 2.015614e-05, 2.015614e-05, 2.015612e-05, 2.01561e-05, 
    2.015608e-05, 2.015607e-05, 2.015605e-05, 2.015607e-05, 2.015604e-05, 
    2.015607e-05, 2.015602e-05, 2.01561e-05, 2.015607e-05, 2.015613e-05, 
    2.015612e-05, 2.015611e-05, 2.015608e-05, 2.01561e-05, 2.015608e-05, 
    2.015612e-05, 2.015614e-05, 2.015615e-05, 2.015616e-05, 2.015615e-05, 
    2.015615e-05, 2.015614e-05, 2.015614e-05, 2.015612e-05, 2.015613e-05, 
    2.015609e-05, 2.015608e-05, 2.015604e-05, 2.015602e-05, 2.0156e-05, 
    2.015599e-05, 2.015598e-05, 2.015598e-05 ;

 LITR2C_TO_SOIL1C =
  1.11921e-13, 1.122242e-13, 1.121653e-13, 1.124096e-13, 1.122741e-13, 
    1.12434e-13, 1.119825e-13, 1.122362e-13, 1.120743e-13, 1.119484e-13, 
    1.12883e-13, 1.124205e-13, 1.133631e-13, 1.130686e-13, 1.138078e-13, 
    1.133172e-13, 1.139066e-13, 1.137937e-13, 1.141336e-13, 1.140363e-13, 
    1.144703e-13, 1.141785e-13, 1.146953e-13, 1.144007e-13, 1.144468e-13, 
    1.141689e-13, 1.125137e-13, 1.128254e-13, 1.124952e-13, 1.125397e-13, 
    1.125198e-13, 1.122769e-13, 1.121544e-13, 1.118979e-13, 1.119445e-13, 
    1.121329e-13, 1.125597e-13, 1.12415e-13, 1.127798e-13, 1.127716e-13, 
    1.131772e-13, 1.129944e-13, 1.136753e-13, 1.13482e-13, 1.140404e-13, 
    1.139e-13, 1.140338e-13, 1.139932e-13, 1.140343e-13, 1.138284e-13, 
    1.139166e-13, 1.137354e-13, 1.130286e-13, 1.132365e-13, 1.12616e-13, 
    1.12242e-13, 1.119936e-13, 1.118172e-13, 1.118421e-13, 1.118897e-13, 
    1.12134e-13, 1.123636e-13, 1.125384e-13, 1.126553e-13, 1.127704e-13, 
    1.131183e-13, 1.133025e-13, 1.137143e-13, 1.136401e-13, 1.137658e-13, 
    1.13886e-13, 1.140876e-13, 1.140545e-13, 1.141432e-13, 1.137626e-13, 
    1.140156e-13, 1.135978e-13, 1.137121e-13, 1.128014e-13, 1.12454e-13, 
    1.12306e-13, 1.121766e-13, 1.118613e-13, 1.120791e-13, 1.119932e-13, 
    1.121974e-13, 1.123271e-13, 1.12263e-13, 1.126585e-13, 1.125048e-13, 
    1.133134e-13, 1.129654e-13, 1.13872e-13, 1.136553e-13, 1.13924e-13, 
    1.137869e-13, 1.140216e-13, 1.138104e-13, 1.141763e-13, 1.142558e-13, 
    1.142014e-13, 1.144104e-13, 1.137987e-13, 1.140337e-13, 1.122612e-13, 
    1.122716e-13, 1.123204e-13, 1.121061e-13, 1.12093e-13, 1.118966e-13, 
    1.120714e-13, 1.121458e-13, 1.123346e-13, 1.124462e-13, 1.125523e-13, 
    1.127854e-13, 1.130454e-13, 1.134087e-13, 1.136694e-13, 1.13844e-13, 
    1.13737e-13, 1.138315e-13, 1.137258e-13, 1.136763e-13, 1.14226e-13, 
    1.139174e-13, 1.143803e-13, 1.143547e-13, 1.141453e-13, 1.143576e-13, 
    1.12279e-13, 1.122188e-13, 1.120097e-13, 1.121734e-13, 1.118752e-13, 
    1.120421e-13, 1.12138e-13, 1.125079e-13, 1.125892e-13, 1.126645e-13, 
    1.128131e-13, 1.130037e-13, 1.133378e-13, 1.136282e-13, 1.138931e-13, 
    1.138737e-13, 1.138805e-13, 1.139396e-13, 1.137931e-13, 1.139636e-13, 
    1.139922e-13, 1.139174e-13, 1.143513e-13, 1.142274e-13, 1.143542e-13, 
    1.142736e-13, 1.122384e-13, 1.123396e-13, 1.122849e-13, 1.123878e-13, 
    1.123153e-13, 1.126373e-13, 1.127338e-13, 1.13185e-13, 1.13e-13, 
    1.132944e-13, 1.130299e-13, 1.130768e-13, 1.133039e-13, 1.130442e-13, 
    1.136121e-13, 1.132271e-13, 1.139419e-13, 1.135578e-13, 1.139659e-13, 
    1.138919e-13, 1.140145e-13, 1.141242e-13, 1.142623e-13, 1.145167e-13, 
    1.144578e-13, 1.146705e-13, 1.124905e-13, 1.126217e-13, 1.126102e-13, 
    1.127474e-13, 1.128489e-13, 1.130687e-13, 1.134209e-13, 1.132885e-13, 
    1.135315e-13, 1.135802e-13, 1.132111e-13, 1.134378e-13, 1.127095e-13, 
    1.128272e-13, 1.127572e-13, 1.125008e-13, 1.133189e-13, 1.128993e-13, 
    1.136737e-13, 1.134468e-13, 1.141086e-13, 1.137796e-13, 1.144254e-13, 
    1.147008e-13, 1.149601e-13, 1.152624e-13, 1.126933e-13, 1.126042e-13, 
    1.127638e-13, 1.129843e-13, 1.131889e-13, 1.134606e-13, 1.134885e-13, 
    1.135393e-13, 1.13671e-13, 1.137817e-13, 1.135553e-13, 1.138095e-13, 
    1.128544e-13, 1.133554e-13, 1.125704e-13, 1.128069e-13, 1.129713e-13, 
    1.128993e-13, 1.132734e-13, 1.133615e-13, 1.137191e-13, 1.135343e-13, 
    1.146328e-13, 1.141473e-13, 1.154926e-13, 1.151173e-13, 1.12573e-13, 
    1.12693e-13, 1.131101e-13, 1.129117e-13, 1.134788e-13, 1.136181e-13, 
    1.137314e-13, 1.138761e-13, 1.138918e-13, 1.139775e-13, 1.13837e-13, 
    1.139719e-13, 1.134612e-13, 1.136895e-13, 1.130625e-13, 1.132152e-13, 
    1.13145e-13, 1.130679e-13, 1.133058e-13, 1.135589e-13, 1.135644e-13, 
    1.136454e-13, 1.138736e-13, 1.134811e-13, 1.146952e-13, 1.139458e-13, 
    1.128238e-13, 1.130545e-13, 1.130876e-13, 1.129982e-13, 1.136041e-13, 
    1.133848e-13, 1.139754e-13, 1.138159e-13, 1.140772e-13, 1.139474e-13, 
    1.139283e-13, 1.137614e-13, 1.136575e-13, 1.133948e-13, 1.131809e-13, 
    1.130112e-13, 1.130506e-13, 1.13237e-13, 1.135744e-13, 1.138931e-13, 
    1.138233e-13, 1.140574e-13, 1.134377e-13, 1.136976e-13, 1.135971e-13, 
    1.138591e-13, 1.13285e-13, 1.137736e-13, 1.131599e-13, 1.132138e-13, 
    1.133804e-13, 1.137152e-13, 1.137893e-13, 1.138683e-13, 1.138196e-13, 
    1.135829e-13, 1.135442e-13, 1.133764e-13, 1.1333e-13, 1.132021e-13, 
    1.130961e-13, 1.131929e-13, 1.132945e-13, 1.13583e-13, 1.138428e-13, 
    1.141258e-13, 1.14195e-13, 1.145249e-13, 1.142562e-13, 1.146993e-13, 
    1.143225e-13, 1.149746e-13, 1.138021e-13, 1.143116e-13, 1.13388e-13, 
    1.134877e-13, 1.136677e-13, 1.140805e-13, 1.138579e-13, 1.141183e-13, 
    1.135427e-13, 1.132434e-13, 1.131661e-13, 1.130215e-13, 1.131694e-13, 
    1.131573e-13, 1.132988e-13, 1.132534e-13, 1.135926e-13, 1.134105e-13, 
    1.139277e-13, 1.141163e-13, 1.146481e-13, 1.149736e-13, 1.153047e-13, 
    1.154507e-13, 1.154951e-13, 1.155137e-13 ;

 LITR2C_vr =
  0.001150942, 0.001150941, 0.001150941, 0.00115094, 0.00115094, 0.00115094, 
    0.001150941, 0.00115094, 0.001150941, 0.001150942, 0.001150938, 
    0.00115094, 0.001150936, 0.001150937, 0.001150934, 0.001150936, 
    0.001150934, 0.001150934, 0.001150933, 0.001150933, 0.001150932, 
    0.001150933, 0.001150931, 0.001150932, 0.001150932, 0.001150933, 
    0.001150939, 0.001150938, 0.001150939, 0.001150939, 0.001150939, 
    0.00115094, 0.001150941, 0.001150942, 0.001150942, 0.001150941, 
    0.001150939, 0.00115094, 0.001150938, 0.001150938, 0.001150937, 
    0.001150937, 0.001150935, 0.001150936, 0.001150933, 0.001150934, 
    0.001150933, 0.001150933, 0.001150933, 0.001150934, 0.001150934, 
    0.001150934, 0.001150937, 0.001150936, 0.001150939, 0.00115094, 
    0.001150941, 0.001150942, 0.001150942, 0.001150942, 0.001150941, 
    0.00115094, 0.001150939, 0.001150939, 0.001150938, 0.001150937, 
    0.001150936, 0.001150935, 0.001150935, 0.001150934, 0.001150934, 
    0.001150933, 0.001150933, 0.001150933, 0.001150934, 0.001150933, 
    0.001150935, 0.001150935, 0.001150938, 0.00115094, 0.00115094, 
    0.001150941, 0.001150942, 0.001150941, 0.001150941, 0.001150941, 
    0.00115094, 0.00115094, 0.001150939, 0.001150939, 0.001150936, 
    0.001150938, 0.001150934, 0.001150935, 0.001150934, 0.001150934, 
    0.001150933, 0.001150934, 0.001150933, 0.001150932, 0.001150933, 
    0.001150932, 0.001150934, 0.001150933, 0.00115094, 0.00115094, 
    0.00115094, 0.001150941, 0.001150941, 0.001150942, 0.001150941, 
    0.001150941, 0.00115094, 0.00115094, 0.001150939, 0.001150938, 
    0.001150937, 0.001150936, 0.001150935, 0.001150934, 0.001150934, 
    0.001150934, 0.001150934, 0.001150935, 0.001150933, 0.001150934, 
    0.001150932, 0.001150932, 0.001150933, 0.001150932, 0.00115094, 
    0.001150941, 0.001150941, 0.001150941, 0.001150942, 0.001150941, 
    0.001150941, 0.001150939, 0.001150939, 0.001150939, 0.001150938, 
    0.001150937, 0.001150936, 0.001150935, 0.001150934, 0.001150934, 
    0.001150934, 0.001150934, 0.001150934, 0.001150934, 0.001150933, 
    0.001150934, 0.001150932, 0.001150933, 0.001150932, 0.001150932, 
    0.00115094, 0.00115094, 0.00115094, 0.00115094, 0.00115094, 0.001150939, 
    0.001150938, 0.001150937, 0.001150937, 0.001150936, 0.001150937, 
    0.001150937, 0.001150936, 0.001150937, 0.001150935, 0.001150936, 
    0.001150934, 0.001150935, 0.001150934, 0.001150934, 0.001150933, 
    0.001150933, 0.001150932, 0.001150931, 0.001150932, 0.001150931, 
    0.001150939, 0.001150939, 0.001150939, 0.001150938, 0.001150938, 
    0.001150937, 0.001150936, 0.001150936, 0.001150935, 0.001150935, 
    0.001150937, 0.001150936, 0.001150939, 0.001150938, 0.001150938, 
    0.001150939, 0.001150936, 0.001150938, 0.001150935, 0.001150936, 
    0.001150933, 0.001150934, 0.001150932, 0.001150931, 0.00115093, 
    0.001150928, 0.001150939, 0.001150939, 0.001150938, 0.001150938, 
    0.001150937, 0.001150936, 0.001150936, 0.001150935, 0.001150935, 
    0.001150934, 0.001150935, 0.001150934, 0.001150938, 0.001150936, 
    0.001150939, 0.001150938, 0.001150938, 0.001150938, 0.001150936, 
    0.001150936, 0.001150935, 0.001150935, 0.001150931, 0.001150933, 
    0.001150928, 0.001150929, 0.001150939, 0.001150939, 0.001150937, 
    0.001150938, 0.001150936, 0.001150935, 0.001150934, 0.001150934, 
    0.001150934, 0.001150934, 0.001150934, 0.001150934, 0.001150936, 
    0.001150935, 0.001150937, 0.001150937, 0.001150937, 0.001150937, 
    0.001150936, 0.001150935, 0.001150935, 0.001150935, 0.001150934, 
    0.001150936, 0.001150931, 0.001150934, 0.001150938, 0.001150937, 
    0.001150937, 0.001150937, 0.001150935, 0.001150936, 0.001150934, 
    0.001150934, 0.001150933, 0.001150934, 0.001150934, 0.001150934, 
    0.001150935, 0.001150936, 0.001150937, 0.001150937, 0.001150937, 
    0.001150936, 0.001150935, 0.001150934, 0.001150934, 0.001150933, 
    0.001150936, 0.001150935, 0.001150935, 0.001150934, 0.001150936, 
    0.001150934, 0.001150937, 0.001150937, 0.001150936, 0.001150935, 
    0.001150934, 0.001150934, 0.001150934, 0.001150935, 0.001150935, 
    0.001150936, 0.001150936, 0.001150937, 0.001150937, 0.001150937, 
    0.001150936, 0.001150935, 0.001150934, 0.001150933, 0.001150933, 
    0.001150931, 0.001150932, 0.001150931, 0.001150932, 0.00115093, 
    0.001150934, 0.001150932, 0.001150936, 0.001150936, 0.001150935, 
    0.001150933, 0.001150934, 0.001150933, 0.001150935, 0.001150936, 
    0.001150937, 0.001150937, 0.001150937, 0.001150937, 0.001150936, 
    0.001150936, 0.001150935, 0.001150936, 0.001150934, 0.001150933, 
    0.001150931, 0.00115093, 0.001150928, 0.001150928, 0.001150928, 
    0.001150927,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N =
  2.789474e-07, 2.789471e-07, 2.789472e-07, 2.78947e-07, 2.789471e-07, 
    2.789469e-07, 2.789474e-07, 2.789471e-07, 2.789473e-07, 2.789474e-07, 
    2.789465e-07, 2.789469e-07, 2.78946e-07, 2.789463e-07, 2.789456e-07, 
    2.789461e-07, 2.789455e-07, 2.789456e-07, 2.789453e-07, 2.789454e-07, 
    2.78945e-07, 2.789453e-07, 2.789448e-07, 2.78945e-07, 2.78945e-07, 
    2.789453e-07, 2.789469e-07, 2.789466e-07, 2.789469e-07, 2.789468e-07, 
    2.789469e-07, 2.789471e-07, 2.789472e-07, 2.789475e-07, 2.789474e-07, 
    2.789472e-07, 2.789468e-07, 2.78947e-07, 2.789466e-07, 2.789466e-07, 
    2.789462e-07, 2.789464e-07, 2.789457e-07, 2.789459e-07, 2.789454e-07, 
    2.789455e-07, 2.789454e-07, 2.789454e-07, 2.789454e-07, 2.789456e-07, 
    2.789455e-07, 2.789457e-07, 2.789464e-07, 2.789462e-07, 2.789468e-07, 
    2.789471e-07, 2.789474e-07, 2.789475e-07, 2.789475e-07, 2.789475e-07, 
    2.789472e-07, 2.78947e-07, 2.789468e-07, 2.789467e-07, 2.789466e-07, 
    2.789463e-07, 2.789461e-07, 2.789457e-07, 2.789458e-07, 2.789457e-07, 
    2.789455e-07, 2.789454e-07, 2.789454e-07, 2.789453e-07, 2.789457e-07, 
    2.789454e-07, 2.789458e-07, 2.789457e-07, 2.789466e-07, 2.789469e-07, 
    2.789471e-07, 2.789472e-07, 2.789475e-07, 2.789473e-07, 2.789474e-07, 
    2.789472e-07, 2.789471e-07, 2.789471e-07, 2.789467e-07, 2.789469e-07, 
    2.789461e-07, 2.789464e-07, 2.789455e-07, 2.789457e-07, 2.789455e-07, 
    2.789456e-07, 2.789454e-07, 2.789456e-07, 2.789453e-07, 2.789452e-07, 
    2.789452e-07, 2.78945e-07, 2.789456e-07, 2.789454e-07, 2.789471e-07, 
    2.789471e-07, 2.789471e-07, 2.789473e-07, 2.789473e-07, 2.789475e-07, 
    2.789473e-07, 2.789472e-07, 2.78947e-07, 2.789469e-07, 2.789468e-07, 
    2.789466e-07, 2.789463e-07, 2.78946e-07, 2.789457e-07, 2.789456e-07, 
    2.789457e-07, 2.789456e-07, 2.789457e-07, 2.789457e-07, 2.789452e-07, 
    2.789455e-07, 2.789451e-07, 2.789451e-07, 2.789453e-07, 2.789451e-07, 
    2.789471e-07, 2.789471e-07, 2.789473e-07, 2.789472e-07, 2.789475e-07, 
    2.789473e-07, 2.789472e-07, 2.789469e-07, 2.789468e-07, 2.789467e-07, 
    2.789466e-07, 2.789464e-07, 2.789461e-07, 2.789458e-07, 2.789455e-07, 
    2.789455e-07, 2.789455e-07, 2.789455e-07, 2.789456e-07, 2.789455e-07, 
    2.789454e-07, 2.789455e-07, 2.789451e-07, 2.789452e-07, 2.789451e-07, 
    2.789452e-07, 2.789471e-07, 2.78947e-07, 2.789471e-07, 2.78947e-07, 
    2.789471e-07, 2.789467e-07, 2.789467e-07, 2.789462e-07, 2.789464e-07, 
    2.789461e-07, 2.789464e-07, 2.789463e-07, 2.789461e-07, 2.789463e-07, 
    2.789458e-07, 2.789462e-07, 2.789455e-07, 2.789459e-07, 2.789455e-07, 
    2.789455e-07, 2.789454e-07, 2.789453e-07, 2.789452e-07, 2.789449e-07, 
    2.78945e-07, 2.789448e-07, 2.789469e-07, 2.789468e-07, 2.789468e-07, 
    2.789466e-07, 2.789465e-07, 2.789463e-07, 2.78946e-07, 2.789461e-07, 
    2.789459e-07, 2.789458e-07, 2.789462e-07, 2.78946e-07, 2.789467e-07, 
    2.789466e-07, 2.789466e-07, 2.789469e-07, 2.789461e-07, 2.789465e-07, 
    2.789457e-07, 2.789459e-07, 2.789453e-07, 2.789456e-07, 2.78945e-07, 
    2.789448e-07, 2.789445e-07, 2.789442e-07, 2.789467e-07, 2.789468e-07, 
    2.789466e-07, 2.789464e-07, 2.789462e-07, 2.789459e-07, 2.789459e-07, 
    2.789459e-07, 2.789457e-07, 2.789456e-07, 2.789459e-07, 2.789456e-07, 
    2.789465e-07, 2.789461e-07, 2.789468e-07, 2.789466e-07, 2.789464e-07, 
    2.789465e-07, 2.789461e-07, 2.78946e-07, 2.789457e-07, 2.789459e-07, 
    2.789448e-07, 2.789453e-07, 2.78944e-07, 2.789444e-07, 2.789468e-07, 
    2.789467e-07, 2.789463e-07, 2.789465e-07, 2.789459e-07, 2.789458e-07, 
    2.789457e-07, 2.789455e-07, 2.789455e-07, 2.789454e-07, 2.789456e-07, 
    2.789455e-07, 2.789459e-07, 2.789457e-07, 2.789463e-07, 2.789462e-07, 
    2.789463e-07, 2.789463e-07, 2.789461e-07, 2.789459e-07, 2.789458e-07, 
    2.789458e-07, 2.789455e-07, 2.789459e-07, 2.789448e-07, 2.789455e-07, 
    2.789466e-07, 2.789463e-07, 2.789463e-07, 2.789464e-07, 2.789458e-07, 
    2.78946e-07, 2.789454e-07, 2.789456e-07, 2.789454e-07, 2.789455e-07, 
    2.789455e-07, 2.789457e-07, 2.789457e-07, 2.78946e-07, 2.789462e-07, 
    2.789464e-07, 2.789463e-07, 2.789462e-07, 2.789458e-07, 2.789455e-07, 
    2.789456e-07, 2.789454e-07, 2.78946e-07, 2.789457e-07, 2.789458e-07, 
    2.789455e-07, 2.789461e-07, 2.789456e-07, 2.789462e-07, 2.789462e-07, 
    2.78946e-07, 2.789457e-07, 2.789456e-07, 2.789455e-07, 2.789456e-07, 
    2.789458e-07, 2.789459e-07, 2.78946e-07, 2.789461e-07, 2.789462e-07, 
    2.789463e-07, 2.789462e-07, 2.789461e-07, 2.789458e-07, 2.789456e-07, 
    2.789453e-07, 2.789452e-07, 2.789449e-07, 2.789452e-07, 2.789448e-07, 
    2.789451e-07, 2.789445e-07, 2.789456e-07, 2.789451e-07, 2.78946e-07, 
    2.789459e-07, 2.789457e-07, 2.789454e-07, 2.789455e-07, 2.789453e-07, 
    2.789459e-07, 2.789461e-07, 2.789462e-07, 2.789464e-07, 2.789462e-07, 
    2.789462e-07, 2.789461e-07, 2.789461e-07, 2.789458e-07, 2.78946e-07, 
    2.789455e-07, 2.789453e-07, 2.789448e-07, 2.789445e-07, 2.789442e-07, 
    2.78944e-07, 2.78944e-07, 2.78944e-07 ;

 LITR2N_TNDNCY_VERT_TRANS =
  1.323489e-25, 1.225453e-26, -2.205815e-25, -6.862535e-26, -1.470543e-26, 
    5.637083e-26, 1.642107e-25, 9.803622e-27, 7.107626e-26, -4.65672e-26, 
    1.985233e-25, 8.82326e-26, -2.941087e-26, 2.941087e-26, 1.127417e-25, 
    1.225453e-26, -7.352717e-27, 3.431268e-26, -1.102908e-25, -1.102908e-25, 
    5.882173e-26, -6.372354e-26, 1.617598e-25, 1.372507e-25, -1.274471e-25, 
    1.274471e-25, 1.102908e-25, -1.960724e-26, -4.901811e-26, -9.803622e-27, 
    1.127417e-25, 7.107626e-26, 1.200944e-25, 2.695996e-26, 4.41163e-26, 
    -2.695996e-25, -3.431268e-26, -9.803622e-26, -2.009742e-25, 
    -1.249962e-25, -1.862688e-25, -1.02938e-25, 4.901811e-27, 8.82326e-26, 
    -2.695996e-26, -2.401887e-25, -2.646978e-25, -1.225453e-25, 3.186177e-26, 
    6.862535e-26, 1.397016e-25, 2.009742e-25, -1.642107e-25, -3.921449e-26, 
    -3.38225e-25, 2.695996e-26, 2.671487e-25, -7.842898e-26, 1.151926e-25, 
    7.352717e-27, 4.65672e-26, -9.313441e-26, 6.372354e-26, -6.617445e-26, 
    6.862535e-26, -9.313441e-26, -1.004871e-25, -3.774394e-25, 8.578169e-26, 
    2.205815e-25, -3.357741e-25, 8.087988e-26, -2.450905e-26, 1.323489e-25, 
    -1.347998e-25, 9.558531e-26, -1.200944e-25, -6.862535e-26, -1.249962e-25, 
    -1.960724e-26, -9.068351e-26, 1.02938e-25, -4.65672e-26, -4.41163e-26, 
    1.02938e-25, 9.558531e-26, 1.225453e-26, 2.695996e-26, 1.911706e-25, 
    -2.254833e-25, -9.313441e-26, -1.691125e-25, -7.107626e-26, 2.254833e-25, 
    1.176435e-25, -9.313441e-26, 1.862688e-25, 4.41163e-26, 2.573451e-25, 
    8.333079e-26, 1.323489e-25, 2.377378e-25, 1.200944e-25, -9.558531e-26, 
    -5.146902e-26, 2.034252e-25, -1.985233e-25, 1.053889e-25, -1.715634e-26, 
    -2.695996e-26, 1.960724e-26, -1.347998e-25, 4.901811e-27, 4.901811e-27, 
    1.81367e-25, 1.617598e-25, 7.352717e-26, 2.941087e-26, -9.068351e-26, 
    1.715634e-25, 1.274471e-25, 1.323489e-25, 9.313441e-26, -1.715634e-26, 
    1.740143e-25, -3.186177e-26, -3.431268e-26, -2.916578e-25, -1.176435e-25, 
    4.901811e-26, -1.838179e-25, -6.862535e-26, -1.56858e-25, 5.391992e-26, 
    -2.843051e-25, -2.867559e-25, 2.695996e-26, -7.597807e-26, 2.205815e-26, 
    -2.205815e-26, 0, 1.960724e-26, 1.372507e-25, 2.205815e-25, 4.901811e-26, 
    1.446034e-25, 4.41163e-26, -3.970467e-25, 1.740143e-25, -2.401887e-25, 
    1.053889e-25, 1.691125e-25, 9.803622e-26, 1.02938e-25, 2.450906e-25, 
    -2.450906e-27, -3.431268e-26, 2.058761e-25, -5.146902e-26, 6.862535e-26, 
    9.558531e-26, -4.901811e-26, 6.862535e-26, -3.431268e-25, -1.274471e-25, 
    3.749886e-25, 7.352717e-27, -1.02938e-25, -1.56858e-25, 1.495052e-25, 
    -3.088141e-25, 8.333079e-26, -7.842898e-26, -2.695996e-26, 6.127264e-26, 
    8.333079e-26, 6.862535e-26, -1.862688e-25, -3.921449e-26, 2.230324e-25, 
    7.597807e-26, 1.053889e-25, 4.901811e-27, 1.470543e-26, 1.29898e-25, 
    -5.637083e-26, -6.862535e-26, -1.078398e-25, -3.186177e-26, 3.553813e-25, 
    -5.637083e-26, 3.186177e-26, -4.901811e-26, -5.637083e-26, 5.637083e-26, 
    -1.446034e-25, 2.695996e-26, -3.235195e-25, 1.249962e-25, -1.960724e-26, 
    2.181306e-25, -4.901811e-27, -7.842898e-26, 3.725376e-25, -1.347998e-25, 
    1.470543e-26, -6.372354e-26, -6.617445e-26, -1.225453e-26, -1.519561e-25, 
    -1.249962e-25, -8.087988e-26, 4.019485e-25, -1.078398e-25, 1.691125e-25, 
    -8.087988e-26, -3.676358e-26, -1.225453e-25, -1.053889e-25, 
    -3.186177e-26, 9.313441e-26, 5.146902e-26, -1.911706e-25, 2.303851e-25, 
    6.127264e-26, 1.81367e-25, -1.960724e-26, 1.691125e-25, 3.431268e-26, 
    6.617445e-26, 7.352717e-27, -2.450905e-26, 2.205815e-26, 1.004871e-25, 
    -7.352717e-27, 4.901811e-27, 6.127264e-26, -1.372507e-25, 1.02938e-25, 
    4.901811e-27, -4.901811e-26, -3.357741e-25, -4.901811e-26, 1.397016e-25, 
    1.225453e-25, 1.470543e-26, 1.593089e-25, -1.838179e-25, 2.303851e-25, 
    8.82326e-26, -2.59796e-25, 9.558531e-26, 2.401887e-25, -4.901811e-27, 
    5.391992e-26, -2.695996e-25, -2.205815e-26, -1.347998e-25, 9.803622e-27, 
    2.524433e-25, 9.803622e-27, 9.558531e-26, 7.352717e-27, -2.426396e-25, 
    -1.053889e-25, 2.450905e-26, 3.431268e-26, 2.450906e-27, 1.642107e-25, 
    -3.921449e-26, -1.274471e-25, -3.431268e-26, -1.960724e-26, 
    -4.166539e-26, 5.391992e-26, 6.862535e-26, -2.695996e-26, 4.41163e-26, 
    -7.597807e-26, -1.29898e-25, -1.960724e-26, -9.803622e-27, -7.597807e-26, 
    1.470543e-26, 1.323489e-25, -2.548942e-25, 1.789161e-25, 1.985233e-25, 
    4.41163e-26, 1.053889e-25, -2.941087e-25, -5.882173e-26, 4.41163e-26, 
    -2.205815e-26, 1.54407e-25, -2.377378e-25, -8.82326e-26, 1.176435e-25, 
    1.225453e-26, -1.323489e-25, -7.352717e-26, -1.323489e-25, -1.176435e-25, 
    -1.691125e-25, 3.063632e-25, -2.695996e-26, 1.789161e-25, -4.191048e-25, 
    -1.053889e-25, 5.391992e-26, -1.176435e-25, 1.960724e-25, 2.941087e-26, 
    8.578169e-26, 4.901811e-26, -4.901811e-27, -1.102908e-25, 3.676358e-26, 
    -3.921449e-26, 4.901811e-26, 1.249962e-25, -3.676358e-26, 2.205815e-26, 
    -4.41163e-26, -7.597807e-26, -1.715634e-25, 1.200944e-25, -7.352717e-26, 
    -3.333231e-25, 1.911706e-25, -1.225453e-25, -2.867559e-25, -7.352717e-27, 
    9.803622e-26, -5.146902e-26, 1.200944e-25, 4.901811e-27, 2.450906e-27,
  2.781949e-32, 2.781946e-32, 2.781947e-32, 2.781944e-32, 2.781946e-32, 
    2.781944e-32, 2.781948e-32, 2.781946e-32, 2.781948e-32, 2.781949e-32, 
    2.78194e-32, 2.781944e-32, 2.781935e-32, 2.781938e-32, 2.781931e-32, 
    2.781936e-32, 2.78193e-32, 2.781931e-32, 2.781928e-32, 2.781929e-32, 
    2.781924e-32, 2.781927e-32, 2.781922e-32, 2.781925e-32, 2.781925e-32, 
    2.781927e-32, 2.781943e-32, 2.781941e-32, 2.781944e-32, 2.781943e-32, 
    2.781943e-32, 2.781946e-32, 2.781947e-32, 2.781949e-32, 2.781949e-32, 
    2.781947e-32, 2.781943e-32, 2.781944e-32, 2.781941e-32, 2.781941e-32, 
    2.781937e-32, 2.781939e-32, 2.781932e-32, 2.781934e-32, 2.781928e-32, 
    2.78193e-32, 2.781929e-32, 2.781929e-32, 2.781929e-32, 2.781931e-32, 
    2.78193e-32, 2.781932e-32, 2.781938e-32, 2.781936e-32, 2.781943e-32, 
    2.781946e-32, 2.781948e-32, 2.78195e-32, 2.78195e-32, 2.78195e-32, 
    2.781947e-32, 2.781945e-32, 2.781943e-32, 2.781942e-32, 2.781941e-32, 
    2.781938e-32, 2.781936e-32, 2.781932e-32, 2.781933e-32, 2.781931e-32, 
    2.78193e-32, 2.781928e-32, 2.781928e-32, 2.781928e-32, 2.781931e-32, 
    2.781929e-32, 2.781933e-32, 2.781932e-32, 2.781941e-32, 2.781944e-32, 
    2.781946e-32, 2.781947e-32, 2.78195e-32, 2.781948e-32, 2.781948e-32, 
    2.781946e-32, 2.781945e-32, 2.781946e-32, 2.781942e-32, 2.781943e-32, 
    2.781936e-32, 2.781939e-32, 2.78193e-32, 2.781932e-32, 2.78193e-32, 
    2.781931e-32, 2.781929e-32, 2.781931e-32, 2.781927e-32, 2.781926e-32, 
    2.781927e-32, 2.781925e-32, 2.781931e-32, 2.781929e-32, 2.781946e-32, 
    2.781946e-32, 2.781945e-32, 2.781947e-32, 2.781948e-32, 2.781949e-32, 
    2.781948e-32, 2.781947e-32, 2.781945e-32, 2.781944e-32, 2.781943e-32, 
    2.781941e-32, 2.781938e-32, 2.781935e-32, 2.781932e-32, 2.781931e-32, 
    2.781931e-32, 2.781931e-32, 2.781932e-32, 2.781932e-32, 2.781927e-32, 
    2.78193e-32, 2.781925e-32, 2.781926e-32, 2.781928e-32, 2.781926e-32, 
    2.781946e-32, 2.781946e-32, 2.781948e-32, 2.781947e-32, 2.78195e-32, 
    2.781948e-32, 2.781947e-32, 2.781943e-32, 2.781943e-32, 2.781942e-32, 
    2.781941e-32, 2.781939e-32, 2.781936e-32, 2.781933e-32, 2.78193e-32, 
    2.78193e-32, 2.78193e-32, 2.78193e-32, 2.781931e-32, 2.781929e-32, 
    2.781929e-32, 2.78193e-32, 2.781926e-32, 2.781927e-32, 2.781926e-32, 
    2.781926e-32, 2.781946e-32, 2.781945e-32, 2.781946e-32, 2.781945e-32, 
    2.781945e-32, 2.781942e-32, 2.781941e-32, 2.781937e-32, 2.781939e-32, 
    2.781936e-32, 2.781938e-32, 2.781938e-32, 2.781936e-32, 2.781938e-32, 
    2.781933e-32, 2.781936e-32, 2.78193e-32, 2.781933e-32, 2.781929e-32, 
    2.78193e-32, 2.781929e-32, 2.781928e-32, 2.781926e-32, 2.781924e-32, 
    2.781925e-32, 2.781923e-32, 2.781944e-32, 2.781942e-32, 2.781943e-32, 
    2.781941e-32, 2.78194e-32, 2.781938e-32, 2.781935e-32, 2.781936e-32, 
    2.781933e-32, 2.781933e-32, 2.781937e-32, 2.781934e-32, 2.781941e-32, 
    2.781941e-32, 2.781941e-32, 2.781943e-32, 2.781936e-32, 2.78194e-32, 
    2.781932e-32, 2.781934e-32, 2.781928e-32, 2.781931e-32, 2.781925e-32, 
    2.781922e-32, 2.78192e-32, 2.781917e-32, 2.781942e-32, 2.781943e-32, 
    2.781941e-32, 2.781939e-32, 2.781937e-32, 2.781934e-32, 2.781934e-32, 
    2.781933e-32, 2.781932e-32, 2.781931e-32, 2.781933e-32, 2.781931e-32, 
    2.78194e-32, 2.781935e-32, 2.781943e-32, 2.781941e-32, 2.781939e-32, 
    2.78194e-32, 2.781936e-32, 2.781935e-32, 2.781932e-32, 2.781933e-32, 
    2.781923e-32, 2.781928e-32, 2.781915e-32, 2.781918e-32, 2.781943e-32, 
    2.781942e-32, 2.781938e-32, 2.78194e-32, 2.781934e-32, 2.781933e-32, 
    2.781932e-32, 2.78193e-32, 2.78193e-32, 2.781929e-32, 2.781931e-32, 
    2.781929e-32, 2.781934e-32, 2.781932e-32, 2.781938e-32, 2.781937e-32, 
    2.781937e-32, 2.781938e-32, 2.781936e-32, 2.781933e-32, 2.781933e-32, 
    2.781933e-32, 2.78193e-32, 2.781934e-32, 2.781922e-32, 2.78193e-32, 
    2.781941e-32, 2.781938e-32, 2.781938e-32, 2.781939e-32, 2.781933e-32, 
    2.781935e-32, 2.781929e-32, 2.781931e-32, 2.781928e-32, 2.78193e-32, 
    2.78193e-32, 2.781931e-32, 2.781932e-32, 2.781935e-32, 2.781937e-32, 
    2.781938e-32, 2.781938e-32, 2.781936e-32, 2.781933e-32, 2.78193e-32, 
    2.781931e-32, 2.781928e-32, 2.781934e-32, 2.781932e-32, 2.781933e-32, 
    2.78193e-32, 2.781936e-32, 2.781931e-32, 2.781937e-32, 2.781937e-32, 
    2.781935e-32, 2.781932e-32, 2.781931e-32, 2.78193e-32, 2.781931e-32, 
    2.781933e-32, 2.781933e-32, 2.781935e-32, 2.781936e-32, 2.781937e-32, 
    2.781938e-32, 2.781937e-32, 2.781936e-32, 2.781933e-32, 2.781931e-32, 
    2.781928e-32, 2.781927e-32, 2.781924e-32, 2.781926e-32, 2.781922e-32, 
    2.781926e-32, 2.78192e-32, 2.781931e-32, 2.781926e-32, 2.781935e-32, 
    2.781934e-32, 2.781932e-32, 2.781928e-32, 2.781931e-32, 2.781928e-32, 
    2.781933e-32, 2.781936e-32, 2.781937e-32, 2.781938e-32, 2.781937e-32, 
    2.781937e-32, 2.781936e-32, 2.781936e-32, 2.781933e-32, 2.781935e-32, 
    2.78193e-32, 2.781928e-32, 2.781923e-32, 2.78192e-32, 2.781916e-32, 
    2.781915e-32, 2.781914e-32, 2.781914e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N_TO_SOIL1N =
  3.097809e-15, 3.1062e-15, 3.10457e-15, 3.111332e-15, 3.107583e-15, 
    3.112009e-15, 3.099512e-15, 3.106533e-15, 3.102052e-15, 3.098566e-15, 
    3.124436e-15, 3.111634e-15, 3.137723e-15, 3.129573e-15, 3.150032e-15, 
    3.136454e-15, 3.152768e-15, 3.149643e-15, 3.159051e-15, 3.156357e-15, 
    3.168371e-15, 3.160293e-15, 3.174596e-15, 3.166444e-15, 3.167719e-15, 
    3.160026e-15, 3.114215e-15, 3.122842e-15, 3.113703e-15, 3.114934e-15, 
    3.114382e-15, 3.10766e-15, 3.104268e-15, 3.097169e-15, 3.098459e-15, 
    3.103674e-15, 3.115487e-15, 3.111481e-15, 3.12158e-15, 3.121352e-15, 
    3.132578e-15, 3.127519e-15, 3.146364e-15, 3.141014e-15, 3.15647e-15, 
    3.152585e-15, 3.156287e-15, 3.155164e-15, 3.156301e-15, 3.150603e-15, 
    3.153045e-15, 3.14803e-15, 3.128466e-15, 3.13422e-15, 3.117044e-15, 
    3.106694e-15, 3.09982e-15, 3.094936e-15, 3.095626e-15, 3.096942e-15, 
    3.103704e-15, 3.110059e-15, 3.114898e-15, 3.118133e-15, 3.121319e-15, 
    3.130949e-15, 3.136047e-15, 3.147445e-15, 3.145391e-15, 3.148871e-15, 
    3.152198e-15, 3.157777e-15, 3.15686e-15, 3.159316e-15, 3.148781e-15, 
    3.155783e-15, 3.14422e-15, 3.147384e-15, 3.122176e-15, 3.112562e-15, 
    3.108465e-15, 3.104883e-15, 3.096157e-15, 3.102184e-15, 3.099808e-15, 
    3.105461e-15, 3.109049e-15, 3.107275e-15, 3.118221e-15, 3.113967e-15, 
    3.13635e-15, 3.126716e-15, 3.15181e-15, 3.145813e-15, 3.153247e-15, 
    3.149455e-15, 3.155951e-15, 3.150105e-15, 3.160231e-15, 3.162433e-15, 
    3.160928e-15, 3.166711e-15, 3.149781e-15, 3.156286e-15, 3.107225e-15, 
    3.107514e-15, 3.108863e-15, 3.102932e-15, 3.102569e-15, 3.097133e-15, 
    3.101971e-15, 3.10403e-15, 3.109257e-15, 3.112346e-15, 3.115282e-15, 
    3.121733e-15, 3.12893e-15, 3.138986e-15, 3.146202e-15, 3.151036e-15, 
    3.148072e-15, 3.150689e-15, 3.147764e-15, 3.146393e-15, 3.161607e-15, 
    3.153067e-15, 3.165879e-15, 3.165171e-15, 3.159374e-15, 3.165251e-15, 
    3.107717e-15, 3.106052e-15, 3.100264e-15, 3.104794e-15, 3.096541e-15, 
    3.10116e-15, 3.103815e-15, 3.114054e-15, 3.116304e-15, 3.118387e-15, 
    3.122501e-15, 3.127778e-15, 3.137024e-15, 3.14506e-15, 3.152392e-15, 
    3.151855e-15, 3.152044e-15, 3.15368e-15, 3.149626e-15, 3.154346e-15, 
    3.155137e-15, 3.153067e-15, 3.165076e-15, 3.161647e-15, 3.165156e-15, 
    3.162924e-15, 3.106593e-15, 3.109395e-15, 3.107881e-15, 3.110728e-15, 
    3.108722e-15, 3.117636e-15, 3.120306e-15, 3.132793e-15, 3.127673e-15, 
    3.135823e-15, 3.128502e-15, 3.129799e-15, 3.136085e-15, 3.128899e-15, 
    3.144616e-15, 3.13396e-15, 3.153744e-15, 3.143112e-15, 3.15441e-15, 
    3.15236e-15, 3.155754e-15, 3.158791e-15, 3.162611e-15, 3.169653e-15, 
    3.168023e-15, 3.17391e-15, 3.113572e-15, 3.117202e-15, 3.116885e-15, 
    3.120683e-15, 3.123491e-15, 3.129576e-15, 3.139323e-15, 3.13566e-15, 
    3.142386e-15, 3.143733e-15, 3.133517e-15, 3.13979e-15, 3.119632e-15, 
    3.122891e-15, 3.120952e-15, 3.113857e-15, 3.136502e-15, 3.124888e-15, 
    3.14632e-15, 3.140041e-15, 3.158357e-15, 3.149251e-15, 3.167125e-15, 
    3.17475e-15, 3.181926e-15, 3.190294e-15, 3.119185e-15, 3.116719e-15, 
    3.121135e-15, 3.127239e-15, 3.132903e-15, 3.140424e-15, 3.141194e-15, 
    3.142601e-15, 3.146246e-15, 3.14931e-15, 3.143044e-15, 3.150078e-15, 
    3.123643e-15, 3.13751e-15, 3.115784e-15, 3.122331e-15, 3.12688e-15, 
    3.124886e-15, 3.135241e-15, 3.137679e-15, 3.147576e-15, 3.142463e-15, 
    3.172867e-15, 3.159429e-15, 3.196666e-15, 3.186277e-15, 3.115856e-15, 
    3.119177e-15, 3.130721e-15, 3.125231e-15, 3.140926e-15, 3.144783e-15, 
    3.147919e-15, 3.151923e-15, 3.152357e-15, 3.154728e-15, 3.150841e-15, 
    3.154576e-15, 3.14044e-15, 3.146759e-15, 3.129405e-15, 3.133632e-15, 
    3.131688e-15, 3.129554e-15, 3.136138e-15, 3.143143e-15, 3.143295e-15, 
    3.145538e-15, 3.151854e-15, 3.14099e-15, 3.174594e-15, 3.153852e-15, 
    3.122797e-15, 3.129182e-15, 3.130097e-15, 3.127624e-15, 3.144396e-15, 
    3.138324e-15, 3.154671e-15, 3.150256e-15, 3.157489e-15, 3.153896e-15, 
    3.153367e-15, 3.148749e-15, 3.145873e-15, 3.138602e-15, 3.13268e-15, 
    3.127983e-15, 3.129076e-15, 3.134235e-15, 3.143572e-15, 3.152395e-15, 
    3.150462e-15, 3.15694e-15, 3.139789e-15, 3.146983e-15, 3.144202e-15, 
    3.151452e-15, 3.135562e-15, 3.149087e-15, 3.1321e-15, 3.133591e-15, 
    3.138203e-15, 3.147469e-15, 3.149522e-15, 3.151708e-15, 3.15036e-15, 
    3.143807e-15, 3.142736e-15, 3.138092e-15, 3.136807e-15, 3.133267e-15, 
    3.130333e-15, 3.133013e-15, 3.135825e-15, 3.143811e-15, 3.151001e-15, 
    3.158833e-15, 3.16075e-15, 3.169882e-15, 3.162445e-15, 3.174709e-15, 
    3.164278e-15, 3.182329e-15, 3.149874e-15, 3.163977e-15, 3.138414e-15, 
    3.141173e-15, 3.146155e-15, 3.157582e-15, 3.151418e-15, 3.158627e-15, 
    3.142695e-15, 3.134411e-15, 3.13227e-15, 3.128268e-15, 3.132362e-15, 
    3.132029e-15, 3.135944e-15, 3.134686e-15, 3.144077e-15, 3.139035e-15, 
    3.153353e-15, 3.158571e-15, 3.173292e-15, 3.182301e-15, 3.191464e-15, 
    3.195505e-15, 3.196734e-15, 3.197248e-15 ;

 LITR2N_vr =
  1.592819e-05, 1.592817e-05, 1.592817e-05, 1.592816e-05, 1.592817e-05, 
    1.592816e-05, 1.592818e-05, 1.592817e-05, 1.592818e-05, 1.592818e-05, 
    1.592813e-05, 1.592816e-05, 1.592811e-05, 1.592812e-05, 1.592808e-05, 
    1.592811e-05, 1.592808e-05, 1.592808e-05, 1.592806e-05, 1.592807e-05, 
    1.592805e-05, 1.592806e-05, 1.592803e-05, 1.592805e-05, 1.592805e-05, 
    1.592806e-05, 1.592815e-05, 1.592814e-05, 1.592816e-05, 1.592815e-05, 
    1.592815e-05, 1.592817e-05, 1.592817e-05, 1.592819e-05, 1.592819e-05, 
    1.592818e-05, 1.592815e-05, 1.592816e-05, 1.592814e-05, 1.592814e-05, 
    1.592812e-05, 1.592813e-05, 1.592809e-05, 1.59281e-05, 1.592807e-05, 
    1.592808e-05, 1.592807e-05, 1.592807e-05, 1.592807e-05, 1.592808e-05, 
    1.592808e-05, 1.592809e-05, 1.592813e-05, 1.592811e-05, 1.592815e-05, 
    1.592817e-05, 1.592818e-05, 1.592819e-05, 1.592819e-05, 1.592819e-05, 
    1.592818e-05, 1.592816e-05, 1.592815e-05, 1.592815e-05, 1.592814e-05, 
    1.592812e-05, 1.592811e-05, 1.592809e-05, 1.592809e-05, 1.592808e-05, 
    1.592808e-05, 1.592807e-05, 1.592807e-05, 1.592806e-05, 1.592808e-05, 
    1.592807e-05, 1.592809e-05, 1.592809e-05, 1.592814e-05, 1.592816e-05, 
    1.592817e-05, 1.592817e-05, 1.592819e-05, 1.592818e-05, 1.592818e-05, 
    1.592817e-05, 1.592816e-05, 1.592817e-05, 1.592815e-05, 1.592816e-05, 
    1.592811e-05, 1.592813e-05, 1.592808e-05, 1.592809e-05, 1.592808e-05, 
    1.592808e-05, 1.592807e-05, 1.592808e-05, 1.592806e-05, 1.592806e-05, 
    1.592806e-05, 1.592805e-05, 1.592808e-05, 1.592807e-05, 1.592817e-05, 
    1.592817e-05, 1.592816e-05, 1.592818e-05, 1.592818e-05, 1.592819e-05, 
    1.592818e-05, 1.592817e-05, 1.592816e-05, 1.592816e-05, 1.592815e-05, 
    1.592814e-05, 1.592812e-05, 1.59281e-05, 1.592809e-05, 1.592808e-05, 
    1.592809e-05, 1.592808e-05, 1.592809e-05, 1.592809e-05, 1.592806e-05, 
    1.592808e-05, 1.592805e-05, 1.592805e-05, 1.592806e-05, 1.592805e-05, 
    1.592817e-05, 1.592817e-05, 1.592818e-05, 1.592817e-05, 1.592819e-05, 
    1.592818e-05, 1.592818e-05, 1.592815e-05, 1.592815e-05, 1.592815e-05, 
    1.592814e-05, 1.592813e-05, 1.592811e-05, 1.592809e-05, 1.592808e-05, 
    1.592808e-05, 1.592808e-05, 1.592808e-05, 1.592808e-05, 1.592807e-05, 
    1.592807e-05, 1.592808e-05, 1.592805e-05, 1.592806e-05, 1.592805e-05, 
    1.592806e-05, 1.592817e-05, 1.592816e-05, 1.592817e-05, 1.592816e-05, 
    1.592816e-05, 1.592815e-05, 1.592814e-05, 1.592812e-05, 1.592813e-05, 
    1.592811e-05, 1.592813e-05, 1.592812e-05, 1.592811e-05, 1.592812e-05, 
    1.592809e-05, 1.592812e-05, 1.592808e-05, 1.59281e-05, 1.592807e-05, 
    1.592808e-05, 1.592807e-05, 1.592806e-05, 1.592806e-05, 1.592804e-05, 
    1.592805e-05, 1.592804e-05, 1.592816e-05, 1.592815e-05, 1.592815e-05, 
    1.592814e-05, 1.592814e-05, 1.592812e-05, 1.59281e-05, 1.592811e-05, 
    1.59281e-05, 1.59281e-05, 1.592812e-05, 1.59281e-05, 1.592814e-05, 
    1.592814e-05, 1.592814e-05, 1.592816e-05, 1.592811e-05, 1.592813e-05, 
    1.592809e-05, 1.59281e-05, 1.592807e-05, 1.592808e-05, 1.592805e-05, 
    1.592803e-05, 1.592802e-05, 1.5928e-05, 1.592814e-05, 1.592815e-05, 
    1.592814e-05, 1.592813e-05, 1.592812e-05, 1.59281e-05, 1.59281e-05, 
    1.59281e-05, 1.592809e-05, 1.592808e-05, 1.59281e-05, 1.592808e-05, 
    1.592814e-05, 1.592811e-05, 1.592815e-05, 1.592814e-05, 1.592813e-05, 
    1.592813e-05, 1.592811e-05, 1.592811e-05, 1.592809e-05, 1.59281e-05, 
    1.592804e-05, 1.592806e-05, 1.592799e-05, 1.592801e-05, 1.592815e-05, 
    1.592814e-05, 1.592812e-05, 1.592813e-05, 1.59281e-05, 1.592809e-05, 
    1.592809e-05, 1.592808e-05, 1.592808e-05, 1.592807e-05, 1.592808e-05, 
    1.592807e-05, 1.59281e-05, 1.592809e-05, 1.592812e-05, 1.592812e-05, 
    1.592812e-05, 1.592812e-05, 1.592811e-05, 1.59281e-05, 1.59281e-05, 
    1.592809e-05, 1.592808e-05, 1.59281e-05, 1.592803e-05, 1.592808e-05, 
    1.592814e-05, 1.592812e-05, 1.592812e-05, 1.592813e-05, 1.592809e-05, 
    1.592811e-05, 1.592807e-05, 1.592808e-05, 1.592807e-05, 1.592808e-05, 
    1.592808e-05, 1.592808e-05, 1.592809e-05, 1.592811e-05, 1.592812e-05, 
    1.592813e-05, 1.592812e-05, 1.592811e-05, 1.59281e-05, 1.592808e-05, 
    1.592808e-05, 1.592807e-05, 1.59281e-05, 1.592809e-05, 1.592809e-05, 
    1.592808e-05, 1.592811e-05, 1.592808e-05, 1.592812e-05, 1.592812e-05, 
    1.592811e-05, 1.592809e-05, 1.592808e-05, 1.592808e-05, 1.592808e-05, 
    1.59281e-05, 1.59281e-05, 1.592811e-05, 1.592811e-05, 1.592812e-05, 
    1.592812e-05, 1.592812e-05, 1.592811e-05, 1.59281e-05, 1.592808e-05, 
    1.592806e-05, 1.592806e-05, 1.592804e-05, 1.592806e-05, 1.592803e-05, 
    1.592805e-05, 1.592802e-05, 1.592808e-05, 1.592806e-05, 1.592811e-05, 
    1.59281e-05, 1.592809e-05, 1.592807e-05, 1.592808e-05, 1.592807e-05, 
    1.59281e-05, 1.592811e-05, 1.592812e-05, 1.592813e-05, 1.592812e-05, 
    1.592812e-05, 1.592811e-05, 1.592811e-05, 1.59281e-05, 1.59281e-05, 
    1.592808e-05, 1.592807e-05, 1.592804e-05, 1.592802e-05, 1.5928e-05, 
    1.592799e-05, 1.592799e-05, 1.592799e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2_HR =
  1.11921e-13, 1.122242e-13, 1.121653e-13, 1.124096e-13, 1.122741e-13, 
    1.12434e-13, 1.119825e-13, 1.122362e-13, 1.120743e-13, 1.119484e-13, 
    1.12883e-13, 1.124205e-13, 1.133631e-13, 1.130686e-13, 1.138078e-13, 
    1.133172e-13, 1.139066e-13, 1.137937e-13, 1.141336e-13, 1.140363e-13, 
    1.144703e-13, 1.141785e-13, 1.146953e-13, 1.144007e-13, 1.144468e-13, 
    1.141689e-13, 1.125137e-13, 1.128254e-13, 1.124952e-13, 1.125397e-13, 
    1.125198e-13, 1.122769e-13, 1.121544e-13, 1.118979e-13, 1.119445e-13, 
    1.121329e-13, 1.125597e-13, 1.12415e-13, 1.127798e-13, 1.127716e-13, 
    1.131772e-13, 1.129944e-13, 1.136753e-13, 1.13482e-13, 1.140404e-13, 
    1.139e-13, 1.140338e-13, 1.139932e-13, 1.140343e-13, 1.138284e-13, 
    1.139166e-13, 1.137354e-13, 1.130286e-13, 1.132365e-13, 1.12616e-13, 
    1.12242e-13, 1.119936e-13, 1.118172e-13, 1.118421e-13, 1.118897e-13, 
    1.12134e-13, 1.123636e-13, 1.125384e-13, 1.126553e-13, 1.127704e-13, 
    1.131183e-13, 1.133025e-13, 1.137143e-13, 1.136401e-13, 1.137658e-13, 
    1.13886e-13, 1.140876e-13, 1.140545e-13, 1.141432e-13, 1.137626e-13, 
    1.140156e-13, 1.135978e-13, 1.137121e-13, 1.128014e-13, 1.12454e-13, 
    1.12306e-13, 1.121766e-13, 1.118613e-13, 1.120791e-13, 1.119932e-13, 
    1.121974e-13, 1.123271e-13, 1.12263e-13, 1.126585e-13, 1.125048e-13, 
    1.133134e-13, 1.129654e-13, 1.13872e-13, 1.136553e-13, 1.13924e-13, 
    1.137869e-13, 1.140216e-13, 1.138104e-13, 1.141763e-13, 1.142558e-13, 
    1.142014e-13, 1.144104e-13, 1.137987e-13, 1.140337e-13, 1.122612e-13, 
    1.122716e-13, 1.123204e-13, 1.121061e-13, 1.12093e-13, 1.118966e-13, 
    1.120714e-13, 1.121458e-13, 1.123346e-13, 1.124462e-13, 1.125523e-13, 
    1.127854e-13, 1.130454e-13, 1.134087e-13, 1.136694e-13, 1.13844e-13, 
    1.13737e-13, 1.138315e-13, 1.137258e-13, 1.136763e-13, 1.14226e-13, 
    1.139174e-13, 1.143803e-13, 1.143547e-13, 1.141453e-13, 1.143576e-13, 
    1.12279e-13, 1.122188e-13, 1.120097e-13, 1.121734e-13, 1.118752e-13, 
    1.120421e-13, 1.12138e-13, 1.125079e-13, 1.125892e-13, 1.126645e-13, 
    1.128131e-13, 1.130037e-13, 1.133378e-13, 1.136282e-13, 1.138931e-13, 
    1.138737e-13, 1.138805e-13, 1.139396e-13, 1.137931e-13, 1.139636e-13, 
    1.139922e-13, 1.139174e-13, 1.143513e-13, 1.142274e-13, 1.143542e-13, 
    1.142736e-13, 1.122384e-13, 1.123396e-13, 1.122849e-13, 1.123878e-13, 
    1.123153e-13, 1.126373e-13, 1.127338e-13, 1.13185e-13, 1.13e-13, 
    1.132944e-13, 1.130299e-13, 1.130768e-13, 1.133039e-13, 1.130442e-13, 
    1.136121e-13, 1.132271e-13, 1.139419e-13, 1.135578e-13, 1.139659e-13, 
    1.138919e-13, 1.140145e-13, 1.141242e-13, 1.142623e-13, 1.145167e-13, 
    1.144578e-13, 1.146705e-13, 1.124905e-13, 1.126217e-13, 1.126102e-13, 
    1.127474e-13, 1.128489e-13, 1.130687e-13, 1.134209e-13, 1.132885e-13, 
    1.135315e-13, 1.135802e-13, 1.132111e-13, 1.134378e-13, 1.127095e-13, 
    1.128272e-13, 1.127572e-13, 1.125008e-13, 1.133189e-13, 1.128993e-13, 
    1.136737e-13, 1.134468e-13, 1.141086e-13, 1.137796e-13, 1.144254e-13, 
    1.147008e-13, 1.149601e-13, 1.152624e-13, 1.126933e-13, 1.126042e-13, 
    1.127638e-13, 1.129843e-13, 1.131889e-13, 1.134606e-13, 1.134885e-13, 
    1.135393e-13, 1.13671e-13, 1.137817e-13, 1.135553e-13, 1.138095e-13, 
    1.128544e-13, 1.133554e-13, 1.125704e-13, 1.128069e-13, 1.129713e-13, 
    1.128993e-13, 1.132734e-13, 1.133615e-13, 1.137191e-13, 1.135343e-13, 
    1.146328e-13, 1.141473e-13, 1.154926e-13, 1.151173e-13, 1.12573e-13, 
    1.12693e-13, 1.131101e-13, 1.129117e-13, 1.134788e-13, 1.136181e-13, 
    1.137314e-13, 1.138761e-13, 1.138918e-13, 1.139775e-13, 1.13837e-13, 
    1.139719e-13, 1.134612e-13, 1.136895e-13, 1.130625e-13, 1.132152e-13, 
    1.13145e-13, 1.130679e-13, 1.133058e-13, 1.135589e-13, 1.135644e-13, 
    1.136454e-13, 1.138736e-13, 1.134811e-13, 1.146952e-13, 1.139458e-13, 
    1.128238e-13, 1.130545e-13, 1.130876e-13, 1.129982e-13, 1.136041e-13, 
    1.133848e-13, 1.139754e-13, 1.138159e-13, 1.140772e-13, 1.139474e-13, 
    1.139283e-13, 1.137614e-13, 1.136575e-13, 1.133948e-13, 1.131809e-13, 
    1.130112e-13, 1.130506e-13, 1.13237e-13, 1.135744e-13, 1.138931e-13, 
    1.138233e-13, 1.140574e-13, 1.134377e-13, 1.136976e-13, 1.135971e-13, 
    1.138591e-13, 1.13285e-13, 1.137736e-13, 1.131599e-13, 1.132138e-13, 
    1.133804e-13, 1.137152e-13, 1.137893e-13, 1.138683e-13, 1.138196e-13, 
    1.135829e-13, 1.135442e-13, 1.133764e-13, 1.1333e-13, 1.132021e-13, 
    1.130961e-13, 1.131929e-13, 1.132945e-13, 1.13583e-13, 1.138428e-13, 
    1.141258e-13, 1.14195e-13, 1.145249e-13, 1.142562e-13, 1.146993e-13, 
    1.143225e-13, 1.149746e-13, 1.138021e-13, 1.143116e-13, 1.13388e-13, 
    1.134877e-13, 1.136677e-13, 1.140805e-13, 1.138579e-13, 1.141183e-13, 
    1.135427e-13, 1.132434e-13, 1.131661e-13, 1.130215e-13, 1.131694e-13, 
    1.131573e-13, 1.132988e-13, 1.132534e-13, 1.135926e-13, 1.134105e-13, 
    1.139277e-13, 1.141163e-13, 1.146481e-13, 1.149736e-13, 1.153047e-13, 
    1.154507e-13, 1.154951e-13, 1.155137e-13 ;

 LITR3C =
  1.007811e-05, 1.00781e-05, 1.00781e-05, 1.00781e-05, 1.00781e-05, 
    1.00781e-05, 1.007811e-05, 1.00781e-05, 1.007811e-05, 1.007811e-05, 
    1.007808e-05, 1.00781e-05, 1.007806e-05, 1.007807e-05, 1.007805e-05, 
    1.007806e-05, 1.007804e-05, 1.007805e-05, 1.007804e-05, 1.007804e-05, 
    1.007802e-05, 1.007803e-05, 1.007802e-05, 1.007803e-05, 1.007803e-05, 
    1.007804e-05, 1.007809e-05, 1.007808e-05, 1.007809e-05, 1.007809e-05, 
    1.007809e-05, 1.00781e-05, 1.007811e-05, 1.007811e-05, 1.007811e-05, 
    1.007811e-05, 1.007809e-05, 1.00781e-05, 1.007808e-05, 1.007808e-05, 
    1.007807e-05, 1.007808e-05, 1.007805e-05, 1.007806e-05, 1.007804e-05, 
    1.007804e-05, 1.007804e-05, 1.007804e-05, 1.007804e-05, 1.007805e-05, 
    1.007804e-05, 1.007805e-05, 1.007807e-05, 1.007807e-05, 1.007809e-05, 
    1.00781e-05, 1.007811e-05, 1.007812e-05, 1.007812e-05, 1.007811e-05, 
    1.007811e-05, 1.00781e-05, 1.007809e-05, 1.007809e-05, 1.007808e-05, 
    1.007807e-05, 1.007807e-05, 1.007805e-05, 1.007805e-05, 1.007805e-05, 
    1.007804e-05, 1.007804e-05, 1.007804e-05, 1.007804e-05, 1.007805e-05, 
    1.007804e-05, 1.007805e-05, 1.007805e-05, 1.007808e-05, 1.007809e-05, 
    1.00781e-05, 1.00781e-05, 1.007812e-05, 1.007811e-05, 1.007811e-05, 
    1.00781e-05, 1.00781e-05, 1.00781e-05, 1.007809e-05, 1.007809e-05, 
    1.007806e-05, 1.007808e-05, 1.007805e-05, 1.007805e-05, 1.007804e-05, 
    1.007805e-05, 1.007804e-05, 1.007805e-05, 1.007803e-05, 1.007803e-05, 
    1.007803e-05, 1.007803e-05, 1.007805e-05, 1.007804e-05, 1.00781e-05, 
    1.00781e-05, 1.00781e-05, 1.007811e-05, 1.007811e-05, 1.007811e-05, 
    1.007811e-05, 1.007811e-05, 1.00781e-05, 1.00781e-05, 1.007809e-05, 
    1.007808e-05, 1.007807e-05, 1.007806e-05, 1.007805e-05, 1.007805e-05, 
    1.007805e-05, 1.007805e-05, 1.007805e-05, 1.007805e-05, 1.007803e-05, 
    1.007804e-05, 1.007803e-05, 1.007803e-05, 1.007804e-05, 1.007803e-05, 
    1.00781e-05, 1.00781e-05, 1.007811e-05, 1.00781e-05, 1.007812e-05, 
    1.007811e-05, 1.007811e-05, 1.007809e-05, 1.007809e-05, 1.007809e-05, 
    1.007808e-05, 1.007808e-05, 1.007806e-05, 1.007805e-05, 1.007804e-05, 
    1.007805e-05, 1.007805e-05, 1.007804e-05, 1.007805e-05, 1.007804e-05, 
    1.007804e-05, 1.007804e-05, 1.007803e-05, 1.007803e-05, 1.007803e-05, 
    1.007803e-05, 1.00781e-05, 1.00781e-05, 1.00781e-05, 1.00781e-05, 
    1.00781e-05, 1.007809e-05, 1.007809e-05, 1.007807e-05, 1.007808e-05, 
    1.007807e-05, 1.007807e-05, 1.007807e-05, 1.007807e-05, 1.007807e-05, 
    1.007805e-05, 1.007807e-05, 1.007804e-05, 1.007806e-05, 1.007804e-05, 
    1.007804e-05, 1.007804e-05, 1.007804e-05, 1.007803e-05, 1.007802e-05, 
    1.007803e-05, 1.007802e-05, 1.007809e-05, 1.007809e-05, 1.007809e-05, 
    1.007808e-05, 1.007808e-05, 1.007807e-05, 1.007806e-05, 1.007807e-05, 
    1.007806e-05, 1.007806e-05, 1.007807e-05, 1.007806e-05, 1.007809e-05, 
    1.007808e-05, 1.007808e-05, 1.007809e-05, 1.007806e-05, 1.007808e-05, 
    1.007805e-05, 1.007806e-05, 1.007804e-05, 1.007805e-05, 1.007803e-05, 
    1.007802e-05, 1.007801e-05, 1.0078e-05, 1.007809e-05, 1.007809e-05, 
    1.007808e-05, 1.007808e-05, 1.007807e-05, 1.007806e-05, 1.007806e-05, 
    1.007806e-05, 1.007805e-05, 1.007805e-05, 1.007806e-05, 1.007805e-05, 
    1.007808e-05, 1.007806e-05, 1.007809e-05, 1.007808e-05, 1.007808e-05, 
    1.007808e-05, 1.007807e-05, 1.007806e-05, 1.007805e-05, 1.007806e-05, 
    1.007802e-05, 1.007804e-05, 1.007799e-05, 1.0078e-05, 1.007809e-05, 
    1.007809e-05, 1.007807e-05, 1.007808e-05, 1.007806e-05, 1.007805e-05, 
    1.007805e-05, 1.007805e-05, 1.007804e-05, 1.007804e-05, 1.007805e-05, 
    1.007804e-05, 1.007806e-05, 1.007805e-05, 1.007807e-05, 1.007807e-05, 
    1.007807e-05, 1.007807e-05, 1.007807e-05, 1.007806e-05, 1.007806e-05, 
    1.007805e-05, 1.007805e-05, 1.007806e-05, 1.007802e-05, 1.007804e-05, 
    1.007808e-05, 1.007807e-05, 1.007807e-05, 1.007808e-05, 1.007805e-05, 
    1.007806e-05, 1.007804e-05, 1.007805e-05, 1.007804e-05, 1.007804e-05, 
    1.007804e-05, 1.007805e-05, 1.007805e-05, 1.007806e-05, 1.007807e-05, 
    1.007808e-05, 1.007807e-05, 1.007807e-05, 1.007806e-05, 1.007804e-05, 
    1.007805e-05, 1.007804e-05, 1.007806e-05, 1.007805e-05, 1.007805e-05, 
    1.007805e-05, 1.007807e-05, 1.007805e-05, 1.007807e-05, 1.007807e-05, 
    1.007806e-05, 1.007805e-05, 1.007805e-05, 1.007805e-05, 1.007805e-05, 
    1.007806e-05, 1.007806e-05, 1.007806e-05, 1.007806e-05, 1.007807e-05, 
    1.007807e-05, 1.007807e-05, 1.007807e-05, 1.007806e-05, 1.007805e-05, 
    1.007804e-05, 1.007803e-05, 1.007802e-05, 1.007803e-05, 1.007802e-05, 
    1.007803e-05, 1.007801e-05, 1.007805e-05, 1.007803e-05, 1.007806e-05, 
    1.007806e-05, 1.007805e-05, 1.007804e-05, 1.007805e-05, 1.007804e-05, 
    1.007806e-05, 1.007807e-05, 1.007807e-05, 1.007808e-05, 1.007807e-05, 
    1.007807e-05, 1.007807e-05, 1.007807e-05, 1.007806e-05, 1.007806e-05, 
    1.007804e-05, 1.007804e-05, 1.007802e-05, 1.007801e-05, 1.0078e-05, 
    1.007799e-05, 1.007799e-05, 1.007799e-05 ;

 LITR3C_TO_SOIL2C =
  5.596049e-14, 5.611208e-14, 5.608263e-14, 5.620478e-14, 5.613705e-14, 
    5.621701e-14, 5.599125e-14, 5.611807e-14, 5.603714e-14, 5.597417e-14, 
    5.644149e-14, 5.621023e-14, 5.668151e-14, 5.653429e-14, 5.690388e-14, 
    5.665858e-14, 5.69533e-14, 5.689685e-14, 5.706679e-14, 5.701813e-14, 
    5.723516e-14, 5.708924e-14, 5.734761e-14, 5.720035e-14, 5.722338e-14, 
    5.708442e-14, 5.625685e-14, 5.641271e-14, 5.62476e-14, 5.626984e-14, 
    5.625987e-14, 5.613843e-14, 5.607717e-14, 5.594892e-14, 5.597223e-14, 
    5.606643e-14, 5.627984e-14, 5.620746e-14, 5.63899e-14, 5.638578e-14, 
    5.658858e-14, 5.649718e-14, 5.683761e-14, 5.674098e-14, 5.702016e-14, 
    5.694998e-14, 5.701686e-14, 5.699659e-14, 5.701712e-14, 5.691419e-14, 
    5.69583e-14, 5.68677e-14, 5.651429e-14, 5.661824e-14, 5.630796e-14, 
    5.6121e-14, 5.599681e-14, 5.590858e-14, 5.592106e-14, 5.594483e-14, 
    5.606698e-14, 5.618178e-14, 5.626919e-14, 5.632763e-14, 5.638519e-14, 
    5.655915e-14, 5.665125e-14, 5.685713e-14, 5.682003e-14, 5.68829e-14, 
    5.6943e-14, 5.704379e-14, 5.702721e-14, 5.707159e-14, 5.688128e-14, 
    5.700777e-14, 5.679889e-14, 5.685604e-14, 5.640067e-14, 5.6227e-14, 
    5.615298e-14, 5.608829e-14, 5.593065e-14, 5.603952e-14, 5.599661e-14, 
    5.609871e-14, 5.616353e-14, 5.613148e-14, 5.632922e-14, 5.625237e-14, 
    5.66567e-14, 5.648269e-14, 5.6936e-14, 5.682765e-14, 5.696196e-14, 
    5.689345e-14, 5.70108e-14, 5.690519e-14, 5.708811e-14, 5.712789e-14, 
    5.710071e-14, 5.720517e-14, 5.689933e-14, 5.701684e-14, 5.613057e-14, 
    5.61358e-14, 5.616017e-14, 5.605303e-14, 5.604648e-14, 5.594828e-14, 
    5.603568e-14, 5.607287e-14, 5.61673e-14, 5.62231e-14, 5.627613e-14, 
    5.639267e-14, 5.652267e-14, 5.670432e-14, 5.683468e-14, 5.6922e-14, 
    5.686847e-14, 5.691573e-14, 5.686289e-14, 5.683813e-14, 5.711298e-14, 
    5.69587e-14, 5.719015e-14, 5.717736e-14, 5.707263e-14, 5.71788e-14, 
    5.613947e-14, 5.610939e-14, 5.600485e-14, 5.608667e-14, 5.593758e-14, 
    5.602103e-14, 5.606898e-14, 5.625394e-14, 5.629459e-14, 5.633222e-14, 
    5.640655e-14, 5.650186e-14, 5.666889e-14, 5.681406e-14, 5.694651e-14, 
    5.693681e-14, 5.694022e-14, 5.696978e-14, 5.689653e-14, 5.69818e-14, 
    5.699609e-14, 5.69587e-14, 5.717565e-14, 5.71137e-14, 5.717708e-14, 
    5.713676e-14, 5.611918e-14, 5.616979e-14, 5.614244e-14, 5.619386e-14, 
    5.615762e-14, 5.631865e-14, 5.636689e-14, 5.659246e-14, 5.649997e-14, 
    5.664719e-14, 5.651495e-14, 5.653838e-14, 5.665192e-14, 5.652211e-14, 
    5.680603e-14, 5.661355e-14, 5.697093e-14, 5.677887e-14, 5.698295e-14, 
    5.694594e-14, 5.700724e-14, 5.706209e-14, 5.713111e-14, 5.725832e-14, 
    5.722887e-14, 5.733521e-14, 5.624524e-14, 5.631082e-14, 5.630508e-14, 
    5.63737e-14, 5.642443e-14, 5.653434e-14, 5.671042e-14, 5.664424e-14, 
    5.676575e-14, 5.679009e-14, 5.660553e-14, 5.671886e-14, 5.635472e-14, 
    5.641358e-14, 5.637856e-14, 5.625039e-14, 5.665945e-14, 5.644965e-14, 
    5.683683e-14, 5.672338e-14, 5.705427e-14, 5.688976e-14, 5.721266e-14, 
    5.735039e-14, 5.748002e-14, 5.763119e-14, 5.634663e-14, 5.630208e-14, 
    5.638187e-14, 5.649213e-14, 5.659444e-14, 5.67303e-14, 5.674421e-14, 
    5.676964e-14, 5.683549e-14, 5.689084e-14, 5.677765e-14, 5.690471e-14, 
    5.642717e-14, 5.667766e-14, 5.628521e-14, 5.640346e-14, 5.648565e-14, 
    5.644963e-14, 5.663669e-14, 5.668073e-14, 5.685951e-14, 5.676715e-14, 
    5.731637e-14, 5.707363e-14, 5.774629e-14, 5.755863e-14, 5.62865e-14, 
    5.63465e-14, 5.655503e-14, 5.645585e-14, 5.673939e-14, 5.680905e-14, 
    5.68657e-14, 5.693804e-14, 5.694587e-14, 5.698872e-14, 5.691849e-14, 
    5.698595e-14, 5.673059e-14, 5.684475e-14, 5.653125e-14, 5.66076e-14, 
    5.65725e-14, 5.653395e-14, 5.665288e-14, 5.677942e-14, 5.678217e-14, 
    5.682269e-14, 5.693678e-14, 5.674053e-14, 5.734758e-14, 5.697289e-14, 
    5.641188e-14, 5.652723e-14, 5.654376e-14, 5.649908e-14, 5.680206e-14, 
    5.669237e-14, 5.698768e-14, 5.690793e-14, 5.703858e-14, 5.697367e-14, 
    5.696411e-14, 5.68807e-14, 5.682873e-14, 5.669739e-14, 5.659042e-14, 
    5.650557e-14, 5.652531e-14, 5.66185e-14, 5.678717e-14, 5.694655e-14, 
    5.691164e-14, 5.702866e-14, 5.671884e-14, 5.684879e-14, 5.679855e-14, 
    5.692952e-14, 5.664248e-14, 5.688679e-14, 5.657993e-14, 5.660688e-14, 
    5.669019e-14, 5.685757e-14, 5.689466e-14, 5.693416e-14, 5.69098e-14, 
    5.679143e-14, 5.677208e-14, 5.668817e-14, 5.666498e-14, 5.660101e-14, 
    5.654801e-14, 5.659643e-14, 5.664724e-14, 5.67915e-14, 5.692138e-14, 
    5.706287e-14, 5.709749e-14, 5.726245e-14, 5.712811e-14, 5.734965e-14, 
    5.716121e-14, 5.748731e-14, 5.690101e-14, 5.715577e-14, 5.6694e-14, 
    5.674383e-14, 5.683384e-14, 5.704026e-14, 5.692891e-14, 5.705914e-14, 
    5.677133e-14, 5.662169e-14, 5.658301e-14, 5.651072e-14, 5.658467e-14, 
    5.657866e-14, 5.664938e-14, 5.662666e-14, 5.679629e-14, 5.670521e-14, 
    5.696386e-14, 5.705812e-14, 5.732406e-14, 5.748679e-14, 5.765233e-14, 
    5.772532e-14, 5.774753e-14, 5.775681e-14 ;

 LITR3C_vr =
  0.0005754707, 0.0005754701, 0.0005754702, 0.0005754697, 0.00057547, 
    0.0005754697, 0.0005754706, 0.00057547, 0.0005754704, 0.0005754706, 
    0.0005754688, 0.0005754697, 0.0005754678, 0.0005754684, 0.000575467, 
    0.0005754679, 0.0005754667, 0.000575467, 0.0005754663, 0.0005754665, 
    0.0005754656, 0.0005754662, 0.0005754652, 0.0005754657, 0.0005754657, 
    0.0005754662, 0.0005754695, 0.0005754689, 0.0005754695, 0.0005754695, 
    0.0005754695, 0.00057547, 0.0005754702, 0.0005754707, 0.0005754706, 
    0.0005754703, 0.0005754694, 0.0005754697, 0.000575469, 0.000575469, 
    0.0005754682, 0.0005754685, 0.0005754672, 0.0005754676, 0.0005754665, 
    0.0005754667, 0.0005754665, 0.0005754665, 0.0005754665, 0.0005754669, 
    0.0005754667, 0.0005754671, 0.0005754685, 0.0005754681, 0.0005754693, 
    0.00057547, 0.0005754706, 0.0005754709, 0.0005754709, 0.0005754707, 
    0.0005754703, 0.0005754698, 0.0005754695, 0.0005754692, 0.000575469, 
    0.0005754683, 0.0005754679, 0.0005754671, 0.0005754672, 0.000575467, 
    0.0005754668, 0.0005754664, 0.0005754664, 0.0005754663, 0.000575467, 
    0.0005754665, 0.0005754674, 0.0005754671, 0.0005754689, 0.0005754696, 
    0.0005754699, 0.0005754702, 0.0005754708, 0.0005754704, 0.0005754706, 
    0.0005754702, 0.0005754699, 0.00057547, 0.0005754692, 0.0005754695, 
    0.0005754679, 0.0005754686, 0.0005754668, 0.0005754672, 0.0005754667, 
    0.000575467, 0.0005754665, 0.0005754669, 0.0005754662, 0.000575466, 
    0.0005754661, 0.0005754657, 0.000575467, 0.0005754665, 0.00057547, 
    0.00057547, 0.0005754699, 0.0005754703, 0.0005754703, 0.0005754707, 
    0.0005754704, 0.0005754702, 0.0005754699, 0.0005754696, 0.0005754694, 
    0.0005754689, 0.0005754685, 0.0005754677, 0.0005754672, 0.0005754668, 
    0.0005754671, 0.0005754669, 0.0005754671, 0.0005754672, 0.0005754661, 
    0.0005754667, 0.0005754658, 0.0005754658, 0.0005754663, 0.0005754658, 
    0.00057547, 0.0005754701, 0.0005754705, 0.0005754702, 0.0005754708, 
    0.0005754704, 0.0005754703, 0.0005754695, 0.0005754693, 0.0005754692, 
    0.0005754689, 0.0005754685, 0.0005754679, 0.0005754673, 0.0005754668, 
    0.0005754668, 0.0005754668, 0.0005754667, 0.000575467, 0.0005754666, 
    0.0005754665, 0.0005754667, 0.0005754658, 0.0005754661, 0.0005754658, 
    0.000575466, 0.00057547, 0.0005754699, 0.00057547, 0.0005754697, 
    0.0005754699, 0.0005754693, 0.0005754691, 0.0005754682, 0.0005754685, 
    0.0005754679, 0.0005754685, 0.0005754684, 0.0005754679, 0.0005754685, 
    0.0005754673, 0.0005754681, 0.0005754667, 0.0005754674, 0.0005754666, 
    0.0005754668, 0.0005754665, 0.0005754663, 0.000575466, 0.0005754655, 
    0.0005754656, 0.0005754652, 0.0005754696, 0.0005754693, 0.0005754693, 
    0.0005754691, 0.0005754688, 0.0005754684, 0.0005754677, 0.0005754679, 
    0.0005754675, 0.0005754674, 0.0005754681, 0.0005754677, 0.0005754691, 
    0.0005754689, 0.000575469, 0.0005754695, 0.0005754679, 0.0005754688, 
    0.0005754672, 0.0005754677, 0.0005754663, 0.000575467, 0.0005754657, 
    0.0005754652, 0.0005754646, 0.000575464, 0.0005754692, 0.0005754693, 
    0.000575469, 0.0005754686, 0.0005754682, 0.0005754676, 0.0005754675, 
    0.0005754675, 0.0005754672, 0.000575467, 0.0005754674, 0.0005754669, 
    0.0005754688, 0.0005754678, 0.0005754694, 0.0005754689, 0.0005754686, 
    0.0005754688, 0.000575468, 0.0005754678, 0.0005754671, 0.0005754675, 
    0.0005754653, 0.0005754663, 0.0005754636, 0.0005754643, 0.0005754694, 
    0.0005754692, 0.0005754683, 0.0005754687, 0.0005754676, 0.0005754673, 
    0.0005754671, 0.0005754668, 0.0005754668, 0.0005754666, 0.0005754669, 
    0.0005754666, 0.0005754676, 0.0005754672, 0.0005754684, 0.0005754681, 
    0.0005754682, 0.0005754684, 0.0005754679, 0.0005754674, 0.0005754674, 
    0.0005754672, 0.0005754668, 0.0005754676, 0.0005754652, 0.0005754667, 
    0.0005754689, 0.0005754684, 0.0005754684, 0.0005754685, 0.0005754673, 
    0.0005754678, 0.0005754666, 0.0005754669, 0.0005754664, 0.0005754667, 
    0.0005754667, 0.000575467, 0.0005754672, 0.0005754678, 0.0005754682, 
    0.0005754685, 0.0005754684, 0.0005754681, 0.0005754674, 0.0005754668, 
    0.0005754669, 0.0005754664, 0.0005754677, 0.0005754671, 0.0005754674, 
    0.0005754668, 0.0005754679, 0.000575467, 0.0005754682, 0.0005754681, 
    0.0005754678, 0.0005754671, 0.000575467, 0.0005754668, 0.0005754669, 
    0.0005754674, 0.0005754675, 0.0005754678, 0.0005754679, 0.0005754681, 
    0.0005754684, 0.0005754682, 0.0005754679, 0.0005754674, 0.0005754668, 
    0.0005754663, 0.0005754661, 0.0005754655, 0.000575466, 0.0005754652, 
    0.0005754659, 0.0005754646, 0.000575467, 0.0005754659, 0.0005754678, 
    0.0005754675, 0.0005754672, 0.0005754664, 0.0005754668, 0.0005754663, 
    0.0005754675, 0.0005754681, 0.0005754682, 0.0005754685, 0.0005754682, 
    0.0005754682, 0.0005754679, 0.000575468, 0.0005754674, 0.0005754677, 
    0.0005754667, 0.0005754663, 0.0005754653, 0.0005754646, 0.0005754639, 
    0.0005754636, 0.0005754636, 0.0005754635,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N =
  1.394737e-07, 1.394736e-07, 1.394736e-07, 1.394735e-07, 1.394735e-07, 
    1.394735e-07, 1.394737e-07, 1.394736e-07, 1.394736e-07, 1.394737e-07, 
    1.394732e-07, 1.394735e-07, 1.39473e-07, 1.394732e-07, 1.394728e-07, 
    1.39473e-07, 1.394727e-07, 1.394728e-07, 1.394726e-07, 1.394727e-07, 
    1.394725e-07, 1.394726e-07, 1.394724e-07, 1.394725e-07, 1.394725e-07, 
    1.394726e-07, 1.394734e-07, 1.394733e-07, 1.394734e-07, 1.394734e-07, 
    1.394734e-07, 1.394735e-07, 1.394736e-07, 1.394737e-07, 1.394737e-07, 
    1.394736e-07, 1.394734e-07, 1.394735e-07, 1.394733e-07, 1.394733e-07, 
    1.394731e-07, 1.394732e-07, 1.394729e-07, 1.39473e-07, 1.394727e-07, 
    1.394728e-07, 1.394727e-07, 1.394727e-07, 1.394727e-07, 1.394728e-07, 
    1.394727e-07, 1.394728e-07, 1.394732e-07, 1.394731e-07, 1.394734e-07, 
    1.394736e-07, 1.394737e-07, 1.394738e-07, 1.394738e-07, 1.394737e-07, 
    1.394736e-07, 1.394735e-07, 1.394734e-07, 1.394734e-07, 1.394733e-07, 
    1.394731e-07, 1.39473e-07, 1.394728e-07, 1.394729e-07, 1.394728e-07, 
    1.394728e-07, 1.394727e-07, 1.394727e-07, 1.394726e-07, 1.394728e-07, 
    1.394727e-07, 1.394729e-07, 1.394728e-07, 1.394733e-07, 1.394735e-07, 
    1.394735e-07, 1.394736e-07, 1.394737e-07, 1.394736e-07, 1.394737e-07, 
    1.394736e-07, 1.394735e-07, 1.394735e-07, 1.394734e-07, 1.394734e-07, 
    1.39473e-07, 1.394732e-07, 1.394728e-07, 1.394729e-07, 1.394727e-07, 
    1.394728e-07, 1.394727e-07, 1.394728e-07, 1.394726e-07, 1.394726e-07, 
    1.394726e-07, 1.394725e-07, 1.394728e-07, 1.394727e-07, 1.394735e-07, 
    1.394735e-07, 1.394735e-07, 1.394736e-07, 1.394736e-07, 1.394737e-07, 
    1.394736e-07, 1.394736e-07, 1.394735e-07, 1.394735e-07, 1.394734e-07, 
    1.394733e-07, 1.394732e-07, 1.39473e-07, 1.394729e-07, 1.394728e-07, 
    1.394728e-07, 1.394728e-07, 1.394728e-07, 1.394729e-07, 1.394726e-07, 
    1.394727e-07, 1.394725e-07, 1.394725e-07, 1.394726e-07, 1.394725e-07, 
    1.394735e-07, 1.394736e-07, 1.394737e-07, 1.394736e-07, 1.394737e-07, 
    1.394737e-07, 1.394736e-07, 1.394734e-07, 1.394734e-07, 1.394734e-07, 
    1.394733e-07, 1.394732e-07, 1.39473e-07, 1.394729e-07, 1.394728e-07, 
    1.394728e-07, 1.394728e-07, 1.394727e-07, 1.394728e-07, 1.394727e-07, 
    1.394727e-07, 1.394727e-07, 1.394725e-07, 1.394726e-07, 1.394725e-07, 
    1.394726e-07, 1.394736e-07, 1.394735e-07, 1.394735e-07, 1.394735e-07, 
    1.394735e-07, 1.394734e-07, 1.394733e-07, 1.394731e-07, 1.394732e-07, 
    1.39473e-07, 1.394732e-07, 1.394732e-07, 1.39473e-07, 1.394732e-07, 
    1.394729e-07, 1.394731e-07, 1.394727e-07, 1.394729e-07, 1.394727e-07, 
    1.394728e-07, 1.394727e-07, 1.394726e-07, 1.394726e-07, 1.394725e-07, 
    1.394725e-07, 1.394724e-07, 1.394734e-07, 1.394734e-07, 1.394734e-07, 
    1.394733e-07, 1.394733e-07, 1.394732e-07, 1.39473e-07, 1.39473e-07, 
    1.394729e-07, 1.394729e-07, 1.394731e-07, 1.39473e-07, 1.394733e-07, 
    1.394733e-07, 1.394733e-07, 1.394734e-07, 1.39473e-07, 1.394732e-07, 
    1.394729e-07, 1.39473e-07, 1.394727e-07, 1.394728e-07, 1.394725e-07, 
    1.394724e-07, 1.394722e-07, 1.394721e-07, 1.394733e-07, 1.394734e-07, 
    1.394733e-07, 1.394732e-07, 1.394731e-07, 1.39473e-07, 1.39473e-07, 
    1.394729e-07, 1.394729e-07, 1.394728e-07, 1.394729e-07, 1.394728e-07, 
    1.394733e-07, 1.39473e-07, 1.394734e-07, 1.394733e-07, 1.394732e-07, 
    1.394732e-07, 1.394731e-07, 1.39473e-07, 1.394728e-07, 1.394729e-07, 
    1.394724e-07, 1.394726e-07, 1.39472e-07, 1.394722e-07, 1.394734e-07, 
    1.394733e-07, 1.394731e-07, 1.394732e-07, 1.39473e-07, 1.394729e-07, 
    1.394728e-07, 1.394728e-07, 1.394728e-07, 1.394727e-07, 1.394728e-07, 
    1.394727e-07, 1.39473e-07, 1.394729e-07, 1.394732e-07, 1.394731e-07, 
    1.394731e-07, 1.394732e-07, 1.39473e-07, 1.394729e-07, 1.394729e-07, 
    1.394729e-07, 1.394728e-07, 1.39473e-07, 1.394724e-07, 1.394727e-07, 
    1.394733e-07, 1.394732e-07, 1.394731e-07, 1.394732e-07, 1.394729e-07, 
    1.39473e-07, 1.394727e-07, 1.394728e-07, 1.394727e-07, 1.394727e-07, 
    1.394727e-07, 1.394728e-07, 1.394729e-07, 1.39473e-07, 1.394731e-07, 
    1.394732e-07, 1.394732e-07, 1.394731e-07, 1.394729e-07, 1.394728e-07, 
    1.394728e-07, 1.394727e-07, 1.39473e-07, 1.394728e-07, 1.394729e-07, 
    1.394728e-07, 1.394731e-07, 1.394728e-07, 1.394731e-07, 1.394731e-07, 
    1.39473e-07, 1.394728e-07, 1.394728e-07, 1.394728e-07, 1.394728e-07, 
    1.394729e-07, 1.394729e-07, 1.39473e-07, 1.39473e-07, 1.394731e-07, 
    1.394731e-07, 1.394731e-07, 1.39473e-07, 1.394729e-07, 1.394728e-07, 
    1.394726e-07, 1.394726e-07, 1.394724e-07, 1.394726e-07, 1.394724e-07, 
    1.394725e-07, 1.394722e-07, 1.394728e-07, 1.394726e-07, 1.39473e-07, 
    1.39473e-07, 1.394729e-07, 1.394727e-07, 1.394728e-07, 1.394726e-07, 
    1.394729e-07, 1.394731e-07, 1.394731e-07, 1.394732e-07, 1.394731e-07, 
    1.394731e-07, 1.39473e-07, 1.394731e-07, 1.394729e-07, 1.39473e-07, 
    1.394727e-07, 1.394726e-07, 1.394724e-07, 1.394722e-07, 1.394721e-07, 
    1.39472e-07, 1.39472e-07, 1.39472e-07 ;

 LITR3N_TNDNCY_VERT_TRANS =
  2.941087e-26, -6.372354e-26, 1.654361e-25, 2.695996e-26, 5.269447e-26, 
    3.798904e-26, 1.225453e-26, -3.553813e-26, -5.146902e-26, 1.397016e-25, 
    -8.455624e-26, 9.558531e-26, 7.352717e-27, -4.901811e-26, -1.02938e-25, 
    -9.068351e-26, 4.901811e-26, 3.676358e-26, 5.882173e-26, 1.139671e-25, 
    -3.063632e-26, -8.700715e-26, 5.514538e-26, 1.090653e-25, 1.470543e-25, 
    -4.901811e-26, -4.289085e-26, -5.759628e-26, -3.431268e-26, 1.115162e-25, 
    3.676358e-26, -8.578169e-26, 2.450906e-27, -2.941087e-26, -1.139671e-25, 
    -1.225453e-26, 1.384762e-25, -4.779266e-26, 7.720352e-26, -1.703379e-25, 
    -6.98508e-26, 7.475262e-26, -1.384762e-25, -4.901811e-26, -2.08327e-26, 
    1.127417e-25, -3.676358e-26, 2.941087e-26, 7.107626e-26, 1.421525e-25, 
    -5.269447e-26, -3.676358e-26, -1.911706e-25, -2.08327e-26, 1.188689e-25, 
    8.578169e-27, -5.269447e-26, 4.534175e-26, -1.838179e-26, -7.352717e-27, 
    -3.063632e-26, 3.553813e-26, 1.593089e-26, -1.593089e-26, 1.715634e-26, 
    1.090653e-25, 1.715634e-26, 1.470543e-26, -4.166539e-26, 1.347998e-26, 
    6.73999e-26, -7.107626e-26, -8.087988e-26, 3.431268e-26, -9.068351e-26, 
    2.32836e-26, 6.127264e-26, -2.695996e-26, 1.384762e-25, 8.333079e-26, 
    6.372354e-26, 4.41163e-26, 2.818541e-26, 4.901811e-27, -1.053889e-25, 
    -7.965443e-26, 2.818541e-26, 3.186177e-26, -2.818541e-26, -4.65672e-26, 
    -6.004719e-26, 4.901811e-27, -9.681077e-26, 4.901811e-27, 2.941087e-26, 
    0, 6.98508e-26, -4.534175e-26, 7.965443e-26, 2.450905e-26, 2.08327e-26, 
    2.450906e-27, -4.901811e-27, 1.004871e-25, -4.901811e-26, -9.803622e-26, 
    3.553813e-26, 5.391992e-26, 8.210533e-26, 5.269447e-26, 3.676358e-26, 
    4.043994e-26, -1.262216e-25, 2.573451e-26, -2.695996e-26, -2.941087e-26, 
    4.043994e-26, -1.335744e-25, 2.205815e-26, -2.573451e-26, 3.798904e-26, 
    -7.352717e-26, -3.921449e-26, 1.115162e-25, -4.534175e-26, -5.882173e-26, 
    -7.230172e-26, -8.210533e-26, 1.470543e-26, 0, -9.313441e-26, 
    5.146902e-26, -6.127264e-26, 1.274471e-25, 4.901811e-26, -9.803622e-27, 
    2.450905e-26, -3.921449e-26, -6.862535e-26, -1.262216e-25, -1.311234e-25, 
    7.842898e-26, -7.475262e-26, -3.063632e-26, 5.269447e-26, -9.681077e-26, 
    7.720352e-26, 9.681077e-26, -4.65672e-26, -2.573451e-26, 6.617445e-26, 
    4.166539e-26, 9.926167e-26, -1.225453e-27, 1.200944e-25, 1.225453e-27, 
    9.068351e-26, 3.431268e-26, 2.205815e-26, -8.82326e-26, -1.715634e-26, 
    -7.352717e-27, -2.818541e-26, 3.921449e-26, 1.16418e-25, 7.352717e-27, 
    -2.32836e-26, 6.617445e-26, -1.004871e-25, -4.166539e-26, -3.553813e-26, 
    5.391992e-26, -1.347998e-26, -5.637083e-26, -1.960724e-26, -6.4949e-26, 
    6.127264e-26, -7.597807e-26, 9.558531e-26, 6.372354e-26, 7.720352e-26, 
    9.681077e-26, -1.311234e-25, -4.043994e-26, 1.347998e-25, 1.960724e-26, 
    6.004719e-26, -1.225453e-26, -6.004719e-26, 4.901811e-27, 2.450905e-26, 
    2.205815e-26, -9.190896e-26, -2.450905e-26, 1.347998e-26, 3.308722e-26, 
    1.850434e-25, -5.269447e-26, 2.818541e-26, -2.450905e-26, 2.205815e-26, 
    8.210533e-26, -2.32836e-26, 1.102908e-25, 2.450906e-27, -6.98508e-26, 
    -9.681077e-26, -1.017126e-25, -4.41163e-26, -3.676358e-26, -4.901811e-26, 
    -2.08327e-26, 6.127264e-26, -9.313441e-26, 5.759628e-26, 2.450905e-26, 
    -6.249809e-26, -1.225453e-26, -7.107626e-26, -1.470543e-26, 3.798904e-26, 
    -3.676358e-27, 1.593089e-25, -1.838179e-26, 4.41163e-26, 9.803622e-26, 
    -1.225453e-27, -1.102908e-26, 5.882173e-26, 6.4949e-26, 4.043994e-26, 
    -4.043994e-26, -1.225453e-26, -8.578169e-27, -7.475262e-26, 5.269447e-26, 
    -6.127264e-27, 4.901811e-26, -1.286725e-25, 4.41163e-26, -3.676358e-27, 
    2.818541e-26, 2.450906e-27, 1.764652e-25, 1.715634e-25, 7.842898e-26, 
    2.573451e-26, 1.225453e-25, 1.237707e-25, -4.043994e-26, -3.676358e-26, 
    -3.921449e-26, -2.695996e-26, 5.024356e-26, -2.941087e-26, 1.151926e-25, 
    3.921449e-26, 4.901811e-27, -7.352717e-27, 1.446034e-25, 1.262216e-25, 
    -5.514538e-26, -1.102908e-26, -1.56858e-25, -2.695996e-26, -1.960724e-26, 
    2.695996e-26, 4.289085e-26, 3.308722e-26, 1.347998e-26, 9.803622e-27, 
    -9.926167e-26, 6.127264e-26, -2.450906e-27, 1.838179e-26, -3.431268e-26, 
    -6.127264e-27, 1.29898e-25, -7.352717e-27, -6.617445e-26, -9.681077e-26, 
    6.617445e-26, -3.676358e-27, -7.230172e-26, -7.965443e-26, 1.347998e-26, 
    4.65672e-26, 4.901811e-27, 6.004719e-26, 7.597807e-26, 3.921449e-26, 
    -1.470543e-26, 1.29898e-25, 1.004871e-25, 5.146902e-26, -1.102908e-26, 
    -5.637083e-26, 7.842898e-26, 3.921449e-26, 1.225453e-27, 5.759628e-26, 
    5.759628e-26, -9.681077e-26, 1.347998e-26, -2.205815e-26, -1.090653e-25, 
    6.127264e-26, -1.225453e-27, -5.269447e-26, -3.676358e-27, 5.759628e-26, 
    1.838179e-26, -3.186177e-26, -1.593089e-26, -3.553813e-26, 1.274471e-25, 
    -4.043994e-26, -5.514538e-26, 7.230172e-26, -3.798904e-26, -7.230172e-26, 
    2.941087e-26, -7.720352e-26, 3.798904e-26, -7.475262e-26, 8.087988e-26, 
    3.431268e-26, 1.102908e-26, 7.842898e-26, 6.127264e-27, 6.98508e-26, 
    1.115162e-25, -2.205815e-26, 9.681077e-26, 1.066144e-25, -8.210533e-26, 
    -6.127264e-27, 6.004719e-26,
  1.390975e-32, 1.390973e-32, 1.390973e-32, 1.390972e-32, 1.390973e-32, 
    1.390972e-32, 1.390974e-32, 1.390973e-32, 1.390974e-32, 1.390974e-32, 
    1.39097e-32, 1.390972e-32, 1.390967e-32, 1.390969e-32, 1.390965e-32, 
    1.390968e-32, 1.390965e-32, 1.390965e-32, 1.390964e-32, 1.390964e-32, 
    1.390962e-32, 1.390963e-32, 1.390961e-32, 1.390962e-32, 1.390962e-32, 
    1.390964e-32, 1.390972e-32, 1.39097e-32, 1.390972e-32, 1.390972e-32, 
    1.390972e-32, 1.390973e-32, 1.390973e-32, 1.390975e-32, 1.390974e-32, 
    1.390973e-32, 1.390971e-32, 1.390972e-32, 1.39097e-32, 1.39097e-32, 
    1.390968e-32, 1.390969e-32, 1.390966e-32, 1.390967e-32, 1.390964e-32, 
    1.390965e-32, 1.390964e-32, 1.390965e-32, 1.390964e-32, 1.390965e-32, 
    1.390965e-32, 1.390966e-32, 1.390969e-32, 1.390968e-32, 1.390971e-32, 
    1.390973e-32, 1.390974e-32, 1.390975e-32, 1.390975e-32, 1.390975e-32, 
    1.390973e-32, 1.390972e-32, 1.390972e-32, 1.390971e-32, 1.39097e-32, 
    1.390969e-32, 1.390968e-32, 1.390966e-32, 1.390966e-32, 1.390966e-32, 
    1.390965e-32, 1.390964e-32, 1.390964e-32, 1.390964e-32, 1.390966e-32, 
    1.390964e-32, 1.390966e-32, 1.390966e-32, 1.39097e-32, 1.390972e-32, 
    1.390973e-32, 1.390973e-32, 1.390975e-32, 1.390974e-32, 1.390974e-32, 
    1.390973e-32, 1.390973e-32, 1.390973e-32, 1.390971e-32, 1.390972e-32, 
    1.390968e-32, 1.39097e-32, 1.390965e-32, 1.390966e-32, 1.390965e-32, 
    1.390965e-32, 1.390964e-32, 1.390965e-32, 1.390964e-32, 1.390963e-32, 
    1.390963e-32, 1.390962e-32, 1.390965e-32, 1.390964e-32, 1.390973e-32, 
    1.390973e-32, 1.390973e-32, 1.390974e-32, 1.390974e-32, 1.390975e-32, 
    1.390974e-32, 1.390973e-32, 1.390972e-32, 1.390972e-32, 1.390971e-32, 
    1.39097e-32, 1.390969e-32, 1.390967e-32, 1.390966e-32, 1.390965e-32, 
    1.390966e-32, 1.390965e-32, 1.390966e-32, 1.390966e-32, 1.390963e-32, 
    1.390965e-32, 1.390963e-32, 1.390963e-32, 1.390964e-32, 1.390963e-32, 
    1.390973e-32, 1.390973e-32, 1.390974e-32, 1.390973e-32, 1.390975e-32, 
    1.390974e-32, 1.390973e-32, 1.390972e-32, 1.390971e-32, 1.390971e-32, 
    1.39097e-32, 1.390969e-32, 1.390968e-32, 1.390966e-32, 1.390965e-32, 
    1.390965e-32, 1.390965e-32, 1.390965e-32, 1.390965e-32, 1.390965e-32, 
    1.390965e-32, 1.390965e-32, 1.390963e-32, 1.390963e-32, 1.390963e-32, 
    1.390963e-32, 1.390973e-32, 1.390972e-32, 1.390973e-32, 1.390972e-32, 
    1.390973e-32, 1.390971e-32, 1.390971e-32, 1.390968e-32, 1.390969e-32, 
    1.390968e-32, 1.390969e-32, 1.390969e-32, 1.390968e-32, 1.390969e-32, 
    1.390966e-32, 1.390968e-32, 1.390965e-32, 1.390967e-32, 1.390965e-32, 
    1.390965e-32, 1.390964e-32, 1.390964e-32, 1.390963e-32, 1.390962e-32, 
    1.390962e-32, 1.390961e-32, 1.390972e-32, 1.390971e-32, 1.390971e-32, 
    1.390971e-32, 1.39097e-32, 1.390969e-32, 1.390967e-32, 1.390968e-32, 
    1.390967e-32, 1.390966e-32, 1.390968e-32, 1.390967e-32, 1.390971e-32, 
    1.39097e-32, 1.39097e-32, 1.390972e-32, 1.390968e-32, 1.39097e-32, 
    1.390966e-32, 1.390967e-32, 1.390964e-32, 1.390966e-32, 1.390962e-32, 
    1.390961e-32, 1.39096e-32, 1.390958e-32, 1.390971e-32, 1.390971e-32, 
    1.39097e-32, 1.390969e-32, 1.390968e-32, 1.390967e-32, 1.390967e-32, 
    1.390967e-32, 1.390966e-32, 1.390966e-32, 1.390967e-32, 1.390965e-32, 
    1.39097e-32, 1.390968e-32, 1.390971e-32, 1.39097e-32, 1.390969e-32, 
    1.39097e-32, 1.390968e-32, 1.390967e-32, 1.390966e-32, 1.390967e-32, 
    1.390961e-32, 1.390964e-32, 1.390957e-32, 1.390959e-32, 1.390971e-32, 
    1.390971e-32, 1.390969e-32, 1.39097e-32, 1.390967e-32, 1.390966e-32, 
    1.390966e-32, 1.390965e-32, 1.390965e-32, 1.390965e-32, 1.390965e-32, 
    1.390965e-32, 1.390967e-32, 1.390966e-32, 1.390969e-32, 1.390968e-32, 
    1.390969e-32, 1.390969e-32, 1.390968e-32, 1.390967e-32, 1.390967e-32, 
    1.390966e-32, 1.390965e-32, 1.390967e-32, 1.390961e-32, 1.390965e-32, 
    1.39097e-32, 1.390969e-32, 1.390969e-32, 1.390969e-32, 1.390966e-32, 
    1.390967e-32, 1.390965e-32, 1.390965e-32, 1.390964e-32, 1.390965e-32, 
    1.390965e-32, 1.390966e-32, 1.390966e-32, 1.390967e-32, 1.390968e-32, 
    1.390969e-32, 1.390969e-32, 1.390968e-32, 1.390966e-32, 1.390965e-32, 
    1.390965e-32, 1.390964e-32, 1.390967e-32, 1.390966e-32, 1.390966e-32, 
    1.390965e-32, 1.390968e-32, 1.390966e-32, 1.390968e-32, 1.390968e-32, 
    1.390967e-32, 1.390966e-32, 1.390965e-32, 1.390965e-32, 1.390965e-32, 
    1.390966e-32, 1.390967e-32, 1.390967e-32, 1.390968e-32, 1.390968e-32, 
    1.390969e-32, 1.390968e-32, 1.390968e-32, 1.390966e-32, 1.390965e-32, 
    1.390964e-32, 1.390963e-32, 1.390962e-32, 1.390963e-32, 1.390961e-32, 
    1.390963e-32, 1.39096e-32, 1.390965e-32, 1.390963e-32, 1.390967e-32, 
    1.390967e-32, 1.390966e-32, 1.390964e-32, 1.390965e-32, 1.390964e-32, 
    1.390967e-32, 1.390968e-32, 1.390968e-32, 1.390969e-32, 1.390968e-32, 
    1.390968e-32, 1.390968e-32, 1.390968e-32, 1.390966e-32, 1.390967e-32, 
    1.390965e-32, 1.390964e-32, 1.390961e-32, 1.39096e-32, 1.390958e-32, 
    1.390957e-32, 1.390957e-32, 1.390957e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N_TO_SOIL2N =
  1.548904e-15, 1.5531e-15, 1.552285e-15, 1.555666e-15, 1.553791e-15, 
    1.556005e-15, 1.549756e-15, 1.553266e-15, 1.551026e-15, 1.549283e-15, 
    1.562218e-15, 1.555817e-15, 1.568861e-15, 1.564786e-15, 1.575016e-15, 
    1.568227e-15, 1.576384e-15, 1.574822e-15, 1.579525e-15, 1.578178e-15, 
    1.584185e-15, 1.580147e-15, 1.587298e-15, 1.583222e-15, 1.583859e-15, 
    1.580013e-15, 1.557107e-15, 1.561421e-15, 1.556851e-15, 1.557467e-15, 
    1.557191e-15, 1.55383e-15, 1.552134e-15, 1.548584e-15, 1.549229e-15, 
    1.551837e-15, 1.557744e-15, 1.55574e-15, 1.56079e-15, 1.560676e-15, 
    1.566289e-15, 1.563759e-15, 1.573182e-15, 1.570507e-15, 1.578235e-15, 
    1.576292e-15, 1.578143e-15, 1.577582e-15, 1.57815e-15, 1.575301e-15, 
    1.576522e-15, 1.574015e-15, 1.564233e-15, 1.56711e-15, 1.558522e-15, 
    1.553347e-15, 1.54991e-15, 1.547468e-15, 1.547813e-15, 1.548471e-15, 
    1.551852e-15, 1.555029e-15, 1.557449e-15, 1.559066e-15, 1.560659e-15, 
    1.565475e-15, 1.568024e-15, 1.573722e-15, 1.572695e-15, 1.574436e-15, 
    1.576099e-15, 1.578889e-15, 1.57843e-15, 1.579658e-15, 1.574391e-15, 
    1.577892e-15, 1.57211e-15, 1.573692e-15, 1.561088e-15, 1.556281e-15, 
    1.554232e-15, 1.552442e-15, 1.548078e-15, 1.551092e-15, 1.549904e-15, 
    1.55273e-15, 1.554524e-15, 1.553637e-15, 1.55911e-15, 1.556983e-15, 
    1.568175e-15, 1.563358e-15, 1.575905e-15, 1.572906e-15, 1.576624e-15, 
    1.574727e-15, 1.577976e-15, 1.575052e-15, 1.580115e-15, 1.581216e-15, 
    1.580464e-15, 1.583355e-15, 1.57489e-15, 1.578143e-15, 1.553612e-15, 
    1.553757e-15, 1.554431e-15, 1.551466e-15, 1.551285e-15, 1.548566e-15, 
    1.550986e-15, 1.552015e-15, 1.554629e-15, 1.556173e-15, 1.557641e-15, 
    1.560866e-15, 1.564465e-15, 1.569493e-15, 1.573101e-15, 1.575518e-15, 
    1.574036e-15, 1.575344e-15, 1.573882e-15, 1.573196e-15, 1.580804e-15, 
    1.576533e-15, 1.58294e-15, 1.582586e-15, 1.579687e-15, 1.582625e-15, 
    1.553858e-15, 1.553026e-15, 1.550132e-15, 1.552397e-15, 1.54827e-15, 
    1.55058e-15, 1.551907e-15, 1.557027e-15, 1.558152e-15, 1.559193e-15, 
    1.561251e-15, 1.563889e-15, 1.568512e-15, 1.57253e-15, 1.576196e-15, 
    1.575928e-15, 1.576022e-15, 1.57684e-15, 1.574813e-15, 1.577173e-15, 
    1.577568e-15, 1.576534e-15, 1.582538e-15, 1.580824e-15, 1.582578e-15, 
    1.581462e-15, 1.553297e-15, 1.554698e-15, 1.553941e-15, 1.555364e-15, 
    1.554361e-15, 1.558818e-15, 1.560153e-15, 1.566397e-15, 1.563837e-15, 
    1.567911e-15, 1.564251e-15, 1.5649e-15, 1.568042e-15, 1.564449e-15, 
    1.572308e-15, 1.56698e-15, 1.576872e-15, 1.571556e-15, 1.577205e-15, 
    1.57618e-15, 1.577877e-15, 1.579395e-15, 1.581305e-15, 1.584826e-15, 
    1.584012e-15, 1.586955e-15, 1.556786e-15, 1.558601e-15, 1.558442e-15, 
    1.560342e-15, 1.561746e-15, 1.564788e-15, 1.569662e-15, 1.56783e-15, 
    1.571193e-15, 1.571866e-15, 1.566758e-15, 1.569895e-15, 1.559816e-15, 
    1.561445e-15, 1.560476e-15, 1.556929e-15, 1.568251e-15, 1.562444e-15, 
    1.57316e-15, 1.57002e-15, 1.579179e-15, 1.574625e-15, 1.583563e-15, 
    1.587375e-15, 1.590963e-15, 1.595147e-15, 1.559592e-15, 1.558359e-15, 
    1.560568e-15, 1.56362e-15, 1.566451e-15, 1.570212e-15, 1.570597e-15, 
    1.571301e-15, 1.573123e-15, 1.574655e-15, 1.571522e-15, 1.575039e-15, 
    1.561821e-15, 1.568755e-15, 1.557892e-15, 1.561165e-15, 1.56344e-15, 
    1.562443e-15, 1.567621e-15, 1.56884e-15, 1.573788e-15, 1.571232e-15, 
    1.586433e-15, 1.579715e-15, 1.598333e-15, 1.593139e-15, 1.557928e-15, 
    1.559589e-15, 1.565361e-15, 1.562615e-15, 1.570463e-15, 1.572391e-15, 
    1.573959e-15, 1.575962e-15, 1.576178e-15, 1.577364e-15, 1.575421e-15, 
    1.577288e-15, 1.57022e-15, 1.57338e-15, 1.564702e-15, 1.566816e-15, 
    1.565844e-15, 1.564777e-15, 1.568069e-15, 1.571571e-15, 1.571648e-15, 
    1.572769e-15, 1.575927e-15, 1.570495e-15, 1.587297e-15, 1.576926e-15, 
    1.561398e-15, 1.564591e-15, 1.565049e-15, 1.563812e-15, 1.572198e-15, 
    1.569162e-15, 1.577336e-15, 1.575128e-15, 1.578745e-15, 1.576948e-15, 
    1.576683e-15, 1.574375e-15, 1.572936e-15, 1.569301e-15, 1.56634e-15, 
    1.563991e-15, 1.564538e-15, 1.567117e-15, 1.571786e-15, 1.576197e-15, 
    1.575231e-15, 1.57847e-15, 1.569895e-15, 1.573491e-15, 1.572101e-15, 
    1.575726e-15, 1.567781e-15, 1.574543e-15, 1.56605e-15, 1.566795e-15, 
    1.569101e-15, 1.573734e-15, 1.574761e-15, 1.575854e-15, 1.57518e-15, 
    1.571904e-15, 1.571368e-15, 1.569046e-15, 1.568404e-15, 1.566633e-15, 
    1.565166e-15, 1.566506e-15, 1.567913e-15, 1.571906e-15, 1.5755e-15, 
    1.579417e-15, 1.580375e-15, 1.584941e-15, 1.581222e-15, 1.587354e-15, 
    1.582139e-15, 1.591164e-15, 1.574937e-15, 1.581988e-15, 1.569207e-15, 
    1.570586e-15, 1.573078e-15, 1.578791e-15, 1.575709e-15, 1.579314e-15, 
    1.571347e-15, 1.567206e-15, 1.566135e-15, 1.564134e-15, 1.566181e-15, 
    1.566014e-15, 1.567972e-15, 1.567343e-15, 1.572038e-15, 1.569517e-15, 
    1.576676e-15, 1.579285e-15, 1.586646e-15, 1.59115e-15, 1.595732e-15, 
    1.597752e-15, 1.598367e-15, 1.598624e-15 ;

 LITR3N_vr =
  7.964093e-06, 7.964085e-06, 7.964086e-06, 7.964079e-06, 7.964083e-06, 
    7.964079e-06, 7.964091e-06, 7.964084e-06, 7.964089e-06, 7.964092e-06, 
    7.964067e-06, 7.964079e-06, 7.964053e-06, 7.964061e-06, 7.964041e-06, 
    7.964055e-06, 7.964039e-06, 7.964041e-06, 7.964032e-06, 7.964035e-06, 
    7.964023e-06, 7.96403e-06, 7.964017e-06, 7.964025e-06, 7.964023e-06, 
    7.964031e-06, 7.964077e-06, 7.964068e-06, 7.964077e-06, 7.964076e-06, 
    7.964077e-06, 7.964083e-06, 7.964087e-06, 7.964094e-06, 7.964092e-06, 
    7.964087e-06, 7.964076e-06, 7.964079e-06, 7.964069e-06, 7.964069e-06, 
    7.964059e-06, 7.964063e-06, 7.964045e-06, 7.96405e-06, 7.964035e-06, 
    7.964039e-06, 7.964035e-06, 7.964036e-06, 7.964035e-06, 7.96404e-06, 
    7.964038e-06, 7.964043e-06, 7.964062e-06, 7.964057e-06, 7.964074e-06, 
    7.964084e-06, 7.964091e-06, 7.964096e-06, 7.964095e-06, 7.964094e-06, 
    7.964087e-06, 7.96408e-06, 7.964076e-06, 7.964073e-06, 7.964069e-06, 
    7.96406e-06, 7.964055e-06, 7.964043e-06, 7.964046e-06, 7.964042e-06, 
    7.964039e-06, 7.964033e-06, 7.964034e-06, 7.964031e-06, 7.964042e-06, 
    7.964035e-06, 7.964047e-06, 7.964044e-06, 7.964069e-06, 7.964079e-06, 
    7.964082e-06, 7.964086e-06, 7.964095e-06, 7.964089e-06, 7.964091e-06, 
    7.964085e-06, 7.964082e-06, 7.964084e-06, 7.964073e-06, 7.964077e-06, 
    7.964055e-06, 7.964064e-06, 7.964039e-06, 7.964045e-06, 7.964038e-06, 
    7.964041e-06, 7.964035e-06, 7.964041e-06, 7.96403e-06, 7.964029e-06, 
    7.96403e-06, 7.964024e-06, 7.964041e-06, 7.964035e-06, 7.964084e-06, 
    7.964083e-06, 7.964082e-06, 7.964088e-06, 7.964089e-06, 7.964094e-06, 
    7.964089e-06, 7.964087e-06, 7.964081e-06, 7.964079e-06, 7.964076e-06, 
    7.964069e-06, 7.964062e-06, 7.964052e-06, 7.964045e-06, 7.96404e-06, 
    7.964043e-06, 7.96404e-06, 7.964043e-06, 7.964045e-06, 7.964029e-06, 
    7.964038e-06, 7.964025e-06, 7.964026e-06, 7.964031e-06, 7.964026e-06, 
    7.964083e-06, 7.964085e-06, 7.96409e-06, 7.964086e-06, 7.964094e-06, 
    7.964089e-06, 7.964087e-06, 7.964077e-06, 7.964075e-06, 7.964072e-06, 
    7.964069e-06, 7.964063e-06, 7.964054e-06, 7.964046e-06, 7.964039e-06, 
    7.964039e-06, 7.964039e-06, 7.964038e-06, 7.964041e-06, 7.964037e-06, 
    7.964036e-06, 7.964038e-06, 7.964026e-06, 7.964029e-06, 7.964026e-06, 
    7.964029e-06, 7.964084e-06, 7.964081e-06, 7.964083e-06, 7.96408e-06, 
    7.964082e-06, 7.964073e-06, 7.96407e-06, 7.964059e-06, 7.964063e-06, 
    7.964055e-06, 7.964062e-06, 7.964061e-06, 7.964055e-06, 7.964062e-06, 
    7.964047e-06, 7.964057e-06, 7.964038e-06, 7.964048e-06, 7.964037e-06, 
    7.964039e-06, 7.964035e-06, 7.964032e-06, 7.964029e-06, 7.964021e-06, 
    7.964023e-06, 7.964017e-06, 7.964078e-06, 7.964074e-06, 7.964074e-06, 
    7.96407e-06, 7.964068e-06, 7.964061e-06, 7.964051e-06, 7.964055e-06, 
    7.964049e-06, 7.964048e-06, 7.964058e-06, 7.964051e-06, 7.964071e-06, 
    7.964068e-06, 7.96407e-06, 7.964077e-06, 7.964054e-06, 7.964066e-06, 
    7.964045e-06, 7.964051e-06, 7.964033e-06, 7.964042e-06, 7.964024e-06, 
    7.964017e-06, 7.964009e-06, 7.964001e-06, 7.964071e-06, 7.964074e-06, 
    7.964069e-06, 7.964064e-06, 7.964058e-06, 7.96405e-06, 7.964049e-06, 
    7.964049e-06, 7.964045e-06, 7.964041e-06, 7.964048e-06, 7.964041e-06, 
    7.964068e-06, 7.964053e-06, 7.964075e-06, 7.964069e-06, 7.964064e-06, 
    7.964066e-06, 7.964056e-06, 7.964053e-06, 7.964043e-06, 7.964049e-06, 
    7.964019e-06, 7.964031e-06, 7.963995e-06, 7.964005e-06, 7.964075e-06, 
    7.964071e-06, 7.96406e-06, 7.964066e-06, 7.96405e-06, 7.964046e-06, 
    7.964043e-06, 7.964039e-06, 7.964039e-06, 7.964037e-06, 7.96404e-06, 
    7.964037e-06, 7.96405e-06, 7.964044e-06, 7.964061e-06, 7.964058e-06, 
    7.964059e-06, 7.964061e-06, 7.964055e-06, 7.964048e-06, 7.964048e-06, 
    7.964046e-06, 7.964039e-06, 7.96405e-06, 7.964017e-06, 7.964037e-06, 
    7.964068e-06, 7.964061e-06, 7.96406e-06, 7.964063e-06, 7.964047e-06, 
    7.964052e-06, 7.964037e-06, 7.96404e-06, 7.964033e-06, 7.964037e-06, 
    7.964038e-06, 7.964042e-06, 7.964045e-06, 7.964052e-06, 7.964059e-06, 
    7.964063e-06, 7.964062e-06, 7.964057e-06, 7.964048e-06, 7.964039e-06, 
    7.96404e-06, 7.964034e-06, 7.964051e-06, 7.964044e-06, 7.964047e-06, 
    7.964039e-06, 7.964056e-06, 7.964042e-06, 7.964059e-06, 7.964058e-06, 
    7.964053e-06, 7.964043e-06, 7.964041e-06, 7.964039e-06, 7.96404e-06, 
    7.964047e-06, 7.964049e-06, 7.964053e-06, 7.964054e-06, 7.964058e-06, 
    7.96406e-06, 7.964058e-06, 7.964055e-06, 7.964047e-06, 7.96404e-06, 
    7.964032e-06, 7.96403e-06, 7.964021e-06, 7.964029e-06, 7.964017e-06, 
    7.964027e-06, 7.964009e-06, 7.964041e-06, 7.964027e-06, 7.964052e-06, 
    7.964049e-06, 7.964045e-06, 7.964033e-06, 7.964039e-06, 7.964032e-06, 
    7.964049e-06, 7.964057e-06, 7.964059e-06, 7.964062e-06, 7.964059e-06, 
    7.964059e-06, 7.964055e-06, 7.964056e-06, 7.964047e-06, 7.964052e-06, 
    7.964038e-06, 7.964032e-06, 7.964018e-06, 7.964009e-06, 7.963999e-06, 
    7.963996e-06, 7.963995e-06, 7.963994e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3_HR =
  5.596049e-14, 5.611208e-14, 5.608263e-14, 5.620478e-14, 5.613705e-14, 
    5.621701e-14, 5.599125e-14, 5.611807e-14, 5.603714e-14, 5.597417e-14, 
    5.644149e-14, 5.621023e-14, 5.668151e-14, 5.653429e-14, 5.690388e-14, 
    5.665858e-14, 5.69533e-14, 5.689685e-14, 5.706679e-14, 5.701813e-14, 
    5.723516e-14, 5.708924e-14, 5.734761e-14, 5.720035e-14, 5.722338e-14, 
    5.708442e-14, 5.625685e-14, 5.641271e-14, 5.62476e-14, 5.626984e-14, 
    5.625987e-14, 5.613843e-14, 5.607717e-14, 5.594892e-14, 5.597223e-14, 
    5.606643e-14, 5.627984e-14, 5.620746e-14, 5.63899e-14, 5.638578e-14, 
    5.658858e-14, 5.649718e-14, 5.683761e-14, 5.674098e-14, 5.702016e-14, 
    5.694998e-14, 5.701686e-14, 5.699659e-14, 5.701712e-14, 5.691419e-14, 
    5.69583e-14, 5.68677e-14, 5.651429e-14, 5.661824e-14, 5.630796e-14, 
    5.6121e-14, 5.599681e-14, 5.590858e-14, 5.592106e-14, 5.594483e-14, 
    5.606698e-14, 5.618178e-14, 5.626919e-14, 5.632763e-14, 5.638519e-14, 
    5.655915e-14, 5.665125e-14, 5.685713e-14, 5.682003e-14, 5.68829e-14, 
    5.6943e-14, 5.704379e-14, 5.702721e-14, 5.707159e-14, 5.688128e-14, 
    5.700777e-14, 5.679889e-14, 5.685604e-14, 5.640067e-14, 5.6227e-14, 
    5.615298e-14, 5.608829e-14, 5.593065e-14, 5.603952e-14, 5.599661e-14, 
    5.609871e-14, 5.616353e-14, 5.613148e-14, 5.632922e-14, 5.625237e-14, 
    5.66567e-14, 5.648269e-14, 5.6936e-14, 5.682765e-14, 5.696196e-14, 
    5.689345e-14, 5.70108e-14, 5.690519e-14, 5.708811e-14, 5.712789e-14, 
    5.710071e-14, 5.720517e-14, 5.689933e-14, 5.701684e-14, 5.613057e-14, 
    5.61358e-14, 5.616017e-14, 5.605303e-14, 5.604648e-14, 5.594828e-14, 
    5.603568e-14, 5.607287e-14, 5.61673e-14, 5.62231e-14, 5.627613e-14, 
    5.639267e-14, 5.652267e-14, 5.670432e-14, 5.683468e-14, 5.6922e-14, 
    5.686847e-14, 5.691573e-14, 5.686289e-14, 5.683813e-14, 5.711298e-14, 
    5.69587e-14, 5.719015e-14, 5.717736e-14, 5.707263e-14, 5.71788e-14, 
    5.613947e-14, 5.610939e-14, 5.600485e-14, 5.608667e-14, 5.593758e-14, 
    5.602103e-14, 5.606898e-14, 5.625394e-14, 5.629459e-14, 5.633222e-14, 
    5.640655e-14, 5.650186e-14, 5.666889e-14, 5.681406e-14, 5.694651e-14, 
    5.693681e-14, 5.694022e-14, 5.696978e-14, 5.689653e-14, 5.69818e-14, 
    5.699609e-14, 5.69587e-14, 5.717565e-14, 5.71137e-14, 5.717708e-14, 
    5.713676e-14, 5.611918e-14, 5.616979e-14, 5.614244e-14, 5.619386e-14, 
    5.615762e-14, 5.631865e-14, 5.636689e-14, 5.659246e-14, 5.649997e-14, 
    5.664719e-14, 5.651495e-14, 5.653838e-14, 5.665192e-14, 5.652211e-14, 
    5.680603e-14, 5.661355e-14, 5.697093e-14, 5.677887e-14, 5.698295e-14, 
    5.694594e-14, 5.700724e-14, 5.706209e-14, 5.713111e-14, 5.725832e-14, 
    5.722887e-14, 5.733521e-14, 5.624524e-14, 5.631082e-14, 5.630508e-14, 
    5.63737e-14, 5.642443e-14, 5.653434e-14, 5.671042e-14, 5.664424e-14, 
    5.676575e-14, 5.679009e-14, 5.660553e-14, 5.671886e-14, 5.635472e-14, 
    5.641358e-14, 5.637856e-14, 5.625039e-14, 5.665945e-14, 5.644965e-14, 
    5.683683e-14, 5.672338e-14, 5.705427e-14, 5.688976e-14, 5.721266e-14, 
    5.735039e-14, 5.748002e-14, 5.763119e-14, 5.634663e-14, 5.630208e-14, 
    5.638187e-14, 5.649213e-14, 5.659444e-14, 5.67303e-14, 5.674421e-14, 
    5.676964e-14, 5.683549e-14, 5.689084e-14, 5.677765e-14, 5.690471e-14, 
    5.642717e-14, 5.667766e-14, 5.628521e-14, 5.640346e-14, 5.648565e-14, 
    5.644963e-14, 5.663669e-14, 5.668073e-14, 5.685951e-14, 5.676715e-14, 
    5.731637e-14, 5.707363e-14, 5.774629e-14, 5.755863e-14, 5.62865e-14, 
    5.63465e-14, 5.655503e-14, 5.645585e-14, 5.673939e-14, 5.680905e-14, 
    5.68657e-14, 5.693804e-14, 5.694587e-14, 5.698872e-14, 5.691849e-14, 
    5.698595e-14, 5.673059e-14, 5.684475e-14, 5.653125e-14, 5.66076e-14, 
    5.65725e-14, 5.653395e-14, 5.665288e-14, 5.677942e-14, 5.678217e-14, 
    5.682269e-14, 5.693678e-14, 5.674053e-14, 5.734758e-14, 5.697289e-14, 
    5.641188e-14, 5.652723e-14, 5.654376e-14, 5.649908e-14, 5.680206e-14, 
    5.669237e-14, 5.698768e-14, 5.690793e-14, 5.703858e-14, 5.697367e-14, 
    5.696411e-14, 5.68807e-14, 5.682873e-14, 5.669739e-14, 5.659042e-14, 
    5.650557e-14, 5.652531e-14, 5.66185e-14, 5.678717e-14, 5.694655e-14, 
    5.691164e-14, 5.702866e-14, 5.671884e-14, 5.684879e-14, 5.679855e-14, 
    5.692952e-14, 5.664248e-14, 5.688679e-14, 5.657993e-14, 5.660688e-14, 
    5.669019e-14, 5.685757e-14, 5.689466e-14, 5.693416e-14, 5.69098e-14, 
    5.679143e-14, 5.677208e-14, 5.668817e-14, 5.666498e-14, 5.660101e-14, 
    5.654801e-14, 5.659643e-14, 5.664724e-14, 5.67915e-14, 5.692138e-14, 
    5.706287e-14, 5.709749e-14, 5.726245e-14, 5.712811e-14, 5.734965e-14, 
    5.716121e-14, 5.748731e-14, 5.690101e-14, 5.715577e-14, 5.6694e-14, 
    5.674383e-14, 5.683384e-14, 5.704026e-14, 5.692891e-14, 5.705914e-14, 
    5.677133e-14, 5.662169e-14, 5.658301e-14, 5.651072e-14, 5.658467e-14, 
    5.657866e-14, 5.664938e-14, 5.662666e-14, 5.679629e-14, 5.670521e-14, 
    5.696386e-14, 5.705812e-14, 5.732406e-14, 5.748679e-14, 5.765233e-14, 
    5.772532e-14, 5.774753e-14, 5.775681e-14 ;

 LITTERC =
  6.210311e-05, 6.210295e-05, 6.210298e-05, 6.210285e-05, 6.210292e-05, 
    6.210284e-05, 6.210307e-05, 6.210294e-05, 6.210303e-05, 6.210309e-05, 
    6.21026e-05, 6.210284e-05, 6.210235e-05, 6.21025e-05, 6.210212e-05, 
    6.210238e-05, 6.210207e-05, 6.210212e-05, 6.210195e-05, 6.2102e-05, 
    6.210178e-05, 6.210193e-05, 6.210166e-05, 6.210181e-05, 6.210179e-05, 
    6.210194e-05, 6.210279e-05, 6.210263e-05, 6.21028e-05, 6.210278e-05, 
    6.210279e-05, 6.210292e-05, 6.210298e-05, 6.210311e-05, 6.210309e-05, 
    6.210299e-05, 6.210277e-05, 6.210284e-05, 6.210266e-05, 6.210266e-05, 
    6.210245e-05, 6.210255e-05, 6.210219e-05, 6.210229e-05, 6.2102e-05, 
    6.210207e-05, 6.2102e-05, 6.210202e-05, 6.2102e-05, 6.210211e-05, 
    6.210207e-05, 6.210216e-05, 6.210252e-05, 6.210242e-05, 6.210274e-05, 
    6.210294e-05, 6.210306e-05, 6.210316e-05, 6.210314e-05, 6.210312e-05, 
    6.210299e-05, 6.210287e-05, 6.210278e-05, 6.210272e-05, 6.210266e-05, 
    6.210248e-05, 6.210239e-05, 6.210217e-05, 6.21022e-05, 6.210214e-05, 
    6.210208e-05, 6.210197e-05, 6.210199e-05, 6.210194e-05, 6.210215e-05, 
    6.210202e-05, 6.210223e-05, 6.210217e-05, 6.210264e-05, 6.210282e-05, 
    6.21029e-05, 6.210297e-05, 6.210314e-05, 6.210302e-05, 6.210306e-05, 
    6.210296e-05, 6.210289e-05, 6.210292e-05, 6.210272e-05, 6.21028e-05, 
    6.210238e-05, 6.210256e-05, 6.210209e-05, 6.21022e-05, 6.210206e-05, 
    6.210213e-05, 6.210201e-05, 6.210212e-05, 6.210193e-05, 6.210188e-05, 
    6.210191e-05, 6.21018e-05, 6.210212e-05, 6.2102e-05, 6.210292e-05, 
    6.210292e-05, 6.21029e-05, 6.2103e-05, 6.210301e-05, 6.210311e-05, 
    6.210303e-05, 6.210298e-05, 6.210289e-05, 6.210283e-05, 6.210277e-05, 
    6.210266e-05, 6.210252e-05, 6.210233e-05, 6.210219e-05, 6.21021e-05, 
    6.210215e-05, 6.210211e-05, 6.210216e-05, 6.210219e-05, 6.21019e-05, 
    6.210207e-05, 6.210182e-05, 6.210183e-05, 6.210194e-05, 6.210183e-05, 
    6.210292e-05, 6.210295e-05, 6.210306e-05, 6.210297e-05, 6.210313e-05, 
    6.210304e-05, 6.210299e-05, 6.210279e-05, 6.210276e-05, 6.210271e-05, 
    6.210264e-05, 6.210254e-05, 6.210236e-05, 6.210221e-05, 6.210207e-05, 
    6.210209e-05, 6.210208e-05, 6.210205e-05, 6.210212e-05, 6.210204e-05, 
    6.210202e-05, 6.210207e-05, 6.210183e-05, 6.21019e-05, 6.210183e-05, 
    6.210188e-05, 6.210294e-05, 6.210289e-05, 6.210291e-05, 6.210286e-05, 
    6.21029e-05, 6.210273e-05, 6.210268e-05, 6.210244e-05, 6.210254e-05, 
    6.210239e-05, 6.210252e-05, 6.21025e-05, 6.210238e-05, 6.210252e-05, 
    6.210222e-05, 6.210242e-05, 6.210205e-05, 6.210225e-05, 6.210204e-05, 
    6.210207e-05, 6.210202e-05, 6.210196e-05, 6.210188e-05, 6.210175e-05, 
    6.210178e-05, 6.210167e-05, 6.210281e-05, 6.210274e-05, 6.210274e-05, 
    6.210267e-05, 6.210262e-05, 6.21025e-05, 6.210232e-05, 6.210239e-05, 
    6.210226e-05, 6.210224e-05, 6.210243e-05, 6.210231e-05, 6.210269e-05, 
    6.210263e-05, 6.210267e-05, 6.21028e-05, 6.210237e-05, 6.210259e-05, 
    6.210219e-05, 6.210231e-05, 6.210196e-05, 6.210213e-05, 6.21018e-05, 
    6.210165e-05, 6.210152e-05, 6.210136e-05, 6.21027e-05, 6.210275e-05, 
    6.210266e-05, 6.210255e-05, 6.210244e-05, 6.21023e-05, 6.210228e-05, 
    6.210226e-05, 6.210219e-05, 6.210213e-05, 6.210225e-05, 6.210212e-05, 
    6.210262e-05, 6.210236e-05, 6.210276e-05, 6.210264e-05, 6.210255e-05, 
    6.210259e-05, 6.21024e-05, 6.210235e-05, 6.210217e-05, 6.210226e-05, 
    6.210169e-05, 6.210194e-05, 6.210124e-05, 6.210144e-05, 6.210276e-05, 
    6.21027e-05, 6.210248e-05, 6.210259e-05, 6.210229e-05, 6.210222e-05, 
    6.210216e-05, 6.210208e-05, 6.210207e-05, 6.210203e-05, 6.21021e-05, 
    6.210204e-05, 6.21023e-05, 6.210218e-05, 6.210251e-05, 6.210243e-05, 
    6.210247e-05, 6.21025e-05, 6.210238e-05, 6.210225e-05, 6.210225e-05, 
    6.21022e-05, 6.210209e-05, 6.210229e-05, 6.210166e-05, 6.210204e-05, 
    6.210263e-05, 6.210251e-05, 6.21025e-05, 6.210254e-05, 6.210223e-05, 
    6.210234e-05, 6.210203e-05, 6.210212e-05, 6.210198e-05, 6.210204e-05, 
    6.210206e-05, 6.210215e-05, 6.21022e-05, 6.210234e-05, 6.210244e-05, 
    6.210253e-05, 6.210252e-05, 6.210242e-05, 6.210224e-05, 6.210207e-05, 
    6.210211e-05, 6.210199e-05, 6.210231e-05, 6.210218e-05, 6.210223e-05, 
    6.21021e-05, 6.210239e-05, 6.210214e-05, 6.210246e-05, 6.210243e-05, 
    6.210234e-05, 6.210217e-05, 6.210213e-05, 6.210209e-05, 6.210212e-05, 
    6.210223e-05, 6.210226e-05, 6.210234e-05, 6.210237e-05, 6.210244e-05, 
    6.210249e-05, 6.210244e-05, 6.210239e-05, 6.210223e-05, 6.21021e-05, 
    6.210196e-05, 6.210192e-05, 6.210175e-05, 6.210188e-05, 6.210166e-05, 
    6.210186e-05, 6.210151e-05, 6.210212e-05, 6.210186e-05, 6.210234e-05, 
    6.210228e-05, 6.210219e-05, 6.210198e-05, 6.21021e-05, 6.210196e-05, 
    6.210226e-05, 6.210242e-05, 6.210245e-05, 6.210253e-05, 6.210245e-05, 
    6.210246e-05, 6.210239e-05, 6.210241e-05, 6.210223e-05, 6.210233e-05, 
    6.210206e-05, 6.210196e-05, 6.210168e-05, 6.210151e-05, 6.210134e-05, 
    6.210127e-05, 6.210124e-05, 6.210123e-05 ;

 LITTERC_HR =
  9.028442e-13, 9.052879e-13, 9.048132e-13, 9.067824e-13, 9.056906e-13, 
    9.069795e-13, 9.033402e-13, 9.053846e-13, 9.040799e-13, 9.030648e-13, 
    9.105982e-13, 9.068703e-13, 9.144674e-13, 9.120941e-13, 9.180519e-13, 
    9.140977e-13, 9.188485e-13, 9.179387e-13, 9.20678e-13, 9.198936e-13, 
    9.233922e-13, 9.2104e-13, 9.252049e-13, 9.22831e-13, 9.232023e-13, 
    9.209622e-13, 9.076217e-13, 9.101342e-13, 9.074726e-13, 9.078311e-13, 
    9.076704e-13, 9.057128e-13, 9.047252e-13, 9.026579e-13, 9.030335e-13, 
    9.045521e-13, 9.079923e-13, 9.068256e-13, 9.097664e-13, 9.097e-13, 
    9.129694e-13, 9.114959e-13, 9.169837e-13, 9.154259e-13, 9.199265e-13, 
    9.187952e-13, 9.198731e-13, 9.195464e-13, 9.198775e-13, 9.182181e-13, 
    9.189291e-13, 9.174688e-13, 9.117717e-13, 9.134475e-13, 9.084456e-13, 
    9.054318e-13, 9.034297e-13, 9.020075e-13, 9.022086e-13, 9.025918e-13, 
    9.045609e-13, 9.064116e-13, 9.078206e-13, 9.087626e-13, 9.096905e-13, 
    9.124949e-13, 9.139795e-13, 9.172984e-13, 9.167003e-13, 9.177138e-13, 
    9.186827e-13, 9.203073e-13, 9.200401e-13, 9.207554e-13, 9.176876e-13, 
    9.197266e-13, 9.163595e-13, 9.172809e-13, 9.099401e-13, 9.071405e-13, 
    9.059473e-13, 9.049044e-13, 9.023632e-13, 9.041183e-13, 9.034265e-13, 
    9.050725e-13, 9.061174e-13, 9.056007e-13, 9.087884e-13, 9.075495e-13, 
    9.140674e-13, 9.112623e-13, 9.185697e-13, 9.168231e-13, 9.189882e-13, 
    9.178838e-13, 9.197755e-13, 9.180731e-13, 9.210217e-13, 9.21663e-13, 
    9.212248e-13, 9.229087e-13, 9.179786e-13, 9.198729e-13, 9.055861e-13, 
    9.056703e-13, 9.060631e-13, 9.043361e-13, 9.042305e-13, 9.026474e-13, 
    9.040563e-13, 9.046559e-13, 9.061781e-13, 9.070776e-13, 9.079325e-13, 
    9.098111e-13, 9.119069e-13, 9.14835e-13, 9.169363e-13, 9.183441e-13, 
    9.174812e-13, 9.18243e-13, 9.173913e-13, 9.169921e-13, 9.214226e-13, 
    9.189356e-13, 9.226666e-13, 9.224604e-13, 9.207722e-13, 9.224837e-13, 
    9.057296e-13, 9.052446e-13, 9.035593e-13, 9.048783e-13, 9.02475e-13, 
    9.038203e-13, 9.045932e-13, 9.075749e-13, 9.082301e-13, 9.088366e-13, 
    9.100349e-13, 9.115713e-13, 9.142639e-13, 9.16604e-13, 9.187392e-13, 
    9.185828e-13, 9.186378e-13, 9.191142e-13, 9.179335e-13, 9.19308e-13, 
    9.195383e-13, 9.189356e-13, 9.224327e-13, 9.214343e-13, 9.22456e-13, 
    9.218059e-13, 9.054023e-13, 9.062184e-13, 9.057774e-13, 9.066063e-13, 
    9.060222e-13, 9.086179e-13, 9.093956e-13, 9.130319e-13, 9.115409e-13, 
    9.13914e-13, 9.117823e-13, 9.1216e-13, 9.139903e-13, 9.118977e-13, 
    9.164746e-13, 9.133717e-13, 9.191327e-13, 9.160368e-13, 9.193266e-13, 
    9.187298e-13, 9.19718e-13, 9.206024e-13, 9.217149e-13, 9.237654e-13, 
    9.232908e-13, 9.250051e-13, 9.074346e-13, 9.084918e-13, 9.083992e-13, 
    9.095054e-13, 9.103231e-13, 9.120951e-13, 9.149334e-13, 9.138666e-13, 
    9.158252e-13, 9.162176e-13, 9.132426e-13, 9.150695e-13, 9.091994e-13, 
    9.101483e-13, 9.095837e-13, 9.075177e-13, 9.141118e-13, 9.107297e-13, 
    9.16971e-13, 9.151424e-13, 9.204762e-13, 9.178244e-13, 9.230294e-13, 
    9.252496e-13, 9.273394e-13, 9.297761e-13, 9.09069e-13, 9.083509e-13, 
    9.096371e-13, 9.114145e-13, 9.130638e-13, 9.152539e-13, 9.154781e-13, 
    9.15888e-13, 9.169495e-13, 9.178416e-13, 9.16017e-13, 9.180653e-13, 
    9.103673e-13, 9.144054e-13, 9.080788e-13, 9.099851e-13, 9.1131e-13, 
    9.107294e-13, 9.137448e-13, 9.144547e-13, 9.173367e-13, 9.158479e-13, 
    9.247014e-13, 9.207883e-13, 9.316315e-13, 9.286064e-13, 9.080998e-13, 
    9.090668e-13, 9.124286e-13, 9.108298e-13, 9.154002e-13, 9.165232e-13, 
    9.174365e-13, 9.186025e-13, 9.187289e-13, 9.194195e-13, 9.182876e-13, 
    9.193749e-13, 9.152585e-13, 9.170989e-13, 9.120451e-13, 9.13276e-13, 
    9.1271e-13, 9.120887e-13, 9.140057e-13, 9.160457e-13, 9.160901e-13, 
    9.167431e-13, 9.185824e-13, 9.154188e-13, 9.252044e-13, 9.191644e-13, 
    9.101208e-13, 9.119803e-13, 9.122468e-13, 9.115266e-13, 9.164106e-13, 
    9.146423e-13, 9.194028e-13, 9.181171e-13, 9.202234e-13, 9.19177e-13, 
    9.190229e-13, 9.176784e-13, 9.168406e-13, 9.147233e-13, 9.12999e-13, 
    9.116311e-13, 9.119493e-13, 9.134516e-13, 9.161706e-13, 9.187399e-13, 
    9.181771e-13, 9.200634e-13, 9.150691e-13, 9.171639e-13, 9.163541e-13, 
    9.184654e-13, 9.13838e-13, 9.177765e-13, 9.128299e-13, 9.132643e-13, 
    9.146073e-13, 9.173055e-13, 9.179033e-13, 9.1854e-13, 9.181473e-13, 
    9.162392e-13, 9.159274e-13, 9.145747e-13, 9.142008e-13, 9.131697e-13, 
    9.123154e-13, 9.130958e-13, 9.139149e-13, 9.162404e-13, 9.18334e-13, 
    9.206148e-13, 9.211729e-13, 9.238321e-13, 9.216665e-13, 9.252378e-13, 
    9.222001e-13, 9.274567e-13, 9.180057e-13, 9.221124e-13, 9.146686e-13, 
    9.154719e-13, 9.169229e-13, 9.202503e-13, 9.184554e-13, 9.205548e-13, 
    9.159151e-13, 9.135031e-13, 9.128796e-13, 9.117142e-13, 9.129063e-13, 
    9.128093e-13, 9.139494e-13, 9.135831e-13, 9.163176e-13, 9.148495e-13, 
    9.190188e-13, 9.205384e-13, 9.248251e-13, 9.274484e-13, 9.301169e-13, 
    9.312933e-13, 9.316515e-13, 9.318011e-13 ;

 LITTERC_LOSS =
  1.672059e-12, 1.676585e-12, 1.675705e-12, 1.679352e-12, 1.67733e-12, 
    1.679717e-12, 1.672977e-12, 1.676764e-12, 1.674347e-12, 1.672467e-12, 
    1.686419e-12, 1.679515e-12, 1.693585e-12, 1.68919e-12, 1.700224e-12, 
    1.692901e-12, 1.701699e-12, 1.700014e-12, 1.705087e-12, 1.703635e-12, 
    1.710114e-12, 1.705758e-12, 1.713471e-12, 1.709075e-12, 1.709762e-12, 
    1.705614e-12, 1.680907e-12, 1.68556e-12, 1.680631e-12, 1.681295e-12, 
    1.680997e-12, 1.677372e-12, 1.675543e-12, 1.671714e-12, 1.672409e-12, 
    1.675222e-12, 1.681593e-12, 1.679432e-12, 1.684879e-12, 1.684756e-12, 
    1.690811e-12, 1.688082e-12, 1.698246e-12, 1.69536e-12, 1.703695e-12, 
    1.7016e-12, 1.703597e-12, 1.702992e-12, 1.703605e-12, 1.700532e-12, 
    1.701848e-12, 1.699144e-12, 1.688593e-12, 1.691696e-12, 1.682433e-12, 
    1.676851e-12, 1.673143e-12, 1.670509e-12, 1.670882e-12, 1.671591e-12, 
    1.675238e-12, 1.678666e-12, 1.681275e-12, 1.68302e-12, 1.684738e-12, 
    1.689932e-12, 1.692682e-12, 1.698828e-12, 1.697721e-12, 1.699598e-12, 
    1.701392e-12, 1.704401e-12, 1.703906e-12, 1.705231e-12, 1.699549e-12, 
    1.703326e-12, 1.697089e-12, 1.698796e-12, 1.685201e-12, 1.680016e-12, 
    1.677806e-12, 1.675874e-12, 1.671168e-12, 1.674418e-12, 1.673137e-12, 
    1.676186e-12, 1.678121e-12, 1.677164e-12, 1.683068e-12, 1.680773e-12, 
    1.692845e-12, 1.687649e-12, 1.701183e-12, 1.697948e-12, 1.701958e-12, 
    1.699912e-12, 1.703416e-12, 1.700263e-12, 1.705724e-12, 1.706912e-12, 
    1.7061e-12, 1.709219e-12, 1.700088e-12, 1.703596e-12, 1.677137e-12, 
    1.677293e-12, 1.67802e-12, 1.674822e-12, 1.674626e-12, 1.671694e-12, 
    1.674304e-12, 1.675414e-12, 1.678233e-12, 1.679899e-12, 1.681482e-12, 
    1.684962e-12, 1.688843e-12, 1.694266e-12, 1.698158e-12, 1.700765e-12, 
    1.699167e-12, 1.700578e-12, 1.699e-12, 1.698261e-12, 1.706466e-12, 
    1.70186e-12, 1.70877e-12, 1.708388e-12, 1.705262e-12, 1.708431e-12, 
    1.677403e-12, 1.676504e-12, 1.673383e-12, 1.675826e-12, 1.671375e-12, 
    1.673866e-12, 1.675298e-12, 1.68082e-12, 1.682034e-12, 1.683157e-12, 
    1.685376e-12, 1.688222e-12, 1.693208e-12, 1.697542e-12, 1.701496e-12, 
    1.701207e-12, 1.701309e-12, 1.702191e-12, 1.700005e-12, 1.70255e-12, 
    1.702977e-12, 1.70186e-12, 1.708337e-12, 1.706488e-12, 1.70838e-12, 
    1.707176e-12, 1.676797e-12, 1.678308e-12, 1.677491e-12, 1.679026e-12, 
    1.677944e-12, 1.682752e-12, 1.684192e-12, 1.690927e-12, 1.688165e-12, 
    1.69256e-12, 1.688612e-12, 1.689312e-12, 1.692702e-12, 1.688826e-12, 
    1.697303e-12, 1.691556e-12, 1.702225e-12, 1.696492e-12, 1.702584e-12, 
    1.701479e-12, 1.703309e-12, 1.704947e-12, 1.707008e-12, 1.710805e-12, 
    1.709926e-12, 1.713101e-12, 1.68056e-12, 1.682518e-12, 1.682347e-12, 
    1.684395e-12, 1.68591e-12, 1.689191e-12, 1.694448e-12, 1.692473e-12, 
    1.6961e-12, 1.696827e-12, 1.691317e-12, 1.6947e-12, 1.683829e-12, 
    1.685586e-12, 1.684541e-12, 1.680714e-12, 1.692927e-12, 1.686663e-12, 
    1.698222e-12, 1.694835e-12, 1.704714e-12, 1.699802e-12, 1.709442e-12, 
    1.713554e-12, 1.717424e-12, 1.721937e-12, 1.683587e-12, 1.682257e-12, 
    1.684639e-12, 1.687931e-12, 1.690986e-12, 1.695042e-12, 1.695457e-12, 
    1.696216e-12, 1.698182e-12, 1.699834e-12, 1.696455e-12, 1.700249e-12, 
    1.685992e-12, 1.69347e-12, 1.681753e-12, 1.685284e-12, 1.687738e-12, 
    1.686662e-12, 1.692247e-12, 1.693562e-12, 1.698899e-12, 1.696142e-12, 
    1.712539e-12, 1.705292e-12, 1.725373e-12, 1.719771e-12, 1.681792e-12, 
    1.683583e-12, 1.689809e-12, 1.686848e-12, 1.695313e-12, 1.697393e-12, 
    1.699084e-12, 1.701244e-12, 1.701477e-12, 1.702757e-12, 1.70066e-12, 
    1.702674e-12, 1.69505e-12, 1.698459e-12, 1.689099e-12, 1.691379e-12, 
    1.69033e-12, 1.68918e-12, 1.69273e-12, 1.696508e-12, 1.69659e-12, 
    1.6978e-12, 1.701206e-12, 1.695347e-12, 1.71347e-12, 1.702284e-12, 
    1.685535e-12, 1.688979e-12, 1.689473e-12, 1.688139e-12, 1.697184e-12, 
    1.693909e-12, 1.702726e-12, 1.700345e-12, 1.704245e-12, 1.702307e-12, 
    1.702022e-12, 1.699532e-12, 1.69798e-12, 1.694059e-12, 1.690866e-12, 
    1.688332e-12, 1.688922e-12, 1.691704e-12, 1.69674e-12, 1.701498e-12, 
    1.700456e-12, 1.703949e-12, 1.6947e-12, 1.698579e-12, 1.697079e-12, 
    1.70099e-12, 1.69242e-12, 1.699714e-12, 1.690552e-12, 1.691357e-12, 
    1.693844e-12, 1.698841e-12, 1.699949e-12, 1.701128e-12, 1.7004e-12, 
    1.696867e-12, 1.696289e-12, 1.693784e-12, 1.693091e-12, 1.691182e-12, 
    1.6896e-12, 1.691045e-12, 1.692562e-12, 1.696869e-12, 1.700746e-12, 
    1.70497e-12, 1.706004e-12, 1.710929e-12, 1.706918e-12, 1.713532e-12, 
    1.707906e-12, 1.717642e-12, 1.700138e-12, 1.707744e-12, 1.693958e-12, 
    1.695446e-12, 1.698133e-12, 1.704295e-12, 1.700971e-12, 1.704859e-12, 
    1.696266e-12, 1.691799e-12, 1.690644e-12, 1.688486e-12, 1.690694e-12, 
    1.690514e-12, 1.692626e-12, 1.691947e-12, 1.697012e-12, 1.694293e-12, 
    1.702015e-12, 1.704829e-12, 1.712768e-12, 1.717626e-12, 1.722568e-12, 
    1.724747e-12, 1.72541e-12, 1.725687e-12 ;

 LIVECROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVECROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 MEG_acetaldehyde =
  4.222116e-18, 4.220624e-18, 4.220907e-18, 4.21972e-18, 4.220368e-18, 
    4.219599e-18, 4.221801e-18, 4.220576e-18, 4.221351e-18, 4.221965e-18, 
    4.217458e-18, 4.219664e-18, 4.215054e-18, 4.216476e-18, 4.212871e-18, 
    4.215291e-18, 4.212378e-18, 4.212912e-18, 4.211238e-18, 4.211715e-18, 
    4.209636e-18, 4.211017e-18, 4.208515e-18, 4.20995e-18, 4.209736e-18, 
    4.211067e-18, 4.219193e-18, 4.217741e-18, 4.219285e-18, 4.219076e-18, 
    4.219164e-18, 4.220364e-18, 4.220989e-18, 4.222212e-18, 4.221984e-18, 
    4.221076e-18, 4.218982e-18, 4.219674e-18, 4.217877e-18, 4.217917e-18, 
    4.21594e-18, 4.216832e-18, 4.213494e-18, 4.214435e-18, 4.211695e-18, 
    4.212387e-18, 4.211732e-18, 4.211927e-18, 4.21173e-18, 4.212744e-18, 
    4.212311e-18, 4.213194e-18, 4.21667e-18, 4.215657e-18, 4.218698e-18, 
    4.220574e-18, 4.221752e-18, 4.222611e-18, 4.22249e-18, 4.222264e-18, 
    4.221071e-18, 4.219926e-18, 4.219063e-18, 4.218491e-18, 4.217923e-18, 
    4.21628e-18, 4.21535e-18, 4.213317e-18, 4.21366e-18, 4.213061e-18, 
    4.212455e-18, 4.211471e-18, 4.211629e-18, 4.211202e-18, 4.213059e-18, 
    4.211833e-18, 4.213861e-18, 4.213309e-18, 4.217864e-18, 4.219482e-18, 
    4.220254e-18, 4.220857e-18, 4.222398e-18, 4.221339e-18, 4.221759e-18, 
    4.22074e-18, 4.220107e-18, 4.220416e-18, 4.218475e-18, 4.219232e-18, 
    4.215295e-18, 4.216988e-18, 4.212526e-18, 4.213588e-18, 4.212268e-18, 
    4.212936e-18, 4.211799e-18, 4.212822e-18, 4.211035e-18, 4.210657e-18, 
    4.210917e-18, 4.209887e-18, 4.212881e-18, 4.211741e-18, 4.220429e-18, 
    4.220379e-18, 4.220136e-18, 4.221207e-18, 4.221268e-18, 4.222222e-18, 
    4.221364e-18, 4.221007e-18, 4.220062e-18, 4.219522e-18, 4.219002e-18, 
    4.217859e-18, 4.2166e-18, 4.214816e-18, 4.21352e-18, 4.212657e-18, 
    4.21318e-18, 4.212719e-18, 4.213237e-18, 4.213476e-18, 4.210805e-18, 
    4.212312e-18, 4.210035e-18, 4.210157e-18, 4.211195e-18, 4.210143e-18, 
    4.220342e-18, 4.220632e-18, 4.22167e-18, 4.220858e-18, 4.222325e-18, 
    4.221515e-18, 4.221057e-18, 4.219238e-18, 4.218815e-18, 4.218454e-18, 
    4.217718e-18, 4.216786e-18, 4.21516e-18, 4.213732e-18, 4.212416e-18, 
    4.212511e-18, 4.212478e-18, 4.212194e-18, 4.21291e-18, 4.212076e-18, 
    4.211945e-18, 4.212301e-18, 4.210174e-18, 4.21078e-18, 4.21016e-18, 
    4.210552e-18, 4.220536e-18, 4.220043e-18, 4.220311e-18, 4.219814e-18, 
    4.220171e-18, 4.218608e-18, 4.21814e-18, 4.215926e-18, 4.21681e-18, 
    4.215377e-18, 4.216657e-18, 4.216435e-18, 4.21537e-18, 4.216581e-18, 
    4.213828e-18, 4.21573e-18, 4.212183e-18, 4.214116e-18, 4.212064e-18, 
    4.212422e-18, 4.21182e-18, 4.211292e-18, 4.210611e-18, 4.209383e-18, 
    4.209663e-18, 4.208622e-18, 4.219301e-18, 4.218673e-18, 4.21871e-18, 
    4.21804e-18, 4.21755e-18, 4.216463e-18, 4.214745e-18, 4.215385e-18, 
    4.21419e-18, 4.213956e-18, 4.215761e-18, 4.21467e-18, 4.218239e-18, 
    4.21768e-18, 4.217999e-18, 4.219262e-18, 4.215262e-18, 4.217324e-18, 
    4.213502e-18, 4.214613e-18, 4.21137e-18, 4.213e-18, 4.209822e-18, 
    4.208513e-18, 4.2072e-18, 4.205763e-18, 4.218311e-18, 4.218739e-18, 
    4.217956e-18, 4.216906e-18, 4.215881e-18, 4.214549e-18, 4.214403e-18, 
    4.214158e-18, 4.213504e-18, 4.212964e-18, 4.214099e-18, 4.212826e-18, 
    4.217586e-18, 4.215075e-18, 4.218918e-18, 4.217784e-18, 4.216959e-18, 
    4.217303e-18, 4.215453e-18, 4.215025e-18, 4.213289e-18, 4.214175e-18, 
    4.208851e-18, 4.211206e-18, 4.204613e-18, 4.206462e-18, 4.218894e-18, 
    4.218303e-18, 4.216279e-18, 4.217239e-18, 4.21445e-18, 4.213773e-18, 
    4.213207e-18, 4.212513e-18, 4.212425e-18, 4.212012e-18, 4.212691e-18, 
    4.212032e-18, 4.214546e-18, 4.213419e-18, 4.216489e-18, 4.215751e-18, 
    4.216084e-18, 4.216463e-18, 4.215297e-18, 4.214085e-18, 4.214031e-18, 
    4.213647e-18, 4.212619e-18, 4.214438e-18, 4.2086e-18, 4.212251e-18, 
    4.217662e-18, 4.216567e-18, 4.216376e-18, 4.216806e-18, 4.213841e-18, 
    4.214918e-18, 4.212019e-18, 4.212795e-18, 4.211515e-18, 4.212153e-18, 
    4.212249e-18, 4.213062e-18, 4.213577e-18, 4.214874e-18, 4.215923e-18, 
    4.21674e-18, 4.216547e-18, 4.215649e-18, 4.214004e-18, 4.212431e-18, 
    4.212779e-18, 4.211612e-18, 4.214653e-18, 4.213391e-18, 4.213888e-18, 
    4.212588e-18, 4.215408e-18, 4.213093e-18, 4.216011e-18, 4.215749e-18, 
    4.214939e-18, 4.213326e-18, 4.212926e-18, 4.212551e-18, 4.212777e-18, 
    4.213957e-18, 4.214138e-18, 4.214952e-18, 4.215192e-18, 4.215803e-18, 
    4.216324e-18, 4.215856e-18, 4.215369e-18, 4.213945e-18, 4.212678e-18, 
    4.211289e-18, 4.210938e-18, 4.20939e-18, 4.210689e-18, 4.208586e-18, 
    4.210433e-18, 4.207207e-18, 4.212916e-18, 4.21043e-18, 4.214893e-18, 
    4.214404e-18, 4.213551e-18, 4.211538e-18, 4.212594e-18, 4.211344e-18, 
    4.214143e-18, 4.215633e-18, 4.215983e-18, 4.216695e-18, 4.215967e-18, 
    4.216025e-18, 4.215329e-18, 4.215551e-18, 4.213897e-18, 4.214784e-18, 
    4.212259e-18, 4.211347e-18, 4.208741e-18, 4.207165e-18, 4.205518e-18, 
    4.204806e-18, 4.204588e-18, 4.204497e-18 ;

 MEG_acetic_acid =
  6.333174e-19, 6.330936e-19, 6.33136e-19, 6.32958e-19, 6.330552e-19, 
    6.329398e-19, 6.332701e-19, 6.330864e-19, 6.332026e-19, 6.332948e-19, 
    6.326186e-19, 6.329496e-19, 6.32258e-19, 6.324713e-19, 6.319306e-19, 
    6.322936e-19, 6.318567e-19, 6.319368e-19, 6.316857e-19, 6.317573e-19, 
    6.314454e-19, 6.316525e-19, 6.312772e-19, 6.314925e-19, 6.314605e-19, 
    6.3166e-19, 6.328789e-19, 6.326611e-19, 6.328928e-19, 6.328615e-19, 
    6.328746e-19, 6.330547e-19, 6.331483e-19, 6.333317e-19, 6.332976e-19, 
    6.331613e-19, 6.328473e-19, 6.32951e-19, 6.326816e-19, 6.326875e-19, 
    6.32391e-19, 6.325247e-19, 6.32024e-19, 6.321652e-19, 6.317542e-19, 
    6.318581e-19, 6.317598e-19, 6.317891e-19, 6.317595e-19, 6.319115e-19, 
    6.318466e-19, 6.319792e-19, 6.325005e-19, 6.323485e-19, 6.328046e-19, 
    6.33086e-19, 6.332629e-19, 6.333916e-19, 6.333735e-19, 6.333396e-19, 
    6.331606e-19, 6.329889e-19, 6.328594e-19, 6.327736e-19, 6.326884e-19, 
    6.32442e-19, 6.323025e-19, 6.319976e-19, 6.32049e-19, 6.319591e-19, 
    6.318682e-19, 6.317207e-19, 6.317444e-19, 6.316802e-19, 6.319589e-19, 
    6.317749e-19, 6.320791e-19, 6.319963e-19, 6.326796e-19, 6.329224e-19, 
    6.33038e-19, 6.331284e-19, 6.333597e-19, 6.332008e-19, 6.332637e-19, 
    6.33111e-19, 6.330159e-19, 6.330623e-19, 6.327712e-19, 6.328848e-19, 
    6.322943e-19, 6.325482e-19, 6.318788e-19, 6.320381e-19, 6.318402e-19, 
    6.319404e-19, 6.317698e-19, 6.319233e-19, 6.316552e-19, 6.315985e-19, 
    6.316375e-19, 6.314829e-19, 6.319322e-19, 6.317612e-19, 6.330643e-19, 
    6.330568e-19, 6.330204e-19, 6.331811e-19, 6.331902e-19, 6.333333e-19, 
    6.332046e-19, 6.33151e-19, 6.330093e-19, 6.329283e-19, 6.328503e-19, 
    6.326789e-19, 6.324901e-19, 6.322223e-19, 6.320279e-19, 6.318985e-19, 
    6.319769e-19, 6.319078e-19, 6.319856e-19, 6.320215e-19, 6.316207e-19, 
    6.318468e-19, 6.315051e-19, 6.315235e-19, 6.316792e-19, 6.315215e-19, 
    6.330514e-19, 6.330948e-19, 6.332505e-19, 6.331286e-19, 6.333487e-19, 
    6.332273e-19, 6.331585e-19, 6.328857e-19, 6.328223e-19, 6.32768e-19, 
    6.326577e-19, 6.32518e-19, 6.32274e-19, 6.320597e-19, 6.318624e-19, 
    6.318765e-19, 6.318717e-19, 6.318291e-19, 6.319365e-19, 6.318114e-19, 
    6.317917e-19, 6.318452e-19, 6.315261e-19, 6.31617e-19, 6.31524e-19, 
    6.315827e-19, 6.330803e-19, 6.330065e-19, 6.330466e-19, 6.32972e-19, 
    6.330257e-19, 6.327912e-19, 6.327209e-19, 6.323889e-19, 6.325215e-19, 
    6.323065e-19, 6.324985e-19, 6.324653e-19, 6.323055e-19, 6.324872e-19, 
    6.320742e-19, 6.323594e-19, 6.318275e-19, 6.321175e-19, 6.318096e-19, 
    6.318632e-19, 6.31773e-19, 6.316938e-19, 6.315916e-19, 6.314074e-19, 
    6.314495e-19, 6.312933e-19, 6.328952e-19, 6.328009e-19, 6.328066e-19, 
    6.327061e-19, 6.326324e-19, 6.324695e-19, 6.322117e-19, 6.323077e-19, 
    6.321285e-19, 6.320934e-19, 6.323641e-19, 6.322004e-19, 6.327358e-19, 
    6.32652e-19, 6.326999e-19, 6.328893e-19, 6.322893e-19, 6.325985e-19, 
    6.320252e-19, 6.321919e-19, 6.317055e-19, 6.319499e-19, 6.314732e-19, 
    6.312769e-19, 6.3108e-19, 6.308645e-19, 6.327466e-19, 6.328109e-19, 
    6.326933e-19, 6.325358e-19, 6.323821e-19, 6.321823e-19, 6.321603e-19, 
    6.321238e-19, 6.320256e-19, 6.319445e-19, 6.321147e-19, 6.31924e-19, 
    6.326379e-19, 6.322612e-19, 6.328377e-19, 6.326675e-19, 6.325439e-19, 
    6.325954e-19, 6.32318e-19, 6.322536e-19, 6.319933e-19, 6.321263e-19, 
    6.313277e-19, 6.316808e-19, 6.306919e-19, 6.309693e-19, 6.32834e-19, 
    6.327455e-19, 6.324418e-19, 6.325858e-19, 6.321675e-19, 6.320659e-19, 
    6.31981e-19, 6.31877e-19, 6.318638e-19, 6.318018e-19, 6.319036e-19, 
    6.318048e-19, 6.321818e-19, 6.320128e-19, 6.324733e-19, 6.323627e-19, 
    6.324126e-19, 6.324694e-19, 6.322945e-19, 6.321128e-19, 6.321045e-19, 
    6.320471e-19, 6.318928e-19, 6.321657e-19, 6.3129e-19, 6.318376e-19, 
    6.326493e-19, 6.32485e-19, 6.324564e-19, 6.325209e-19, 6.320762e-19, 
    6.322377e-19, 6.318027e-19, 6.319193e-19, 6.317273e-19, 6.31823e-19, 
    6.318373e-19, 6.319594e-19, 6.320366e-19, 6.322312e-19, 6.323884e-19, 
    6.325109e-19, 6.324821e-19, 6.323474e-19, 6.321006e-19, 6.318646e-19, 
    6.319168e-19, 6.317418e-19, 6.321979e-19, 6.320087e-19, 6.320831e-19, 
    6.318882e-19, 6.323111e-19, 6.31964e-19, 6.324016e-19, 6.323623e-19, 
    6.322409e-19, 6.319988e-19, 6.319388e-19, 6.318827e-19, 6.319165e-19, 
    6.320935e-19, 6.321207e-19, 6.322428e-19, 6.322787e-19, 6.323705e-19, 
    6.324486e-19, 6.323783e-19, 6.323054e-19, 6.320917e-19, 6.319017e-19, 
    6.316934e-19, 6.316408e-19, 6.314085e-19, 6.316034e-19, 6.312878e-19, 
    6.315649e-19, 6.310811e-19, 6.319375e-19, 6.315645e-19, 6.322339e-19, 
    6.321606e-19, 6.320327e-19, 6.317306e-19, 6.318891e-19, 6.317017e-19, 
    6.321214e-19, 6.323449e-19, 6.323974e-19, 6.325043e-19, 6.32395e-19, 
    6.324037e-19, 6.322994e-19, 6.323326e-19, 6.320845e-19, 6.322176e-19, 
    6.318388e-19, 6.31702e-19, 6.313111e-19, 6.310748e-19, 6.308276e-19, 
    6.307209e-19, 6.306881e-19, 6.306746e-19 ;

 MEG_acetone =
  1.325753e-16, 1.325506e-16, 1.325552e-16, 1.325356e-16, 1.325463e-16, 
    1.325336e-16, 1.325701e-16, 1.325498e-16, 1.325626e-16, 1.325728e-16, 
    1.324981e-16, 1.325347e-16, 1.324584e-16, 1.324819e-16, 1.324222e-16, 
    1.324623e-16, 1.324141e-16, 1.324229e-16, 1.323952e-16, 1.324031e-16, 
    1.323688e-16, 1.323916e-16, 1.323502e-16, 1.32374e-16, 1.323704e-16, 
    1.323924e-16, 1.325269e-16, 1.325028e-16, 1.325284e-16, 1.325249e-16, 
    1.325264e-16, 1.325463e-16, 1.325566e-16, 1.325768e-16, 1.325731e-16, 
    1.32558e-16, 1.325234e-16, 1.325348e-16, 1.325051e-16, 1.325057e-16, 
    1.32473e-16, 1.324878e-16, 1.324325e-16, 1.324481e-16, 1.324028e-16, 
    1.324142e-16, 1.324034e-16, 1.324066e-16, 1.324034e-16, 1.324201e-16, 
    1.32413e-16, 1.324276e-16, 1.324851e-16, 1.324683e-16, 1.325187e-16, 
    1.325497e-16, 1.325692e-16, 1.325835e-16, 1.325815e-16, 1.325777e-16, 
    1.325579e-16, 1.32539e-16, 1.325247e-16, 1.325152e-16, 1.325058e-16, 
    1.324787e-16, 1.324633e-16, 1.324296e-16, 1.324353e-16, 1.324254e-16, 
    1.324154e-16, 1.323991e-16, 1.324017e-16, 1.323946e-16, 1.324254e-16, 
    1.324051e-16, 1.324386e-16, 1.324295e-16, 1.325049e-16, 1.325317e-16, 
    1.325444e-16, 1.325544e-16, 1.325799e-16, 1.325624e-16, 1.325693e-16, 
    1.325525e-16, 1.32542e-16, 1.325471e-16, 1.32515e-16, 1.325275e-16, 
    1.324624e-16, 1.324904e-16, 1.324165e-16, 1.324341e-16, 1.324123e-16, 
    1.324233e-16, 1.324045e-16, 1.324214e-16, 1.323919e-16, 1.323856e-16, 
    1.323899e-16, 1.323729e-16, 1.324224e-16, 1.324036e-16, 1.325473e-16, 
    1.325465e-16, 1.325425e-16, 1.325602e-16, 1.325612e-16, 1.32577e-16, 
    1.325628e-16, 1.325569e-16, 1.325413e-16, 1.325323e-16, 1.325237e-16, 
    1.325048e-16, 1.32484e-16, 1.324544e-16, 1.32433e-16, 1.324187e-16, 
    1.324273e-16, 1.324197e-16, 1.324283e-16, 1.324323e-16, 1.323881e-16, 
    1.32413e-16, 1.323754e-16, 1.323774e-16, 1.323945e-16, 1.323772e-16, 
    1.325459e-16, 1.325507e-16, 1.325679e-16, 1.325544e-16, 1.325787e-16, 
    1.325653e-16, 1.325577e-16, 1.325276e-16, 1.325206e-16, 1.325146e-16, 
    1.325024e-16, 1.32487e-16, 1.324601e-16, 1.324365e-16, 1.324147e-16, 
    1.324163e-16, 1.324157e-16, 1.32411e-16, 1.324229e-16, 1.324091e-16, 
    1.324069e-16, 1.324128e-16, 1.323777e-16, 1.323877e-16, 1.323774e-16, 
    1.323839e-16, 1.325491e-16, 1.325409e-16, 1.325454e-16, 1.325371e-16, 
    1.325431e-16, 1.325172e-16, 1.325094e-16, 1.324728e-16, 1.324874e-16, 
    1.324637e-16, 1.324849e-16, 1.324812e-16, 1.324636e-16, 1.324836e-16, 
    1.324381e-16, 1.324695e-16, 1.324109e-16, 1.324428e-16, 1.324089e-16, 
    1.324148e-16, 1.324049e-16, 1.323961e-16, 1.323849e-16, 1.323646e-16, 
    1.323692e-16, 1.32352e-16, 1.325287e-16, 1.325183e-16, 1.325189e-16, 
    1.325078e-16, 1.324997e-16, 1.324817e-16, 1.324532e-16, 1.324638e-16, 
    1.324441e-16, 1.324402e-16, 1.324701e-16, 1.32452e-16, 1.325111e-16, 
    1.325018e-16, 1.325071e-16, 1.32528e-16, 1.324618e-16, 1.324959e-16, 
    1.324327e-16, 1.324511e-16, 1.323974e-16, 1.324244e-16, 1.323718e-16, 
    1.323502e-16, 1.323286e-16, 1.323049e-16, 1.325123e-16, 1.325194e-16, 
    1.325064e-16, 1.32489e-16, 1.32472e-16, 1.3245e-16, 1.324476e-16, 
    1.324436e-16, 1.324327e-16, 1.324238e-16, 1.324425e-16, 1.324215e-16, 
    1.325003e-16, 1.324587e-16, 1.325223e-16, 1.325035e-16, 1.324899e-16, 
    1.324956e-16, 1.32465e-16, 1.324579e-16, 1.324291e-16, 1.324438e-16, 
    1.323558e-16, 1.323947e-16, 1.322859e-16, 1.323164e-16, 1.325219e-16, 
    1.325121e-16, 1.324786e-16, 1.324945e-16, 1.324484e-16, 1.324371e-16, 
    1.324278e-16, 1.324163e-16, 1.324149e-16, 1.32408e-16, 1.324193e-16, 
    1.324084e-16, 1.3245e-16, 1.324313e-16, 1.324821e-16, 1.324699e-16, 
    1.324754e-16, 1.324817e-16, 1.324624e-16, 1.324423e-16, 1.324414e-16, 
    1.324351e-16, 1.324181e-16, 1.324482e-16, 1.323517e-16, 1.32412e-16, 
    1.325015e-16, 1.324834e-16, 1.324802e-16, 1.324874e-16, 1.324383e-16, 
    1.324561e-16, 1.324081e-16, 1.32421e-16, 1.323998e-16, 1.324104e-16, 
    1.324119e-16, 1.324254e-16, 1.324339e-16, 1.324554e-16, 1.324727e-16, 
    1.324863e-16, 1.324831e-16, 1.324682e-16, 1.32441e-16, 1.32415e-16, 
    1.324207e-16, 1.324014e-16, 1.324517e-16, 1.324308e-16, 1.324391e-16, 
    1.324176e-16, 1.324642e-16, 1.324259e-16, 1.324742e-16, 1.324699e-16, 
    1.324565e-16, 1.324297e-16, 1.324231e-16, 1.32417e-16, 1.324207e-16, 
    1.324402e-16, 1.324432e-16, 1.324567e-16, 1.324606e-16, 1.324708e-16, 
    1.324794e-16, 1.324716e-16, 1.324636e-16, 1.3244e-16, 1.32419e-16, 
    1.323961e-16, 1.323903e-16, 1.323647e-16, 1.323862e-16, 1.323514e-16, 
    1.323819e-16, 1.323287e-16, 1.32423e-16, 1.323819e-16, 1.324557e-16, 
    1.324476e-16, 1.324335e-16, 1.324002e-16, 1.324177e-16, 1.32397e-16, 
    1.324433e-16, 1.324679e-16, 1.324737e-16, 1.324855e-16, 1.324735e-16, 
    1.324744e-16, 1.324629e-16, 1.324666e-16, 1.324392e-16, 1.324539e-16, 
    1.324121e-16, 1.32397e-16, 1.32354e-16, 1.32328e-16, 1.323008e-16, 
    1.322891e-16, 1.322854e-16, 1.32284e-16 ;

 MEG_carene_3 =
  5.257901e-17, 5.256874e-17, 5.257069e-17, 5.256252e-17, 5.256698e-17, 
    5.256169e-17, 5.257684e-17, 5.256841e-17, 5.257374e-17, 5.257797e-17, 
    5.254696e-17, 5.256213e-17, 5.253043e-17, 5.254021e-17, 5.251541e-17, 
    5.253206e-17, 5.251203e-17, 5.25157e-17, 5.25042e-17, 5.250748e-17, 
    5.24932e-17, 5.250268e-17, 5.24855e-17, 5.249536e-17, 5.249389e-17, 
    5.250303e-17, 5.255889e-17, 5.25489e-17, 5.255953e-17, 5.255809e-17, 
    5.25587e-17, 5.256695e-17, 5.257125e-17, 5.257966e-17, 5.25781e-17, 
    5.257184e-17, 5.255744e-17, 5.25622e-17, 5.254984e-17, 5.255012e-17, 
    5.253652e-17, 5.254265e-17, 5.25197e-17, 5.252617e-17, 5.250734e-17, 
    5.25121e-17, 5.250759e-17, 5.250893e-17, 5.250758e-17, 5.251454e-17, 
    5.251157e-17, 5.251764e-17, 5.254154e-17, 5.253457e-17, 5.255549e-17, 
    5.256839e-17, 5.25765e-17, 5.258241e-17, 5.258158e-17, 5.258002e-17, 
    5.257181e-17, 5.256394e-17, 5.2558e-17, 5.255406e-17, 5.255016e-17, 
    5.253886e-17, 5.253246e-17, 5.251848e-17, 5.252084e-17, 5.251672e-17, 
    5.251256e-17, 5.25058e-17, 5.250689e-17, 5.250395e-17, 5.251671e-17, 
    5.250828e-17, 5.252222e-17, 5.251843e-17, 5.254975e-17, 5.256088e-17, 
    5.256619e-17, 5.257034e-17, 5.258095e-17, 5.257365e-17, 5.257654e-17, 
    5.256953e-17, 5.256518e-17, 5.25673e-17, 5.255395e-17, 5.255917e-17, 
    5.253209e-17, 5.254373e-17, 5.251305e-17, 5.252034e-17, 5.251127e-17, 
    5.251587e-17, 5.250805e-17, 5.251508e-17, 5.25028e-17, 5.250021e-17, 
    5.250199e-17, 5.249492e-17, 5.251549e-17, 5.250766e-17, 5.256739e-17, 
    5.256705e-17, 5.256538e-17, 5.257275e-17, 5.257317e-17, 5.257974e-17, 
    5.257383e-17, 5.257137e-17, 5.256487e-17, 5.256116e-17, 5.255758e-17, 
    5.254972e-17, 5.254106e-17, 5.252879e-17, 5.251988e-17, 5.251395e-17, 
    5.251754e-17, 5.251437e-17, 5.251794e-17, 5.251958e-17, 5.250122e-17, 
    5.251158e-17, 5.249594e-17, 5.249678e-17, 5.25039e-17, 5.249668e-17, 
    5.25668e-17, 5.256879e-17, 5.257594e-17, 5.257035e-17, 5.258044e-17, 
    5.257487e-17, 5.257172e-17, 5.25592e-17, 5.255629e-17, 5.255381e-17, 
    5.254875e-17, 5.254234e-17, 5.253116e-17, 5.252133e-17, 5.251229e-17, 
    5.251294e-17, 5.251272e-17, 5.251077e-17, 5.251569e-17, 5.250995e-17, 
    5.250905e-17, 5.25115e-17, 5.249689e-17, 5.250105e-17, 5.24968e-17, 
    5.249949e-17, 5.256813e-17, 5.256474e-17, 5.256658e-17, 5.256316e-17, 
    5.256562e-17, 5.255487e-17, 5.255164e-17, 5.253642e-17, 5.254251e-17, 
    5.253265e-17, 5.254145e-17, 5.253993e-17, 5.25326e-17, 5.254093e-17, 
    5.2522e-17, 5.253507e-17, 5.251069e-17, 5.252398e-17, 5.250988e-17, 
    5.251233e-17, 5.25082e-17, 5.250457e-17, 5.249989e-17, 5.249146e-17, 
    5.249338e-17, 5.248624e-17, 5.255964e-17, 5.255531e-17, 5.255558e-17, 
    5.255097e-17, 5.254759e-17, 5.254012e-17, 5.25283e-17, 5.25327e-17, 
    5.252449e-17, 5.252288e-17, 5.253529e-17, 5.252779e-17, 5.255233e-17, 
    5.254849e-17, 5.255069e-17, 5.255937e-17, 5.253186e-17, 5.254604e-17, 
    5.251976e-17, 5.25274e-17, 5.250511e-17, 5.25163e-17, 5.249447e-17, 
    5.248549e-17, 5.247648e-17, 5.246663e-17, 5.255282e-17, 5.255577e-17, 
    5.255038e-17, 5.254316e-17, 5.253611e-17, 5.252695e-17, 5.252595e-17, 
    5.252427e-17, 5.251977e-17, 5.251605e-17, 5.252386e-17, 5.251511e-17, 
    5.254784e-17, 5.253057e-17, 5.2557e-17, 5.25492e-17, 5.254353e-17, 
    5.254589e-17, 5.253318e-17, 5.253023e-17, 5.251829e-17, 5.252439e-17, 
    5.248781e-17, 5.250398e-17, 5.245874e-17, 5.247142e-17, 5.255683e-17, 
    5.255278e-17, 5.253885e-17, 5.254545e-17, 5.252628e-17, 5.252161e-17, 
    5.251773e-17, 5.251296e-17, 5.251235e-17, 5.250952e-17, 5.251418e-17, 
    5.250966e-17, 5.252694e-17, 5.251918e-17, 5.25403e-17, 5.253523e-17, 
    5.253752e-17, 5.254012e-17, 5.25321e-17, 5.252377e-17, 5.252339e-17, 
    5.252075e-17, 5.251368e-17, 5.252619e-17, 5.248609e-17, 5.251115e-17, 
    5.254837e-17, 5.254083e-17, 5.253952e-17, 5.254248e-17, 5.252209e-17, 
    5.25295e-17, 5.250956e-17, 5.251489e-17, 5.25061e-17, 5.251049e-17, 
    5.251114e-17, 5.251673e-17, 5.252027e-17, 5.252919e-17, 5.25364e-17, 
    5.254202e-17, 5.25407e-17, 5.253453e-17, 5.252321e-17, 5.251239e-17, 
    5.251478e-17, 5.250677e-17, 5.252767e-17, 5.251899e-17, 5.252241e-17, 
    5.251348e-17, 5.253286e-17, 5.251694e-17, 5.253701e-17, 5.253521e-17, 
    5.252964e-17, 5.251854e-17, 5.251579e-17, 5.251322e-17, 5.251477e-17, 
    5.252288e-17, 5.252413e-17, 5.252973e-17, 5.253138e-17, 5.253558e-17, 
    5.253917e-17, 5.253594e-17, 5.25326e-17, 5.25228e-17, 5.251409e-17, 
    5.250455e-17, 5.250214e-17, 5.249151e-17, 5.250043e-17, 5.248598e-17, 
    5.249866e-17, 5.247653e-17, 5.251573e-17, 5.249865e-17, 5.252932e-17, 
    5.252596e-17, 5.252009e-17, 5.250626e-17, 5.251351e-17, 5.250493e-17, 
    5.252417e-17, 5.253441e-17, 5.253682e-17, 5.254172e-17, 5.253671e-17, 
    5.253711e-17, 5.253232e-17, 5.253385e-17, 5.252247e-17, 5.252857e-17, 
    5.251121e-17, 5.250495e-17, 5.248706e-17, 5.247624e-17, 5.246495e-17, 
    5.246007e-17, 5.245857e-17, 5.245795e-17 ;

 MEG_ethanol =
  4.222116e-18, 4.220624e-18, 4.220907e-18, 4.21972e-18, 4.220368e-18, 
    4.219599e-18, 4.221801e-18, 4.220576e-18, 4.221351e-18, 4.221965e-18, 
    4.217458e-18, 4.219664e-18, 4.215054e-18, 4.216476e-18, 4.212871e-18, 
    4.215291e-18, 4.212378e-18, 4.212912e-18, 4.211238e-18, 4.211715e-18, 
    4.209636e-18, 4.211017e-18, 4.208515e-18, 4.20995e-18, 4.209736e-18, 
    4.211067e-18, 4.219193e-18, 4.217741e-18, 4.219285e-18, 4.219076e-18, 
    4.219164e-18, 4.220364e-18, 4.220989e-18, 4.222212e-18, 4.221984e-18, 
    4.221076e-18, 4.218982e-18, 4.219674e-18, 4.217877e-18, 4.217917e-18, 
    4.21594e-18, 4.216832e-18, 4.213494e-18, 4.214435e-18, 4.211695e-18, 
    4.212387e-18, 4.211732e-18, 4.211927e-18, 4.21173e-18, 4.212744e-18, 
    4.212311e-18, 4.213194e-18, 4.21667e-18, 4.215657e-18, 4.218698e-18, 
    4.220574e-18, 4.221752e-18, 4.222611e-18, 4.22249e-18, 4.222264e-18, 
    4.221071e-18, 4.219926e-18, 4.219063e-18, 4.218491e-18, 4.217923e-18, 
    4.21628e-18, 4.21535e-18, 4.213317e-18, 4.21366e-18, 4.213061e-18, 
    4.212455e-18, 4.211471e-18, 4.211629e-18, 4.211202e-18, 4.213059e-18, 
    4.211833e-18, 4.213861e-18, 4.213309e-18, 4.217864e-18, 4.219482e-18, 
    4.220254e-18, 4.220857e-18, 4.222398e-18, 4.221339e-18, 4.221759e-18, 
    4.22074e-18, 4.220107e-18, 4.220416e-18, 4.218475e-18, 4.219232e-18, 
    4.215295e-18, 4.216988e-18, 4.212526e-18, 4.213588e-18, 4.212268e-18, 
    4.212936e-18, 4.211799e-18, 4.212822e-18, 4.211035e-18, 4.210657e-18, 
    4.210917e-18, 4.209887e-18, 4.212881e-18, 4.211741e-18, 4.220429e-18, 
    4.220379e-18, 4.220136e-18, 4.221207e-18, 4.221268e-18, 4.222222e-18, 
    4.221364e-18, 4.221007e-18, 4.220062e-18, 4.219522e-18, 4.219002e-18, 
    4.217859e-18, 4.2166e-18, 4.214816e-18, 4.21352e-18, 4.212657e-18, 
    4.21318e-18, 4.212719e-18, 4.213237e-18, 4.213476e-18, 4.210805e-18, 
    4.212312e-18, 4.210035e-18, 4.210157e-18, 4.211195e-18, 4.210143e-18, 
    4.220342e-18, 4.220632e-18, 4.22167e-18, 4.220858e-18, 4.222325e-18, 
    4.221515e-18, 4.221057e-18, 4.219238e-18, 4.218815e-18, 4.218454e-18, 
    4.217718e-18, 4.216786e-18, 4.21516e-18, 4.213732e-18, 4.212416e-18, 
    4.212511e-18, 4.212478e-18, 4.212194e-18, 4.21291e-18, 4.212076e-18, 
    4.211945e-18, 4.212301e-18, 4.210174e-18, 4.21078e-18, 4.21016e-18, 
    4.210552e-18, 4.220536e-18, 4.220043e-18, 4.220311e-18, 4.219814e-18, 
    4.220171e-18, 4.218608e-18, 4.21814e-18, 4.215926e-18, 4.21681e-18, 
    4.215377e-18, 4.216657e-18, 4.216435e-18, 4.21537e-18, 4.216581e-18, 
    4.213828e-18, 4.21573e-18, 4.212183e-18, 4.214116e-18, 4.212064e-18, 
    4.212422e-18, 4.21182e-18, 4.211292e-18, 4.210611e-18, 4.209383e-18, 
    4.209663e-18, 4.208622e-18, 4.219301e-18, 4.218673e-18, 4.21871e-18, 
    4.21804e-18, 4.21755e-18, 4.216463e-18, 4.214745e-18, 4.215385e-18, 
    4.21419e-18, 4.213956e-18, 4.215761e-18, 4.21467e-18, 4.218239e-18, 
    4.21768e-18, 4.217999e-18, 4.219262e-18, 4.215262e-18, 4.217324e-18, 
    4.213502e-18, 4.214613e-18, 4.21137e-18, 4.213e-18, 4.209822e-18, 
    4.208513e-18, 4.2072e-18, 4.205763e-18, 4.218311e-18, 4.218739e-18, 
    4.217956e-18, 4.216906e-18, 4.215881e-18, 4.214549e-18, 4.214403e-18, 
    4.214158e-18, 4.213504e-18, 4.212964e-18, 4.214099e-18, 4.212826e-18, 
    4.217586e-18, 4.215075e-18, 4.218918e-18, 4.217784e-18, 4.216959e-18, 
    4.217303e-18, 4.215453e-18, 4.215025e-18, 4.213289e-18, 4.214175e-18, 
    4.208851e-18, 4.211206e-18, 4.204613e-18, 4.206462e-18, 4.218894e-18, 
    4.218303e-18, 4.216279e-18, 4.217239e-18, 4.21445e-18, 4.213773e-18, 
    4.213207e-18, 4.212513e-18, 4.212425e-18, 4.212012e-18, 4.212691e-18, 
    4.212032e-18, 4.214546e-18, 4.213419e-18, 4.216489e-18, 4.215751e-18, 
    4.216084e-18, 4.216463e-18, 4.215297e-18, 4.214085e-18, 4.214031e-18, 
    4.213647e-18, 4.212619e-18, 4.214438e-18, 4.2086e-18, 4.212251e-18, 
    4.217662e-18, 4.216567e-18, 4.216376e-18, 4.216806e-18, 4.213841e-18, 
    4.214918e-18, 4.212019e-18, 4.212795e-18, 4.211515e-18, 4.212153e-18, 
    4.212249e-18, 4.213062e-18, 4.213577e-18, 4.214874e-18, 4.215923e-18, 
    4.21674e-18, 4.216547e-18, 4.215649e-18, 4.214004e-18, 4.212431e-18, 
    4.212779e-18, 4.211612e-18, 4.214653e-18, 4.213391e-18, 4.213888e-18, 
    4.212588e-18, 4.215408e-18, 4.213093e-18, 4.216011e-18, 4.215749e-18, 
    4.214939e-18, 4.213326e-18, 4.212926e-18, 4.212551e-18, 4.212777e-18, 
    4.213957e-18, 4.214138e-18, 4.214952e-18, 4.215192e-18, 4.215803e-18, 
    4.216324e-18, 4.215856e-18, 4.215369e-18, 4.213945e-18, 4.212678e-18, 
    4.211289e-18, 4.210938e-18, 4.20939e-18, 4.210689e-18, 4.208586e-18, 
    4.210433e-18, 4.207207e-18, 4.212916e-18, 4.21043e-18, 4.214893e-18, 
    4.214404e-18, 4.213551e-18, 4.211538e-18, 4.212594e-18, 4.211344e-18, 
    4.214143e-18, 4.215633e-18, 4.215983e-18, 4.216695e-18, 4.215967e-18, 
    4.216025e-18, 4.215329e-18, 4.215551e-18, 4.213897e-18, 4.214784e-18, 
    4.212259e-18, 4.211347e-18, 4.208741e-18, 4.207165e-18, 4.205518e-18, 
    4.204806e-18, 4.204588e-18, 4.204497e-18 ;

 MEG_formaldehyde =
  8.444232e-19, 8.441248e-19, 8.441814e-19, 8.43944e-19, 8.440736e-19, 
    8.439198e-19, 8.443602e-19, 8.441152e-19, 8.442701e-19, 8.443929e-19, 
    8.434915e-19, 8.439328e-19, 8.430107e-19, 8.432951e-19, 8.425741e-19, 
    8.430581e-19, 8.424756e-19, 8.425824e-19, 8.422476e-19, 8.42343e-19, 
    8.419272e-19, 8.422033e-19, 8.417029e-19, 8.4199e-19, 8.419473e-19, 
    8.422134e-19, 8.438385e-19, 8.435481e-19, 8.43857e-19, 8.438153e-19, 
    8.438328e-19, 8.440729e-19, 8.441977e-19, 8.444423e-19, 8.443968e-19, 
    8.442151e-19, 8.437964e-19, 8.439347e-19, 8.435754e-19, 8.435833e-19, 
    8.43188e-19, 8.433663e-19, 8.426987e-19, 8.42887e-19, 8.42339e-19, 
    8.424775e-19, 8.423464e-19, 8.423854e-19, 8.423459e-19, 8.425487e-19, 
    8.424622e-19, 8.426389e-19, 8.43334e-19, 8.431313e-19, 8.437395e-19, 
    8.441147e-19, 8.443505e-19, 8.445222e-19, 8.444979e-19, 8.444528e-19, 
    8.442141e-19, 8.439852e-19, 8.438126e-19, 8.436981e-19, 8.435845e-19, 
    8.43256e-19, 8.4307e-19, 8.426635e-19, 8.42732e-19, 8.426122e-19, 
    8.42491e-19, 8.422942e-19, 8.423258e-19, 8.422403e-19, 8.426118e-19, 
    8.423666e-19, 8.427721e-19, 8.426618e-19, 8.435728e-19, 8.438964e-19, 
    8.440507e-19, 8.441713e-19, 8.444796e-19, 8.442677e-19, 8.443516e-19, 
    8.441479e-19, 8.440213e-19, 8.440831e-19, 8.43695e-19, 8.438465e-19, 
    8.430591e-19, 8.433976e-19, 8.425051e-19, 8.427175e-19, 8.424536e-19, 
    8.425872e-19, 8.423597e-19, 8.425644e-19, 8.42207e-19, 8.421314e-19, 
    8.421834e-19, 8.419772e-19, 8.425763e-19, 8.423483e-19, 8.440857e-19, 
    8.440758e-19, 8.440272e-19, 8.442415e-19, 8.442536e-19, 8.444444e-19, 
    8.442728e-19, 8.442014e-19, 8.440124e-19, 8.439044e-19, 8.438004e-19, 
    8.435719e-19, 8.4332e-19, 8.429631e-19, 8.427039e-19, 8.425314e-19, 
    8.426359e-19, 8.425437e-19, 8.426475e-19, 8.426953e-19, 8.42161e-19, 
    8.424624e-19, 8.420069e-19, 8.420314e-19, 8.42239e-19, 8.420286e-19, 
    8.440685e-19, 8.441264e-19, 8.44334e-19, 8.441715e-19, 8.44465e-19, 
    8.443031e-19, 8.442114e-19, 8.438475e-19, 8.43763e-19, 8.436907e-19, 
    8.435436e-19, 8.433573e-19, 8.430319e-19, 8.427463e-19, 8.424831e-19, 
    8.425021e-19, 8.424956e-19, 8.424388e-19, 8.42582e-19, 8.424152e-19, 
    8.423889e-19, 8.424602e-19, 8.420348e-19, 8.42156e-19, 8.42032e-19, 
    8.421103e-19, 8.441071e-19, 8.440087e-19, 8.440621e-19, 8.439627e-19, 
    8.440342e-19, 8.437215e-19, 8.436279e-19, 8.431852e-19, 8.43362e-19, 
    8.430754e-19, 8.433314e-19, 8.432871e-19, 8.43074e-19, 8.433163e-19, 
    8.427656e-19, 8.431459e-19, 8.424366e-19, 8.428233e-19, 8.424128e-19, 
    8.424843e-19, 8.42364e-19, 8.422585e-19, 8.421222e-19, 8.418766e-19, 
    8.419326e-19, 8.417244e-19, 8.438603e-19, 8.437346e-19, 8.437421e-19, 
    8.436081e-19, 8.435098e-19, 8.432926e-19, 8.429489e-19, 8.430769e-19, 
    8.42838e-19, 8.427912e-19, 8.431522e-19, 8.42934e-19, 8.436477e-19, 
    8.43536e-19, 8.435998e-19, 8.438524e-19, 8.430523e-19, 8.434647e-19, 
    8.427003e-19, 8.429225e-19, 8.42274e-19, 8.425998e-19, 8.419643e-19, 
    8.417025e-19, 8.4144e-19, 8.411527e-19, 8.436621e-19, 8.437479e-19, 
    8.43591e-19, 8.43381e-19, 8.431761e-19, 8.429097e-19, 8.428804e-19, 
    8.428317e-19, 8.427008e-19, 8.425926e-19, 8.428197e-19, 8.425652e-19, 
    8.435172e-19, 8.43015e-19, 8.437836e-19, 8.435567e-19, 8.433918e-19, 
    8.434605e-19, 8.430907e-19, 8.430048e-19, 8.426577e-19, 8.428351e-19, 
    8.417702e-19, 8.422411e-19, 8.409226e-19, 8.412925e-19, 8.437787e-19, 
    8.436607e-19, 8.432557e-19, 8.434477e-19, 8.4289e-19, 8.427545e-19, 
    8.426413e-19, 8.425026e-19, 8.42485e-19, 8.424024e-19, 8.425382e-19, 
    8.424064e-19, 8.429091e-19, 8.426837e-19, 8.432977e-19, 8.431502e-19, 
    8.432168e-19, 8.432925e-19, 8.430593e-19, 8.42817e-19, 8.428061e-19, 
    8.427294e-19, 8.425237e-19, 8.428876e-19, 8.417201e-19, 8.424501e-19, 
    8.435324e-19, 8.433134e-19, 8.432751e-19, 8.433611e-19, 8.427683e-19, 
    8.429836e-19, 8.424036e-19, 8.42559e-19, 8.42303e-19, 8.424307e-19, 
    8.424497e-19, 8.426125e-19, 8.427155e-19, 8.429749e-19, 8.431845e-19, 
    8.433479e-19, 8.433095e-19, 8.431298e-19, 8.428008e-19, 8.42486e-19, 
    8.425557e-19, 8.423224e-19, 8.429305e-19, 8.426783e-19, 8.427776e-19, 
    8.425176e-19, 8.430816e-19, 8.426186e-19, 8.432021e-19, 8.431497e-19, 
    8.429878e-19, 8.426651e-19, 8.425851e-19, 8.425103e-19, 8.425553e-19, 
    8.427913e-19, 8.428276e-19, 8.429904e-19, 8.430382e-19, 8.431607e-19, 
    8.432648e-19, 8.431711e-19, 8.430739e-19, 8.427889e-19, 8.425356e-19, 
    8.422579e-19, 8.421876e-19, 8.41878e-19, 8.421378e-19, 8.417171e-19, 
    8.420865e-19, 8.414415e-19, 8.425832e-19, 8.42086e-19, 8.429786e-19, 
    8.428809e-19, 8.427102e-19, 8.423075e-19, 8.425188e-19, 8.422689e-19, 
    8.428285e-19, 8.431265e-19, 8.431965e-19, 8.43339e-19, 8.431933e-19, 
    8.432049e-19, 8.430658e-19, 8.431101e-19, 8.427793e-19, 8.429568e-19, 
    8.424517e-19, 8.422694e-19, 8.417482e-19, 8.41433e-19, 8.411035e-19, 
    8.409612e-19, 8.409174e-19, 8.408995e-19 ;

 MEG_isoprene =
  6.66767e-19, 6.6649e-19, 6.665425e-19, 6.663222e-19, 6.664424e-19, 
    6.662997e-19, 6.667085e-19, 6.664811e-19, 6.666249e-19, 6.667389e-19, 
    6.659022e-19, 6.663117e-19, 6.654558e-19, 6.657198e-19, 6.650505e-19, 
    6.654998e-19, 6.649591e-19, 6.650582e-19, 6.647473e-19, 6.64836e-19, 
    6.644498e-19, 6.647063e-19, 6.642416e-19, 6.645083e-19, 6.644686e-19, 
    6.647156e-19, 6.662242e-19, 6.659547e-19, 6.662414e-19, 6.662027e-19, 
    6.662189e-19, 6.664418e-19, 6.665577e-19, 6.667846e-19, 6.667424e-19, 
    6.665738e-19, 6.661852e-19, 6.663135e-19, 6.6598e-19, 6.659874e-19, 
    6.656204e-19, 6.657858e-19, 6.651662e-19, 6.653409e-19, 6.648322e-19, 
    6.649608e-19, 6.648391e-19, 6.648753e-19, 6.648387e-19, 6.650269e-19, 
    6.649466e-19, 6.651106e-19, 6.657559e-19, 6.655677e-19, 6.661324e-19, 
    6.664806e-19, 6.666995e-19, 6.668588e-19, 6.668364e-19, 6.667944e-19, 
    6.665729e-19, 6.663604e-19, 6.662002e-19, 6.66094e-19, 6.659885e-19, 
    6.656835e-19, 6.655109e-19, 6.651334e-19, 6.65197e-19, 6.650859e-19, 
    6.649733e-19, 6.647907e-19, 6.6482e-19, 6.647406e-19, 6.650855e-19, 
    6.648578e-19, 6.652344e-19, 6.651319e-19, 6.659776e-19, 6.66278e-19, 
    6.664212e-19, 6.665331e-19, 6.668193e-19, 6.666226e-19, 6.667005e-19, 
    6.665114e-19, 6.663939e-19, 6.664513e-19, 6.66091e-19, 6.662316e-19, 
    6.655007e-19, 6.65815e-19, 6.649865e-19, 6.651836e-19, 6.649386e-19, 
    6.650627e-19, 6.648515e-19, 6.650415e-19, 6.647097e-19, 6.646395e-19, 
    6.646878e-19, 6.644964e-19, 6.650525e-19, 6.648408e-19, 6.664537e-19, 
    6.664445e-19, 6.663993e-19, 6.665983e-19, 6.666095e-19, 6.667867e-19, 
    6.666273e-19, 6.66561e-19, 6.663857e-19, 6.662854e-19, 6.661889e-19, 
    6.659767e-19, 6.65743e-19, 6.654116e-19, 6.65171e-19, 6.650109e-19, 
    6.651079e-19, 6.650223e-19, 6.651187e-19, 6.65163e-19, 6.64667e-19, 
    6.649468e-19, 6.645239e-19, 6.645466e-19, 6.647394e-19, 6.645441e-19, 
    6.664377e-19, 6.664915e-19, 6.666842e-19, 6.665333e-19, 6.668057e-19, 
    6.666555e-19, 6.665704e-19, 6.662326e-19, 6.661542e-19, 6.660871e-19, 
    6.659505e-19, 6.657775e-19, 6.654755e-19, 6.652104e-19, 6.649661e-19, 
    6.649836e-19, 6.649776e-19, 6.649249e-19, 6.650579e-19, 6.649029e-19, 
    6.648786e-19, 6.649448e-19, 6.645498e-19, 6.646623e-19, 6.645471e-19, 
    6.646199e-19, 6.664735e-19, 6.663822e-19, 6.664318e-19, 6.663395e-19, 
    6.664059e-19, 6.661157e-19, 6.660287e-19, 6.656178e-19, 6.657819e-19, 
    6.655159e-19, 6.657535e-19, 6.657123e-19, 6.655146e-19, 6.657395e-19, 
    6.652283e-19, 6.655813e-19, 6.649229e-19, 6.652818e-19, 6.649008e-19, 
    6.649671e-19, 6.648555e-19, 6.647575e-19, 6.646309e-19, 6.644029e-19, 
    6.644549e-19, 6.642615e-19, 6.662445e-19, 6.661278e-19, 6.661348e-19, 
    6.660103e-19, 6.659191e-19, 6.657175e-19, 6.653984e-19, 6.655173e-19, 
    6.652955e-19, 6.652521e-19, 6.655872e-19, 6.653846e-19, 6.660471e-19, 
    6.659434e-19, 6.660027e-19, 6.662372e-19, 6.654945e-19, 6.658772e-19, 
    6.651677e-19, 6.65374e-19, 6.647719e-19, 6.650744e-19, 6.644844e-19, 
    6.642413e-19, 6.639974e-19, 6.637307e-19, 6.660605e-19, 6.661401e-19, 
    6.659945e-19, 6.657996e-19, 6.656093e-19, 6.653621e-19, 6.653349e-19, 
    6.652896e-19, 6.651681e-19, 6.650677e-19, 6.652785e-19, 6.650423e-19, 
    6.659259e-19, 6.654598e-19, 6.661733e-19, 6.659626e-19, 6.658096e-19, 
    6.658733e-19, 6.6553e-19, 6.654504e-19, 6.651282e-19, 6.652928e-19, 
    6.643041e-19, 6.647414e-19, 6.635169e-19, 6.638604e-19, 6.661687e-19, 
    6.660592e-19, 6.656833e-19, 6.658615e-19, 6.653438e-19, 6.65218e-19, 
    6.651129e-19, 6.649841e-19, 6.649678e-19, 6.648911e-19, 6.650172e-19, 
    6.648949e-19, 6.653615e-19, 6.651523e-19, 6.657222e-19, 6.655853e-19, 
    6.656471e-19, 6.657174e-19, 6.655009e-19, 6.65276e-19, 6.652658e-19, 
    6.651947e-19, 6.650038e-19, 6.653415e-19, 6.642576e-19, 6.649354e-19, 
    6.659401e-19, 6.657368e-19, 6.657013e-19, 6.657811e-19, 6.652307e-19, 
    6.654307e-19, 6.648923e-19, 6.650365e-19, 6.647989e-19, 6.649173e-19, 
    6.649351e-19, 6.650861e-19, 6.651818e-19, 6.654225e-19, 6.656171e-19, 
    6.657688e-19, 6.657332e-19, 6.655664e-19, 6.65261e-19, 6.649687e-19, 
    6.650334e-19, 6.648168e-19, 6.653814e-19, 6.651472e-19, 6.652394e-19, 
    6.649981e-19, 6.655216e-19, 6.650919e-19, 6.656335e-19, 6.655848e-19, 
    6.654346e-19, 6.651349e-19, 6.650608e-19, 6.649912e-19, 6.65033e-19, 
    6.652522e-19, 6.652859e-19, 6.65437e-19, 6.654814e-19, 6.65595e-19, 
    6.656917e-19, 6.656047e-19, 6.655145e-19, 6.652499e-19, 6.650147e-19, 
    6.647569e-19, 6.646917e-19, 6.644042e-19, 6.646455e-19, 6.642548e-19, 
    6.645978e-19, 6.639988e-19, 6.65059e-19, 6.645974e-19, 6.65426e-19, 
    6.653353e-19, 6.651769e-19, 6.64803e-19, 6.649991e-19, 6.647672e-19, 
    6.652867e-19, 6.655633e-19, 6.656283e-19, 6.657606e-19, 6.656253e-19, 
    6.656361e-19, 6.65507e-19, 6.655481e-19, 6.65241e-19, 6.654057e-19, 
    6.649369e-19, 6.647676e-19, 6.642837e-19, 6.63991e-19, 6.63685e-19, 
    6.635528e-19, 6.635121e-19, 6.634954e-19 ;

 MEG_methanol =
  9.49351e-17, 9.491948e-17, 9.492244e-17, 9.491002e-17, 9.49168e-17, 
    9.490875e-17, 9.49318e-17, 9.491898e-17, 9.492709e-17, 9.493352e-17, 
    9.488634e-17, 9.490943e-17, 9.486119e-17, 9.487608e-17, 9.483835e-17, 
    9.486367e-17, 9.48332e-17, 9.483879e-17, 9.482129e-17, 9.482628e-17, 
    9.480455e-17, 9.481898e-17, 9.479285e-17, 9.480784e-17, 9.48056e-17, 
    9.48195e-17, 9.49045e-17, 9.48893e-17, 9.490547e-17, 9.490328e-17, 
    9.49042e-17, 9.491676e-17, 9.49233e-17, 9.49361e-17, 9.493372e-17, 
    9.49242e-17, 9.490229e-17, 9.490953e-17, 9.489074e-17, 9.489115e-17, 
    9.487047e-17, 9.48798e-17, 9.484487e-17, 9.485473e-17, 9.482607e-17, 
    9.48333e-17, 9.482645e-17, 9.482849e-17, 9.482643e-17, 9.483702e-17, 
    9.48325e-17, 9.484174e-17, 9.487811e-17, 9.48675e-17, 9.489932e-17, 
    9.491895e-17, 9.493129e-17, 9.494028e-17, 9.493901e-17, 9.493665e-17, 
    9.492415e-17, 9.491218e-17, 9.490315e-17, 9.489716e-17, 9.489122e-17, 
    9.487402e-17, 9.48643e-17, 9.484302e-17, 9.484661e-17, 9.484034e-17, 
    9.483401e-17, 9.482372e-17, 9.482538e-17, 9.482091e-17, 9.484033e-17, 
    9.48275e-17, 9.484871e-17, 9.484293e-17, 9.489059e-17, 9.490753e-17, 
    9.491559e-17, 9.492191e-17, 9.493805e-17, 9.492696e-17, 9.493136e-17, 
    9.492069e-17, 9.491407e-17, 9.49173e-17, 9.489699e-17, 9.490491e-17, 
    9.486373e-17, 9.488144e-17, 9.483475e-17, 9.484585e-17, 9.483206e-17, 
    9.483904e-17, 9.482715e-17, 9.483785e-17, 9.481916e-17, 9.481522e-17, 
    9.481793e-17, 9.480717e-17, 9.483847e-17, 9.482655e-17, 9.491743e-17, 
    9.491692e-17, 9.491437e-17, 9.492559e-17, 9.492622e-17, 9.493621e-17, 
    9.492723e-17, 9.492348e-17, 9.49136e-17, 9.490794e-17, 9.49025e-17, 
    9.489055e-17, 9.487738e-17, 9.48587e-17, 9.484514e-17, 9.483612e-17, 
    9.484158e-17, 9.483677e-17, 9.484219e-17, 9.484469e-17, 9.481676e-17, 
    9.483251e-17, 9.480872e-17, 9.481e-17, 9.482084e-17, 9.480985e-17, 
    9.491653e-17, 9.491956e-17, 9.493043e-17, 9.492193e-17, 9.493729e-17, 
    9.492881e-17, 9.492401e-17, 9.490497e-17, 9.490055e-17, 9.489677e-17, 
    9.488908e-17, 9.487933e-17, 9.48623e-17, 9.484735e-17, 9.48336e-17, 
    9.483459e-17, 9.483425e-17, 9.483128e-17, 9.483877e-17, 9.483004e-17, 
    9.482867e-17, 9.48324e-17, 9.481018e-17, 9.48165e-17, 9.481003e-17, 
    9.481412e-17, 9.491855e-17, 9.49134e-17, 9.49162e-17, 9.491099e-17, 
    9.491474e-17, 9.489838e-17, 9.489348e-17, 9.487032e-17, 9.487958e-17, 
    9.486458e-17, 9.487797e-17, 9.487566e-17, 9.48645e-17, 9.487719e-17, 
    9.484837e-17, 9.486827e-17, 9.483117e-17, 9.485138e-17, 9.482992e-17, 
    9.483366e-17, 9.482738e-17, 9.482186e-17, 9.481474e-17, 9.480191e-17, 
    9.480484e-17, 9.479397e-17, 9.490564e-17, 9.489906e-17, 9.489945e-17, 
    9.489245e-17, 9.488731e-17, 9.487595e-17, 9.485796e-17, 9.486466e-17, 
    9.485217e-17, 9.484971e-17, 9.48686e-17, 9.485718e-17, 9.489452e-17, 
    9.488867e-17, 9.489202e-17, 9.490522e-17, 9.486338e-17, 9.488494e-17, 
    9.484495e-17, 9.485659e-17, 9.482267e-17, 9.48397e-17, 9.480649e-17, 
    9.479282e-17, 9.477913e-17, 9.476414e-17, 9.489527e-17, 9.489976e-17, 
    9.489156e-17, 9.488057e-17, 9.486985e-17, 9.485591e-17, 9.485438e-17, 
    9.485183e-17, 9.484498e-17, 9.483933e-17, 9.48512e-17, 9.483789e-17, 
    9.488768e-17, 9.486142e-17, 9.490162e-17, 9.488975e-17, 9.488114e-17, 
    9.488473e-17, 9.486538e-17, 9.486089e-17, 9.484272e-17, 9.485201e-17, 
    9.479635e-17, 9.482094e-17, 9.475215e-17, 9.477143e-17, 9.490137e-17, 
    9.48952e-17, 9.487402e-17, 9.488406e-17, 9.485489e-17, 9.484778e-17, 
    9.484187e-17, 9.483462e-17, 9.48337e-17, 9.482938e-17, 9.483648e-17, 
    9.482959e-17, 9.485588e-17, 9.484409e-17, 9.487621e-17, 9.48685e-17, 
    9.487198e-17, 9.487595e-17, 9.486374e-17, 9.485107e-17, 9.485049e-17, 
    9.484647e-17, 9.483571e-17, 9.485476e-17, 9.479373e-17, 9.483186e-17, 
    9.488849e-17, 9.487703e-17, 9.487504e-17, 9.487954e-17, 9.484851e-17, 
    9.485978e-17, 9.482945e-17, 9.483756e-17, 9.482419e-17, 9.483086e-17, 
    9.483186e-17, 9.484036e-17, 9.484575e-17, 9.485932e-17, 9.487029e-17, 
    9.487884e-17, 9.487683e-17, 9.486743e-17, 9.485021e-17, 9.483375e-17, 
    9.483739e-17, 9.48252e-17, 9.4857e-17, 9.484379e-17, 9.484899e-17, 
    9.48354e-17, 9.48649e-17, 9.484067e-17, 9.487121e-17, 9.486847e-17, 
    9.486e-17, 9.484311e-17, 9.483893e-17, 9.483501e-17, 9.483737e-17, 
    9.484971e-17, 9.485162e-17, 9.486014e-17, 9.486264e-17, 9.486905e-17, 
    9.487449e-17, 9.486959e-17, 9.48645e-17, 9.484958e-17, 9.483634e-17, 
    9.482182e-17, 9.481816e-17, 9.480198e-17, 9.481555e-17, 9.479357e-17, 
    9.481286e-17, 9.47792e-17, 9.483882e-17, 9.481284e-17, 9.485952e-17, 
    9.48544e-17, 9.484547e-17, 9.482441e-17, 9.483546e-17, 9.48224e-17, 
    9.485167e-17, 9.486725e-17, 9.487092e-17, 9.487838e-17, 9.487075e-17, 
    9.487136e-17, 9.486408e-17, 9.48664e-17, 9.484909e-17, 9.485838e-17, 
    9.483196e-17, 9.482243e-17, 9.479521e-17, 9.477876e-17, 9.476158e-17, 
    9.475416e-17, 9.475188e-17, 9.475095e-17 ;

 MEG_pinene_a =
  8.100169e-17, 8.098464e-17, 8.098787e-17, 8.097431e-17, 8.098171e-17, 
    8.097293e-17, 8.099809e-17, 8.098409e-17, 8.099294e-17, 8.099996e-17, 
    8.094847e-17, 8.097367e-17, 8.092102e-17, 8.093726e-17, 8.089609e-17, 
    8.092373e-17, 8.089047e-17, 8.089656e-17, 8.087747e-17, 8.088291e-17, 
    8.085919e-17, 8.087494e-17, 8.084641e-17, 8.086277e-17, 8.086034e-17, 
    8.087551e-17, 8.096828e-17, 8.09517e-17, 8.096934e-17, 8.096696e-17, 
    8.096796e-17, 8.098167e-17, 8.09888e-17, 8.100277e-17, 8.100018e-17, 
    8.09898e-17, 8.096588e-17, 8.097378e-17, 8.095326e-17, 8.095372e-17, 
    8.093115e-17, 8.094132e-17, 8.090321e-17, 8.091396e-17, 8.088268e-17, 
    8.089057e-17, 8.08831e-17, 8.088533e-17, 8.088308e-17, 8.089464e-17, 
    8.08897e-17, 8.089979e-17, 8.093948e-17, 8.09279e-17, 8.096263e-17, 
    8.098406e-17, 8.099753e-17, 8.100734e-17, 8.100596e-17, 8.100338e-17, 
    8.098974e-17, 8.097667e-17, 8.096681e-17, 8.096027e-17, 8.095378e-17, 
    8.093502e-17, 8.09244e-17, 8.090119e-17, 8.09051e-17, 8.089826e-17, 
    8.089135e-17, 8.088013e-17, 8.088193e-17, 8.087705e-17, 8.089824e-17, 
    8.088425e-17, 8.09074e-17, 8.09011e-17, 8.095311e-17, 8.09716e-17, 
    8.09804e-17, 8.098729e-17, 8.100491e-17, 8.09928e-17, 8.09976e-17, 
    8.098596e-17, 8.097873e-17, 8.098225e-17, 8.096009e-17, 8.096874e-17, 
    8.092378e-17, 8.094311e-17, 8.089216e-17, 8.090427e-17, 8.088922e-17, 
    8.089684e-17, 8.088386e-17, 8.089554e-17, 8.087515e-17, 8.087083e-17, 
    8.087381e-17, 8.086205e-17, 8.089622e-17, 8.08832e-17, 8.09824e-17, 
    8.098184e-17, 8.097906e-17, 8.09913e-17, 8.099199e-17, 8.10029e-17, 
    8.099309e-17, 8.098901e-17, 8.097822e-17, 8.097205e-17, 8.096611e-17, 
    8.095306e-17, 8.093868e-17, 8.09183e-17, 8.09035e-17, 8.089366e-17, 
    8.089962e-17, 8.089436e-17, 8.090028e-17, 8.090301e-17, 8.087252e-17, 
    8.088972e-17, 8.086374e-17, 8.086514e-17, 8.087698e-17, 8.086498e-17, 
    8.098142e-17, 8.098473e-17, 8.099659e-17, 8.098731e-17, 8.100408e-17, 
    8.099482e-17, 8.098958e-17, 8.09688e-17, 8.096398e-17, 8.095985e-17, 
    8.095145e-17, 8.094081e-17, 8.092223e-17, 8.090592e-17, 8.089091e-17, 
    8.089198e-17, 8.089161e-17, 8.088837e-17, 8.089654e-17, 8.088702e-17, 
    8.088553e-17, 8.08896e-17, 8.086533e-17, 8.087224e-17, 8.086516e-17, 
    8.086964e-17, 8.098362e-17, 8.0978e-17, 8.098106e-17, 8.097538e-17, 
    8.097946e-17, 8.096161e-17, 8.095626e-17, 8.093098e-17, 8.094108e-17, 
    8.092471e-17, 8.093933e-17, 8.09368e-17, 8.092463e-17, 8.093847e-17, 
    8.090703e-17, 8.092874e-17, 8.088825e-17, 8.091031e-17, 8.088689e-17, 
    8.089097e-17, 8.088411e-17, 8.087809e-17, 8.087031e-17, 8.085631e-17, 
    8.08595e-17, 8.084763e-17, 8.096953e-17, 8.096235e-17, 8.096278e-17, 
    8.095513e-17, 8.094952e-17, 8.093712e-17, 8.091749e-17, 8.09248e-17, 
    8.091116e-17, 8.090849e-17, 8.09291e-17, 8.091664e-17, 8.095739e-17, 
    8.095101e-17, 8.095466e-17, 8.096908e-17, 8.09234e-17, 8.094694e-17, 
    8.09033e-17, 8.091599e-17, 8.087897e-17, 8.089756e-17, 8.086131e-17, 
    8.084638e-17, 8.083142e-17, 8.081506e-17, 8.095821e-17, 8.096311e-17, 
    8.095415e-17, 8.094216e-17, 8.093046e-17, 8.091526e-17, 8.091359e-17, 
    8.09108e-17, 8.090333e-17, 8.089715e-17, 8.091012e-17, 8.089559e-17, 
    8.094993e-17, 8.092127e-17, 8.096515e-17, 8.095219e-17, 8.094278e-17, 
    8.09467e-17, 8.092559e-17, 8.092069e-17, 8.090086e-17, 8.0911e-17, 
    8.085024e-17, 8.087709e-17, 8.080195e-17, 8.082302e-17, 8.096487e-17, 
    8.095813e-17, 8.093501e-17, 8.094598e-17, 8.091413e-17, 8.090639e-17, 
    8.089993e-17, 8.089202e-17, 8.089101e-17, 8.08863e-17, 8.089404e-17, 
    8.088652e-17, 8.091522e-17, 8.090235e-17, 8.093741e-17, 8.092899e-17, 
    8.093279e-17, 8.093711e-17, 8.09238e-17, 8.090996e-17, 8.090934e-17, 
    8.090495e-17, 8.089321e-17, 8.091399e-17, 8.084738e-17, 8.088901e-17, 
    8.095081e-17, 8.093831e-17, 8.093612e-17, 8.094103e-17, 8.090717e-17, 
    8.091948e-17, 8.088637e-17, 8.089523e-17, 8.088063e-17, 8.088791e-17, 
    8.0889e-17, 8.089828e-17, 8.090416e-17, 8.091898e-17, 8.093095e-17, 
    8.094028e-17, 8.093808e-17, 8.092782e-17, 8.090904e-17, 8.089107e-17, 
    8.089504e-17, 8.088173e-17, 8.091645e-17, 8.090204e-17, 8.09077e-17, 
    8.089287e-17, 8.092506e-17, 8.089863e-17, 8.093195e-17, 8.092896e-17, 
    8.091972e-17, 8.090128e-17, 8.089672e-17, 8.089245e-17, 8.089502e-17, 
    8.090849e-17, 8.091057e-17, 8.091986e-17, 8.09226e-17, 8.092958e-17, 
    8.093553e-17, 8.093018e-17, 8.092463e-17, 8.090836e-17, 8.08939e-17, 
    8.087805e-17, 8.087404e-17, 8.085638e-17, 8.08712e-17, 8.084721e-17, 
    8.086827e-17, 8.08315e-17, 8.089661e-17, 8.086825e-17, 8.091919e-17, 
    8.091361e-17, 8.090386e-17, 8.088088e-17, 8.089294e-17, 8.087868e-17, 
    8.091063e-17, 8.092763e-17, 8.093164e-17, 8.093977e-17, 8.093145e-17, 
    8.093211e-17, 8.092417e-17, 8.09267e-17, 8.090781e-17, 8.091794e-17, 
    8.088911e-17, 8.08787e-17, 8.084899e-17, 8.083102e-17, 8.081226e-17, 
    8.080415e-17, 8.080166e-17, 8.080064e-17 ;

 MEG_thujene_a =
  1.951996e-18, 1.951614e-18, 1.951687e-18, 1.951384e-18, 1.951549e-18, 
    1.951353e-18, 1.951915e-18, 1.951602e-18, 1.9518e-18, 1.951957e-18, 
    1.950806e-18, 1.951369e-18, 1.950192e-18, 1.950555e-18, 1.949635e-18, 
    1.950253e-18, 1.949509e-18, 1.949645e-18, 1.949218e-18, 1.94934e-18, 
    1.94881e-18, 1.949162e-18, 1.948524e-18, 1.94889e-18, 1.948835e-18, 
    1.949175e-18, 1.951249e-18, 1.950878e-18, 1.951273e-18, 1.951219e-18, 
    1.951242e-18, 1.951548e-18, 1.951707e-18, 1.95202e-18, 1.951962e-18, 
    1.95173e-18, 1.951195e-18, 1.951372e-18, 1.950913e-18, 1.950923e-18, 
    1.950418e-18, 1.950646e-18, 1.949794e-18, 1.950034e-18, 1.949335e-18, 
    1.949511e-18, 1.949344e-18, 1.949394e-18, 1.949344e-18, 1.949602e-18, 
    1.949492e-18, 1.949717e-18, 1.950605e-18, 1.950346e-18, 1.951122e-18, 
    1.951601e-18, 1.951903e-18, 1.952122e-18, 1.952091e-18, 1.952033e-18, 
    1.951729e-18, 1.951436e-18, 1.951216e-18, 1.95107e-18, 1.950924e-18, 
    1.950505e-18, 1.950268e-18, 1.949749e-18, 1.949836e-18, 1.949683e-18, 
    1.949529e-18, 1.949278e-18, 1.949318e-18, 1.949209e-18, 1.949683e-18, 
    1.94937e-18, 1.949887e-18, 1.949747e-18, 1.950909e-18, 1.951323e-18, 
    1.95152e-18, 1.951674e-18, 1.952068e-18, 1.951797e-18, 1.951904e-18, 
    1.951644e-18, 1.951482e-18, 1.951561e-18, 1.951066e-18, 1.951259e-18, 
    1.950254e-18, 1.950686e-18, 1.949547e-18, 1.949818e-18, 1.949481e-18, 
    1.949651e-18, 1.949361e-18, 1.949622e-18, 1.949167e-18, 1.94907e-18, 
    1.949137e-18, 1.948874e-18, 1.949638e-18, 1.949347e-18, 1.951565e-18, 
    1.951552e-18, 1.95149e-18, 1.951763e-18, 1.951779e-18, 1.952023e-18, 
    1.951803e-18, 1.951712e-18, 1.951471e-18, 1.951333e-18, 1.9512e-18, 
    1.950908e-18, 1.950587e-18, 1.950131e-18, 1.9498e-18, 1.94958e-18, 
    1.949714e-18, 1.949596e-18, 1.949728e-18, 1.949789e-18, 1.949108e-18, 
    1.949492e-18, 1.948912e-18, 1.948943e-18, 1.949207e-18, 1.948939e-18, 
    1.951542e-18, 1.951616e-18, 1.951882e-18, 1.951674e-18, 1.952049e-18, 
    1.951842e-18, 1.951725e-18, 1.95126e-18, 1.951152e-18, 1.95106e-18, 
    1.950872e-18, 1.950635e-18, 1.950219e-18, 1.949855e-18, 1.949519e-18, 
    1.949543e-18, 1.949535e-18, 1.949462e-18, 1.949645e-18, 1.949432e-18, 
    1.949399e-18, 1.94949e-18, 1.948947e-18, 1.949102e-18, 1.948944e-18, 
    1.949043e-18, 1.951592e-18, 1.951466e-18, 1.951534e-18, 1.951407e-18, 
    1.951499e-18, 1.951099e-18, 1.95098e-18, 1.950415e-18, 1.950641e-18, 
    1.950275e-18, 1.950601e-18, 1.950545e-18, 1.950273e-18, 1.950582e-18, 
    1.949879e-18, 1.950365e-18, 1.949459e-18, 1.949953e-18, 1.949429e-18, 
    1.94952e-18, 1.949367e-18, 1.949232e-18, 1.949059e-18, 1.948745e-18, 
    1.948817e-18, 1.948552e-18, 1.951277e-18, 1.951116e-18, 1.951126e-18, 
    1.950955e-18, 1.950829e-18, 1.950552e-18, 1.950113e-18, 1.950277e-18, 
    1.949972e-18, 1.949912e-18, 1.950373e-18, 1.950094e-18, 1.951005e-18, 
    1.950863e-18, 1.950944e-18, 1.951267e-18, 1.950245e-18, 1.950771e-18, 
    1.949796e-18, 1.95008e-18, 1.949252e-18, 1.949668e-18, 1.948857e-18, 
    1.948524e-18, 1.948189e-18, 1.947824e-18, 1.951024e-18, 1.951133e-18, 
    1.950933e-18, 1.950665e-18, 1.950403e-18, 1.950063e-18, 1.950026e-18, 
    1.949964e-18, 1.949796e-18, 1.949658e-18, 1.949948e-18, 1.949624e-18, 
    1.950838e-18, 1.950198e-18, 1.951179e-18, 1.950889e-18, 1.950679e-18, 
    1.950766e-18, 1.950294e-18, 1.950185e-18, 1.949741e-18, 1.949968e-18, 
    1.94861e-18, 1.94921e-18, 1.947531e-18, 1.948001e-18, 1.951172e-18, 
    1.951022e-18, 1.950505e-18, 1.95075e-18, 1.950038e-18, 1.949865e-18, 
    1.949721e-18, 1.949544e-18, 1.949521e-18, 1.949416e-18, 1.949589e-18, 
    1.949421e-18, 1.950062e-18, 1.949775e-18, 1.950558e-18, 1.95037e-18, 
    1.950455e-18, 1.950552e-18, 1.950254e-18, 1.949945e-18, 1.949931e-18, 
    1.949833e-18, 1.94957e-18, 1.950035e-18, 1.948546e-18, 1.949477e-18, 
    1.950858e-18, 1.950579e-18, 1.95053e-18, 1.95064e-18, 1.949882e-18, 
    1.950157e-18, 1.949417e-18, 1.949615e-18, 1.949289e-18, 1.949452e-18, 
    1.949476e-18, 1.949684e-18, 1.949815e-18, 1.950146e-18, 1.950414e-18, 
    1.950623e-18, 1.950574e-18, 1.950344e-18, 1.949924e-18, 1.949522e-18, 
    1.949611e-18, 1.949314e-18, 1.95009e-18, 1.949768e-18, 1.949894e-18, 
    1.949563e-18, 1.950283e-18, 1.949691e-18, 1.950436e-18, 1.950369e-18, 
    1.950163e-18, 1.949751e-18, 1.949649e-18, 1.949553e-18, 1.949611e-18, 
    1.949912e-18, 1.949958e-18, 1.950166e-18, 1.950227e-18, 1.950384e-18, 
    1.950516e-18, 1.950397e-18, 1.950273e-18, 1.949909e-18, 1.949586e-18, 
    1.949231e-18, 1.949142e-18, 1.948747e-18, 1.949078e-18, 1.948542e-18, 
    1.949013e-18, 1.948191e-18, 1.949646e-18, 1.949012e-18, 1.950151e-18, 
    1.950026e-18, 1.949808e-18, 1.949295e-18, 1.949564e-18, 1.949246e-18, 
    1.94996e-18, 1.95034e-18, 1.950429e-18, 1.950611e-18, 1.950425e-18, 
    1.95044e-18, 1.950263e-18, 1.950319e-18, 1.949897e-18, 1.950123e-18, 
    1.949479e-18, 1.949246e-18, 1.948582e-18, 1.94818e-18, 1.947761e-18, 
    1.94758e-18, 1.947524e-18, 1.947501e-18 ;

 MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 M_LITR1C_TO_LEACHING =
  -5.329227e-25, -1.648206e-26, -1.758095e-25, -1.867976e-25, -1.483393e-25, 
    -2.637143e-25, -4.450179e-25, 1.977859e-25, -1.538333e-25, 1.04387e-25, 
    -3.516191e-25, 2.747033e-26, -4.944636e-26, 9.339893e-26, -6.043446e-26, 
    8.241083e-26, -1.428452e-25, -3.131607e-25, 2.747026e-25, -3.351369e-25, 
    2.472323e-25, 3.626074e-25, -1.703155e-25, -2.142678e-25, 1.538335e-25, 
    -4.450179e-25, -1.15375e-25, -3.296429e-25, 3.845843e-26, -5.493964e-27, 
    4.395241e-25, 3.18655e-25, -1.098809e-25, 1.648216e-25, 1.153751e-25, 
    2.362442e-25, -3.296421e-26, -2.032797e-25, -1.648214e-25, -4.724882e-25, 
    -1.098801e-26, 5.494135e-27, 7.142273e-26, -4.395239e-25, 3.076669e-25, 
    -5.494041e-26, 1.703156e-25, 2.252561e-25, -2.527262e-25, 2.747033e-26, 
    1.098819e-26, 1.593275e-25, -3.955715e-25, -3.790893e-25, -3.955715e-25, 
    -3.790893e-25, -7.691661e-26, 2.032799e-25, -1.483393e-25, 7.691678e-26, 
    3.571133e-25, 9.339893e-26, -1.428452e-25, -1.758095e-25, 2.747033e-26, 
    6.592868e-26, 1.813037e-25, 1.977859e-25, -5.493964e-27, -1.20869e-25, 
    5.988515e-25, -3.46125e-25, 5.494135e-27, 5.494058e-26, -3.516191e-25, 
    -3.845834e-25, -1.922916e-25, 3.076669e-25, -7.142256e-26, 1.098811e-25, 
    -1.428452e-25, -4.010655e-25, -7.691661e-26, 3.626074e-25, 5.109467e-25, 
    4.010657e-25, 8.590251e-32, 1.318573e-25, -4.065596e-25, 6.53792e-25, 
    -1.648206e-26, 1.153751e-25, 4.395248e-26, 6.592868e-26, -6.043446e-26, 
    -1.15375e-25, -6.592851e-26, -3.131607e-25, -6.043446e-26, -3.351369e-25, 
    2.197628e-26, -1.593273e-25, 1.318573e-25, 2.197628e-26, 5.109467e-25, 
    -2.032797e-25, 2.197628e-26, 2.197621e-25, -1.648214e-25, -3.40631e-25, 
    -1.758095e-25, 1.703156e-25, 2.637145e-25, 9.339893e-26, -3.845826e-26, 
    9.339893e-26, 2.582204e-25, -1.15375e-25, 3.021728e-25, -3.076667e-25, 
    9.339893e-26, 3.626074e-25, -1.098809e-25, -3.681012e-25, -4.395231e-26, 
    -2.966786e-25, -2.747016e-26, -3.186548e-25, 3.516193e-25, 2.307502e-25, 
    -2.692083e-25, -2.142678e-25, 2.582204e-25, -1.373511e-25, 2.032799e-25, 
    1.648216e-25, 1.208692e-25, -6.373097e-25, -7.142256e-26, 2.307502e-25, 
    5.384169e-25, 2.856907e-25, -1.977857e-25, -2.692083e-25, -2.637143e-25, 
    -3.681012e-25, -2.197611e-26, 2.032799e-25, 5.494058e-26, -2.087738e-25, 
    -1.648214e-25, -2.856905e-25, -2.472321e-25, -5.384167e-25, 
    -3.296429e-25, -1.648206e-26, 7.691678e-26, -2.36244e-25, -3.076667e-25, 
    1.593275e-25, -2.417381e-25, -1.922916e-25, -1.813035e-25, 8.590151e-32, 
    2.911847e-25, -2.747024e-25, 1.922918e-25, -6.043446e-26, 1.593275e-25, 
    -4.889703e-25, 3.076669e-25, -1.428452e-25, 5.494135e-27, 4.3403e-25, 
    4.944653e-26, 4.395248e-26, -1.703155e-25, -3.186548e-25, -8.790471e-26, 
    -6.043446e-26, 4.669943e-25, 1.098819e-26, 2.197621e-25, 9.889298e-26, 
    -1.043869e-25, 3.516193e-25, 1.208692e-25, 1.922918e-25, 1.977859e-25, 
    -2.747016e-26, -5.768751e-25, 1.977859e-25, -6.592851e-26, 1.483394e-25, 
    -4.724882e-25, -5.494049e-25, -2.801964e-25, 2.032799e-25, -1.538333e-25, 
    2.527264e-25, -3.845826e-26, -4.944644e-25, -2.417381e-25, -1.703155e-25, 
    4.395248e-26, -3.46125e-25, -2.3075e-25, 1.483394e-25, 1.867978e-25, 
    1.263632e-25, 5.494058e-26, -6.592851e-26, 1.208692e-25, -1.20869e-25, 
    1.648223e-26, -3.735953e-25, 2.252561e-25, 1.593275e-25, 6.592868e-26, 
    2.747026e-25, -6.043446e-26, -2.197619e-25, 1.648223e-26, 1.153751e-25, 
    -2.197611e-26, 2.801966e-25, 4.944653e-26, 1.648216e-25, 2.856907e-25, 
    5.164408e-25, -2.966786e-25, 5.494058e-26, 2.582204e-25, -4.615001e-25, 
    -2.197619e-25, -2.527262e-25, -8.241066e-26, 3.681014e-25, 5.494135e-27, 
    -2.417381e-25, -2.3075e-25, 2.747026e-25, 1.538335e-25, 1.04387e-25, 
    1.648223e-26, 2.856907e-25, -1.15375e-25, -4.669941e-25, -2.25256e-25, 
    7.691678e-26, -2.966786e-25, -1.098801e-26, 3.076669e-25, 2.307502e-25, 
    -5.493964e-27, 1.813037e-25, 3.845843e-26, 8.790488e-26, 1.648223e-26, 
    -2.747016e-26, 1.318573e-25, -2.966786e-25, -4.944636e-26, -2.801964e-25, 
    1.318573e-25, 4.395248e-26, -1.648206e-26, 7.691678e-26, 1.263632e-25, 
    3.406311e-25, 2.197621e-25, -1.098801e-26, -3.186548e-25, -1.977857e-25, 
    -1.098809e-25, -6.043446e-26, -6.592851e-26, -5.494041e-26, 
    -2.747016e-26, -1.098801e-26, -1.20869e-25, 2.801966e-25, -2.472321e-25, 
    -2.472321e-25, -3.351369e-25, 3.681014e-25, 5.713812e-25, -2.801964e-25, 
    -1.813035e-25, -2.36244e-25, -5.60393e-25, -1.648214e-25, 1.483394e-25, 
    4.120538e-25, -1.593273e-25, 5.768753e-25, 3.296438e-26, -4.230417e-25, 
    -1.648214e-25, -1.648206e-26, 7.856492e-25, 1.813037e-25, -4.120536e-25, 
    -2.527262e-25, -5.493964e-27, -2.087738e-25, 8.241083e-26, -4.944644e-25, 
    1.318573e-25, 3.296438e-26, 1.263632e-25, -2.032797e-25, 1.922918e-25, 
    -6.043446e-26, -1.648206e-26, -2.527262e-25, 3.131609e-25, -4.724882e-25, 
    8.590074e-32, -1.703155e-25, -2.197611e-26, -2.032797e-25, 8.590154e-32, 
    1.153751e-25, -2.3075e-25, -2.197619e-25, 2.032799e-25, -1.263631e-25, 
    1.208692e-25, -1.813035e-25, 2.692085e-25, -2.856905e-25, 7.691678e-26, 
    -1.593273e-25, -1.703155e-25, -1.648206e-26, 1.318573e-25, -1.648206e-26 ;

 M_LITR2C_TO_LEACHING =
  -8.790474e-26, 1.64822e-26, 5.494105e-27, 1.318572e-25, 2.74703e-26, 
    1.593275e-25, -2.197619e-25, -3.021727e-25, -3.296429e-25, 1.318572e-25, 
    1.04387e-25, 8.790485e-26, -1.648209e-26, 2.307501e-25, 9.889295e-26, 
    6.04346e-26, -1.373512e-25, 8.790485e-26, -9.889284e-26, -2.087738e-25, 
    3.29643e-25, 6.04346e-26, -7.142259e-26, -8.790474e-26, 2.74703e-26, 
    -2.197614e-26, 2.252561e-25, 2.362442e-25, 2.032799e-25, -1.098804e-26, 
    5.494105e-27, -1.098809e-25, -4.944639e-26, -6.592854e-26, -2.087738e-25, 
    -3.021727e-25, -1.373512e-25, -1.648209e-26, -9.889284e-26, 1.977858e-25, 
    1.098815e-26, 3.131609e-25, 3.296435e-26, -3.40631e-25, -1.648209e-26, 
    -8.241069e-26, 5.494055e-26, 1.373513e-25, -6.043449e-26, 1.813037e-25, 
    -1.758095e-25, -6.592854e-26, -3.296424e-26, -1.758095e-25, 
    -3.076667e-25, 1.758096e-25, 1.867977e-25, -1.648209e-26, -2.362441e-25, 
    1.428453e-25, 1.318572e-25, -2.142679e-25, 1.703156e-25, -8.790474e-26, 
    -6.043449e-26, -1.758095e-25, -5.494044e-26, -3.845829e-26, 1.483394e-25, 
    -3.296429e-25, 6.04346e-26, 1.04387e-25, -3.296424e-26, -2.527262e-25, 
    -9.889284e-26, -1.318571e-25, -2.747024e-25, -3.35137e-25, 4.395245e-26, 
    -7.142259e-26, 3.131609e-25, 1.813037e-25, -5.493994e-27, 3.571133e-25, 
    -3.131608e-25, 1.813037e-25, -3.900775e-25, -1.20869e-25, -9.339879e-26, 
    3.296435e-26, 3.84584e-26, 4.94465e-26, 1.318572e-25, -1.263631e-25, 
    -2.417381e-25, -6.043449e-26, -4.944639e-26, 1.648215e-25, -1.648214e-25, 
    -8.241069e-26, -1.703155e-25, 2.527263e-25, -5.493994e-27, 1.208691e-25, 
    5.562093e-32, 1.977858e-25, -2.582203e-25, 3.021728e-25, -1.373512e-25, 
    -1.263631e-25, 8.24108e-26, -2.692084e-25, -1.318571e-25, -2.087738e-25, 
    -1.428452e-25, 1.64822e-26, -2.087738e-25, -1.043869e-25, -1.098804e-26, 
    -7.691664e-26, -1.648209e-26, -1.263631e-25, -3.296424e-26, 1.318572e-25, 
    -4.944639e-26, -3.296424e-26, -1.15375e-25, 1.318572e-25, -1.648214e-25, 
    -4.395234e-26, -1.813036e-25, 2.74703e-26, -5.494044e-26, -1.483393e-25, 
    1.648215e-25, 1.098811e-25, 1.153751e-25, 1.648215e-25, -3.131608e-25, 
    1.373513e-25, -1.483393e-25, -8.790474e-26, -1.428452e-25, -8.241069e-26, 
    5.494055e-26, 1.373513e-25, 1.867977e-25, 4.39524e-25, -8.241069e-26, 
    -3.845829e-26, -1.813036e-25, 3.296435e-26, 3.296435e-26, 2.856906e-25, 
    -1.867976e-25, -4.340298e-25, -5.493994e-27, 1.153751e-25, 7.691675e-26, 
    -3.241489e-25, -2.747019e-26, 5.494105e-27, -9.889284e-26, -2.747019e-26, 
    -2.692084e-25, -1.263631e-25, 9.889295e-26, -1.373512e-25, 1.593275e-25, 
    -4.944639e-26, -8.241069e-26, 9.33989e-26, 5.562061e-32, -6.043449e-26, 
    1.373513e-25, -1.922917e-25, -5.494044e-26, 1.428453e-25, -3.296429e-25, 
    5.494105e-27, -7.142259e-26, 2.19762e-25, -9.889284e-26, -4.285358e-25, 
    1.428453e-25, -1.813036e-25, -1.20869e-25, -1.538333e-25, 2.74703e-26, 
    -2.747019e-26, 6.04346e-26, -7.142259e-26, -3.900775e-25, -2.417381e-25, 
    -1.593274e-25, -1.098804e-26, 1.098815e-26, 2.197625e-26, -1.648209e-26, 
    7.14227e-26, -1.20869e-25, -6.043449e-26, 7.691675e-26, -2.637143e-25, 
    1.04387e-25, -1.043869e-25, 3.735954e-25, 1.538334e-25, -1.20869e-25, 
    4.94465e-26, 2.252561e-25, 1.977858e-25, -4.944639e-26, 3.516192e-25, 
    2.197625e-26, -7.691664e-26, 8.24108e-26, 2.197625e-26, -3.296424e-26, 
    9.33989e-26, 2.417382e-25, 7.691675e-26, 1.483394e-25, -1.813036e-25, 
    -1.813036e-25, -2.197614e-26, -1.098804e-26, -1.098804e-26, 9.33989e-26, 
    -3.131608e-25, 1.153751e-25, 2.197625e-26, 1.483394e-25, 7.691675e-26, 
    7.691675e-26, 1.64822e-26, -2.197614e-26, -2.197619e-25, -1.483393e-25, 
    2.307501e-25, -1.263631e-25, -1.538333e-25, 1.64822e-26, -2.3075e-25, 
    -1.098804e-26, -7.691664e-26, 1.373513e-25, 5.494055e-26, -1.098804e-26, 
    -1.098809e-25, -1.593274e-25, 7.691675e-26, 8.790485e-26, -9.889284e-26, 
    2.417382e-25, -1.043869e-25, 6.592865e-26, -2.197614e-26, 1.483394e-25, 
    8.790485e-26, 1.758096e-25, 7.691675e-26, -5.494044e-26, -2.472322e-25, 
    -2.527262e-25, 3.461252e-25, -1.098804e-26, 1.208691e-25, -1.867976e-25, 
    -2.472322e-25, 1.758096e-25, 8.24108e-26, -1.483393e-25, -2.362441e-25, 
    -1.813036e-25, 6.04346e-26, -1.428452e-25, -1.703155e-25, 1.04387e-25, 
    1.813037e-25, -1.593274e-25, -9.339879e-26, 6.04346e-26, 2.74703e-26, 
    -8.241069e-26, -1.373512e-25, -3.461251e-25, 1.977858e-25, -9.339879e-26, 
    1.593275e-25, -2.3075e-25, 1.428453e-25, -2.692084e-25, 6.04346e-26, 
    -4.944639e-26, -3.296429e-25, -2.747019e-26, 3.84584e-26, -3.296424e-26, 
    -7.142259e-26, 1.153751e-25, -2.911846e-25, 5.562073e-32, -1.428452e-25, 
    -2.032798e-25, 5.562057e-32, 2.252561e-25, 7.691675e-26, 3.84584e-26, 
    1.428453e-25, 2.087739e-25, 1.64822e-26, -1.977857e-25, -7.142259e-26, 
    9.889295e-26, 1.263632e-25, -1.648214e-25, -1.318571e-25, -1.15375e-25, 
    2.032799e-25, -2.032798e-25, -2.747019e-26, -2.087738e-25, 4.94465e-26, 
    -3.900775e-25, -1.538333e-25, 1.922918e-25, 2.472323e-25, -1.098804e-26, 
    -1.867976e-25, -2.966786e-25, -7.691664e-26, -4.889704e-25, 5.494055e-26, 
    2.856906e-25, -1.043869e-25, 8.790485e-26, -3.296424e-26 ;

 M_LITR3C_TO_LEACHING =
  -3.845832e-26, -5.494047e-26, -6.318154e-26, -7.966369e-26, -2.746997e-27, 
    4.944647e-26, -6.867559e-26, 4.669945e-26, -6.318154e-26, -2.47232e-26, 
    -8.241047e-27, -9.614584e-26, -1.236161e-25, -1.648212e-26, 2.664614e-25, 
    -6.318154e-26, 1.12628e-25, -1.37351e-26, -5.768749e-26, -5.494022e-27, 
    3.845837e-26, 1.153751e-25, -7.691667e-26, 4.944647e-26, 2.197623e-26, 
    -9.065179e-26, -4.944642e-26, -7.416964e-26, 8.241102e-27, 6.867565e-26, 
    -1.758096e-25, -7.416964e-26, -7.416964e-26, -1.620744e-25, 1.208691e-25, 
    -8.515774e-26, -5.494047e-26, 7.691672e-26, 2.664614e-25, 9.339887e-26, 
    -3.57113e-26, -1.263631e-25, 2.747052e-27, 3.845837e-26, -4.120535e-26, 
    4.669945e-26, 5.494053e-26, 1.373515e-26, 7.416969e-26, -6.318154e-26, 
    -1.346042e-25, 1.92292e-26, -1.922915e-26, 6.867565e-26, -2.47232e-26, 
    6.592862e-26, -1.455923e-25, -3.57113e-26, -8.241047e-27, 1.648218e-26, 
    -1.15375e-25, 1.07134e-25, 9.065185e-26, -1.867977e-25, 8.515779e-26, 
    8.515779e-26, -8.241047e-27, 1.373515e-26, -2.747022e-26, -9.065179e-26, 
    -1.071339e-25, -5.494022e-27, 4.669945e-26, -3.57113e-26, -6.867559e-26, 
    1.373515e-26, 5.494053e-26, -6.043452e-26, -3.296427e-26, 4.669945e-26, 
    -2.747022e-26, -8.515774e-26, 7.142267e-26, -6.318154e-26, 4.395242e-26, 
    -3.021725e-26, -1.455923e-25, -9.339881e-26, -6.318154e-26, 
    -1.922915e-26, -1.098807e-26, 1.648218e-26, 1.07134e-25, 5.21935e-26, 
    1.648218e-26, -8.241047e-27, -1.922915e-26, 8.515779e-26, -1.648212e-26, 
    2.280031e-25, 1.483394e-25, -8.790477e-26, 1.098813e-26, 1.318572e-25, 
    -1.098807e-26, -6.867559e-26, -9.889287e-26, -1.648212e-26, 9.339887e-26, 
    -6.318154e-26, 1.813037e-25, -8.241047e-27, -7.416964e-26, 7.142267e-26, 
    -2.47232e-26, -8.515774e-26, 5.494053e-26, -5.768749e-26, -1.098807e-26, 
    1.373515e-26, -1.043869e-25, 7.416969e-26, -1.208691e-25, 1.813037e-25, 
    -7.142262e-26, -2.747022e-26, -6.318154e-26, -4.669939e-26, 
    -1.071339e-25, -1.12628e-25, -5.494022e-27, 4.12054e-26, 3.845837e-26, 
    -1.37351e-26, 1.098813e-26, 1.92292e-26, -7.416964e-26, -6.592857e-26, 
    6.043457e-26, 4.12054e-26, -1.922917e-25, -5.494047e-26, 7.966375e-26, 
    -4.120535e-26, 6.592862e-26, 1.098813e-26, -2.47232e-26, -9.614584e-26, 
    5.494077e-27, -2.47232e-26, -3.296427e-26, -8.241071e-26, 8.790482e-26, 
    -8.241071e-26, -2.47232e-26, -4.395237e-26, 1.318572e-25, -1.09881e-25, 
    -1.483393e-25, 6.592862e-26, -7.691667e-26, 1.675685e-25, -7.142262e-26, 
    -9.889287e-26, 2.747052e-27, 8.241102e-27, -1.538334e-25, -6.043452e-26, 
    1.538334e-25, 3.02173e-26, -2.747022e-26, 8.241102e-27, -1.346042e-25, 
    -7.691667e-26, -1.538334e-25, 2.472325e-26, -6.318154e-26, 1.373515e-26, 
    -2.197617e-26, 2.781024e-32, 6.31816e-26, -3.57113e-26, -2.197617e-26, 
    -1.016399e-25, 3.296432e-26, 5.494053e-26, -1.840506e-25, -5.219344e-26, 
    -1.37351e-26, -1.18122e-25, -1.016399e-25, -6.592857e-26, -9.889287e-26, 
    9.065185e-26, 2.747028e-26, -5.219344e-26, 1.373515e-26, -3.021725e-26, 
    -5.219344e-26, -3.296427e-26, 5.494077e-27, -7.142262e-26, 2.747028e-26, 
    -4.944642e-26, 8.241077e-26, -1.37351e-26, 1.098813e-26, -7.691667e-26, 
    -3.845832e-26, 3.571135e-26, -2.032798e-25, -9.065179e-26, -2.746997e-27, 
    8.241077e-26, 6.592862e-26, 2.781033e-32, -8.241071e-26, -5.494022e-27, 
    -5.219344e-26, 2.781031e-32, -7.966369e-26, -1.12628e-25, -1.12628e-25, 
    5.494077e-27, -9.614584e-26, -2.747022e-26, -9.065179e-26, -6.867559e-26, 
    -1.291101e-25, -5.494022e-27, -1.263631e-25, -9.339881e-26, 2.781015e-32, 
    -7.142262e-26, 6.043457e-26, -6.867559e-26, 1.593275e-25, -3.296427e-26, 
    4.395242e-26, -7.416964e-26, 2.472325e-26, 2.747028e-26, -8.241071e-26, 
    6.043457e-26, -2.032798e-25, -3.845832e-26, -1.538334e-25, -6.867559e-26, 
    2.747052e-27, -4.120535e-26, 7.966375e-26, 7.691672e-26, -4.395237e-26, 
    -1.648212e-26, -1.15375e-25, -3.296427e-26, -7.416964e-26, -1.922915e-26, 
    -1.373512e-25, -8.241071e-26, 4.12054e-26, 2.747052e-27, -4.944642e-26, 
    -2.197617e-26, 1.373513e-25, -8.790477e-26, -1.37351e-26, -3.845832e-26, 
    5.494077e-27, -8.241071e-26, 7.416969e-26, -2.197617e-26, -1.071339e-25, 
    2.472325e-26, 2.781037e-32, -3.021725e-26, 1.236161e-25, 8.515779e-26, 
    -8.515774e-26, -2.829435e-25, -1.648212e-26, 2.747028e-26, -3.57113e-26, 
    -2.747022e-26, 3.296432e-26, 1.016399e-25, 2.747052e-27, -3.021725e-26, 
    -1.263631e-25, -9.889287e-26, -9.339881e-26, 3.571135e-26, -2.746997e-27, 
    -1.922917e-25, 4.944647e-26, -1.455923e-25, 1.510864e-25, -3.57113e-26, 
    -1.565804e-25, -1.455923e-25, -6.318154e-26, 4.944647e-26, -6.592857e-26, 
    1.098813e-26, -3.296427e-26, 6.31816e-26, 1.373515e-26, -4.944642e-26, 
    1.400983e-25, 1.373515e-26, -1.400982e-25, -8.241047e-27, -7.691667e-26, 
    9.065185e-26, 1.09881e-25, 3.02173e-26, 6.867565e-26, 9.889292e-26, 
    -7.966369e-26, -4.944642e-26, -7.966369e-26, 2.781036e-32, -2.47232e-26, 
    6.043457e-26, -1.37351e-26, 1.92292e-26, 1.098813e-26, -9.065179e-26, 
    6.31816e-26, -3.57113e-26, -4.120535e-26, 9.065185e-26, -1.09881e-25, 
    -7.966369e-26, -3.021725e-26, -1.675685e-25, -9.889287e-26, -7.142262e-26 ;

 M_SOIL1C_TO_LEACHING =
  5.486405e-21, -1.063493e-20, 3.763798e-20, 5.013102e-21, 7.461537e-21, 
    5.161253e-21, -1.253742e-20, -1.340512e-20, 3.120472e-20, 2.678875e-20, 
    -2.732027e-20, 2.596458e-20, 3.272605e-21, -5.106293e-22, 1.977983e-20, 
    -8.194382e-21, -2.183275e-20, 2.520122e-20, -1.976007e-20, -1.674727e-20, 
    -2.248643e-20, 1.815617e-20, -5.027829e-20, -2.376156e-20, 5.202416e-20, 
    2.076362e-21, 3.055492e-21, 2.304312e-20, -2.684529e-20, -1.797574e-20, 
    1.999753e-20, -2.557356e-20, -2.537962e-20, 2.290978e-21, -1.923814e-20, 
    6.096531e-21, -1.695564e-20, -3.018575e-20, 4.938465e-21, 3.044532e-20, 
    1.519821e-20, -2.155089e-20, 1.585843e-21, 1.249416e-20, 5.259086e-21, 
    2.038374e-20, 6.514212e-22, -3.141591e-20, -2.737201e-20, 7.07873e-21, 
    1.343962e-20, 2.530453e-21, -3.717062e-20, -3.925915e-20, 6.482189e-21, 
    3.096467e-20, -3.231274e-20, 1.346448e-20, 3.158669e-20, 1.951435e-20, 
    -8.190414e-21, 8.310282e-21, 4.225142e-21, -4.136935e-21, -6.059776e-21, 
    -4.72364e-20, -7.704147e-21, 1.245514e-20, 4.567226e-21, 2.288253e-20, 
    1.995232e-20, 2.037189e-20, -1.013194e-20, 2.473045e-20, -5.810674e-21, 
    -8.498616e-21, 1.579901e-20, -4.545012e-20, -9.287999e-21, -2.32187e-20, 
    1.828477e-20, 7.904868e-21, 2.531997e-20, 3.132432e-20, 1.105281e-20, 
    1.90552e-20, -3.870698e-20, -3.514766e-20, -8.616795e-21, -2.409941e-20, 
    1.719512e-20, 4.80898e-21, 1.121989e-20, -4.066601e-20, -1.791809e-20, 
    -6.51421e-22, -1.290299e-20, -1.828137e-20, 5.022346e-20, 2.295493e-20, 
    -2.69516e-20, -9.304948e-21, -1.059591e-20, -1.099824e-20, 3.357709e-21, 
    -1.901847e-20, -1.544077e-20, 1.785727e-20, -4.057753e-20, 1.324678e-20, 
    -3.008088e-20, 9.816536e-22, 7.723637e-21, -5.596084e-21, 1.251987e-20, 
    1.740181e-20, -1.677359e-20, 3.987325e-20, -2.19454e-21, 4.33514e-20, 
    2.313925e-20, 1.754231e-20, -1.460326e-21, 5.90631e-22, -2.683792e-20, 
    6.880256e-21, -2.29125e-20, -1.137962e-20, -4.144608e-20, 1.456375e-20, 
    7.710345e-21, 3.794727e-20, 8.558257e-21, -2.569544e-20, -1.506964e-22, 
    -8.066259e-22, 2.248812e-20, -1.389903e-20, 9.236842e-21, -3.710218e-20, 
    1.085741e-20, 1.891695e-20, -1.061366e-21, -2.932682e-20, 2.124129e-20, 
    4.667178e-20, -3.007633e-20, -4.459514e-21, 2.014994e-20, 8.137272e-21, 
    1.911343e-20, 1.413003e-20, 2.762365e-20, -1.407009e-20, 1.48609e-20, 
    -6.991085e-21, -3.061691e-20, 1.982395e-20, -2.0211e-20, 3.121376e-20, 
    -1.189337e-20, 1.44389e-21, -2.501518e-20, 1.399575e-20, -6.325817e-21, 
    3.023919e-20, -2.174964e-20, -2.170835e-20, 1.786847e-21, 3.172608e-20, 
    -1.883638e-20, -1.351962e-20, -3.147727e-20, -1.349531e-20, 3.951359e-20, 
    -7.300962e-21, -1.624089e-20, -9.668544e-21, 2.692614e-20, 2.606184e-20, 
    1.72135e-20, -2.122403e-20, -1.613997e-20, -1.789403e-20, -1.350717e-20, 
    -7.34024e-21, -5.839812e-21, 3.001131e-20, 2.227466e-20, 3.118462e-20, 
    -2.716365e-20, -9.49071e-21, -4.296828e-20, -9.297878e-21, 4.005108e-20, 
    -1.943264e-20, 1.195524e-20, -1.61636e-21, 4.994431e-21, -7.475122e-21, 
    -3.362292e-20, 1.039854e-20, 2.939551e-20, -1.345795e-21, 1.422672e-20, 
    -1.768281e-20, -6.641352e-21, 5.278036e-21, 7.097107e-21, -1.611283e-20, 
    3.440297e-20, -9.722559e-21, 2.488512e-20, 4.12757e-21, 4.234759e-21, 
    3.784635e-20, -6.504502e-21, 6.589328e-21, 2.400751e-20, -2.774704e-21, 
    2.598466e-20, -1.205549e-21, -2.332869e-20, -1.94708e-20, -1.999445e-20, 
    -1.181222e-20, -2.234675e-20, -4.292441e-21, -2.824188e-21, -4.06624e-21, 
    3.459296e-20, -1.180689e-21, -1.675194e-21, 2.612745e-20, -1.24639e-20, 
    3.581946e-20, 2.057984e-21, 1.282465e-21, -1.54928e-20, -5.05729e-20, 
    -8.386936e-21, -3.551805e-20, 3.361677e-21, 2.1547e-21, 2.456932e-20, 
    -1.683604e-20, -5.625795e-21, 8.458717e-21, 2.889282e-20, 1.25866e-20, 
    -1.822737e-20, 1.544869e-20, -6.706111e-21, -4.476757e-21, 1.125836e-20, 
    4.436584e-20, -2.872517e-20, 3.161919e-20, 4.058902e-21, 2.354308e-21, 
    -2.194184e-20, -1.992375e-20, 9.059537e-21, -2.914726e-20, 8.057925e-22, 
    -1.219332e-20, -9.230579e-21, 1.662458e-20, 8.703589e-21, 3.242782e-20, 
    -2.925989e-21, 2.744693e-20, 9.265081e-21, -1.839165e-21, -7.058091e-21, 
    -3.471029e-20, -1.769614e-21, -2.349494e-20, -3.056871e-21, 4.984536e-21, 
    3.221661e-20, 1.441643e-20, -3.500801e-20, -2.822219e-21, 7.924935e-21, 
    2.279742e-20, 2.580738e-20, -6.421944e-21, 5.340795e-21, 2.222349e-20, 
    -1.49717e-20, 5.202076e-20, 3.516048e-21, 4.04531e-20, -3.91206e-20, 
    6.059288e-20, -1.527821e-20, -2.448745e-21, -5.146245e-21, -1.5188e-20, 
    2.129501e-20, -4.707014e-20, -2.854563e-20, -1.339918e-20, -1.559769e-20, 
    2.25359e-20, -3.733486e-20, -2.628286e-21, 3.927962e-21, -1.256286e-20, 
    -9.993385e-21, -1.379641e-20, 1.599039e-20, -1.394173e-20, 1.071975e-20, 
    1.755786e-20, -1.559994e-20, -3.38112e-20, 1.494373e-20, 1.522512e-21, 
    6.907949e-21, 2.01228e-20, 1.153006e-20, 8.188761e-24, 1.366713e-21, 
    1.950818e-21, -2.220282e-21, 4.244925e-21, 2.039817e-20, -2.747583e-21, 
    -1.04797e-20, -4.401015e-20, -3.692238e-20, -2.012872e-20, 6.280302e-21, 
    1.599776e-20, -1.348003e-20, 1.339775e-20 ;

 M_SOIL2C_TO_LEACHING =
  -1.250771e-20, -3.583301e-20, 8.624851e-23, -7.694792e-21, -2.547406e-20, 
    3.448178e-21, 1.133636e-20, -1.756491e-20, 2.310589e-20, -9.513056e-21, 
    -2.564199e-20, 5.935939e-21, -2.734091e-20, 1.175084e-20, 9.253497e-21, 
    -1.116362e-20, -2.169137e-20, -9.635597e-22, -9.123178e-21, 
    -1.419196e-20, -3.528197e-20, -6.172311e-21, -3.293445e-20, 
    -2.479547e-20, 7.105868e-21, -2.495378e-21, -2.395775e-20, -1.775182e-20, 
    3.028416e-20, -4.76232e-21, 1.702916e-20, 6.618728e-21, 1.267316e-20, 
    -9.411264e-21, 3.642165e-20, -6.38408e-22, -4.043322e-21, -1.223262e-20, 
    6.870933e-21, -4.487797e-21, 3.395004e-20, 2.19563e-20, 2.593404e-20, 
    3.198534e-20, 8.02756e-21, 1.390414e-20, -4.205084e-20, 3.070201e-20, 
    2.769574e-20, 8.155104e-21, -1.528783e-20, 4.994725e-21, 6.563586e-21, 
    -5.10411e-20, -2.231596e-20, 4.370752e-21, -2.69776e-20, -2.135947e-20, 
    -1.313933e-20, -9.122321e-21, 2.868983e-20, -2.141716e-20, -6.509588e-21, 
    1.45253e-20, 2.176009e-20, 1.18023e-20, -1.1007e-20, 1.636389e-20, 
    2.010385e-20, 2.546552e-21, -1.257615e-20, -6.549739e-21, 5.891516e-20, 
    -7.141488e-21, 1.311841e-20, -1.992544e-20, -2.418056e-20, 3.706799e-20, 
    -8.008921e-21, 3.333227e-20, 1.770159e-21, 4.950764e-22, -3.313181e-20, 
    -1.67012e-20, -1.771423e-20, 1.873855e-20, 4.931394e-21, -1.148567e-20, 
    2.857294e-21, -3.824189e-20, 3.562776e-20, 1.862913e-20, 5.499108e-21, 
    2.677433e-20, 3.16418e-20, -7.175991e-21, 1.635371e-20, 3.353178e-21, 
    -2.225571e-20, -9.017434e-21, -6.842667e-21, 1.913551e-20, 1.816836e-21, 
    -2.309091e-20, -1.958053e-20, -2.222518e-20, 2.868308e-21, 1.221142e-20, 
    -1.059703e-20, 3.25194e-20, 1.294255e-20, 1.697938e-20, -1.754176e-20, 
    -5.779594e-21, -1.654004e-20, -1.261206e-20, -1.913691e-20, 2.013269e-20, 
    -7.974419e-21, -3.545515e-22, -2.950152e-20, -6.257384e-21, 1.409187e-20, 
    -1.478428e-20, 1.068497e-20, 9.11071e-21, 2.483817e-20, -8.032101e-21, 
    4.411165e-21, 1.484393e-20, 1.291226e-21, -2.946619e-21, 8.018241e-22, 
    5.03402e-21, 3.732867e-21, -1.30305e-20, 2.226248e-20, -1.634917e-20, 
    2.328146e-20, 1.763384e-21, 7.944692e-22, 1.924322e-20, 1.419479e-20, 
    1.805377e-20, 8.24838e-21, 1.159564e-20, 2.486502e-20, -2.521903e-20, 
    9.67222e-21, 1.733394e-20, -7.937091e-21, 3.029161e-21, 3.125876e-21, 
    -1.13706e-20, -3.015886e-21, 3.034464e-20, 1.483628e-20, -2.361115e-20, 
    2.565526e-20, -2.309355e-21, -1.946093e-20, -8.3038e-21, -5.647542e-21, 
    5.718499e-21, 9.723115e-21, 1.07774e-20, -2.168715e-20, 8.640259e-21, 
    -2.212736e-20, -3.960689e-20, 2.257916e-20, -1.986743e-21, 3.919298e-20, 
    4.143164e-20, -1.665623e-20, 1.47885e-20, 4.617282e-21, -1.561267e-20, 
    -5.312512e-21, -3.112881e-22, 1.272062e-20, 1.880754e-20, -6.694189e-21, 
    -1.592935e-20, -2.297104e-20, -1.355552e-20, -1.375231e-20, 2.862195e-20, 
    -1.660677e-20, 2.624729e-20, -3.395455e-20, 6.563586e-21, 1.521431e-20, 
    -1.150657e-20, 4.236436e-20, 1.775522e-20, -2.699372e-20, 4.175e-20, 
    1.328437e-20, 9.508498e-21, -3.699927e-20, -3.71282e-20, 1.830144e-20, 
    -6.01425e-21, -6.321025e-21, 2.841558e-20, 4.228946e-20, 3.182505e-20, 
    -2.65851e-21, 2.643477e-20, -1.824746e-21, -5.572905e-21, -2.372083e-20, 
    -1.318768e-20, 3.06706e-21, -3.005796e-20, -2.436261e-20, 1.49768e-20, 
    -1.032842e-20, -4.175658e-21, -1.23262e-20, 4.734098e-20, -1.338729e-20, 
    2.27553e-20, 1.136518e-20, -4.231009e-20, 2.461227e-20, 1.081134e-20, 
    -3.631948e-21, 6.145159e-21, 5.715413e-21, -3.394179e-21, 5.087734e-21, 
    2.681137e-20, -8.401633e-21, 2.772736e-21, 1.447864e-20, -2.138377e-20, 
    -1.121224e-20, 1.824972e-20, 7.613368e-21, -4.702386e-21, 1.929271e-20, 
    -1.411365e-20, -6.804768e-21, -8.076482e-21, 1.513966e-20, 7.981174e-22, 
    8.629498e-21, -3.393023e-20, 2.272702e-20, -7.229704e-21, 2.581627e-21, 
    -1.346899e-20, -4.670554e-22, -1.960172e-20, -1.203613e-20, 
    -1.034794e-20, -1.134315e-20, 2.46202e-21, -4.053708e-20, -6.747096e-21, 
    -1.471729e-20, 5.490608e-21, 1.744053e-20, -1.283675e-22, -4.668456e-21, 
    -1.026314e-20, 1.959917e-20, -2.222178e-20, 2.549092e-21, 2.453311e-20, 
    -6.135237e-21, 1.862913e-20, 3.593196e-20, -2.874073e-20, -1.392648e-20, 
    -3.264891e-20, -1.337741e-20, -5.479023e-21, -6.0236e-21, 3.049025e-20, 
    3.350302e-22, 2.528715e-20, -7.832214e-21, 9.986626e-21, 5.718499e-21, 
    -2.40322e-21, 7.577747e-21, 2.106351e-21, -4.432948e-21, -3.452453e-20, 
    1.02586e-20, 1.882428e-21, -1.403759e-20, 7.528281e-21, 2.322549e-20, 
    1.57029e-21, 2.487468e-21, -9.101656e-21, -2.570558e-20, 1.387839e-20, 
    1.828931e-20, 1.532202e-20, -9.570712e-21, 1.478824e-20, -5.882486e-21, 
    2.216185e-20, -2.074139e-20, 3.608436e-20, 1.61982e-20, -5.589521e-22, 
    -2.85182e-20, -2.404053e-21, 1.779231e-21, 1.585158e-20, 7.608394e-22, 
    7.916353e-22, -3.71026e-21, 2.141402e-20, -8.536567e-23, 9.642803e-21, 
    -2.269028e-20, -1.185857e-20, 2.226561e-20, -1.979512e-20, -2.049401e-20, 
    -2.87359e-20, -3.26809e-21, 4.514656e-21, 3.629162e-20, 7.201732e-21, 
    9.993386e-21, -1.650017e-20, 1.52505e-20, 5.281666e-20, 7.52121e-21, 
    -1.618663e-20 ;

 M_SOIL3C_TO_LEACHING =
  -1.5216e-20, -5.559613e-21, -4.39208e-20, -1.570861e-21, 3.026687e-20, 
    1.814849e-20, -2.004702e-20, 9.435552e-21, -3.18327e-21, 3.6539e-20, 
    -2.224866e-20, 2.311323e-21, -5.230533e-22, 3.236412e-21, 3.107919e-20, 
    2.273045e-20, -2.785265e-20, 2.284917e-20, 6.147983e-21, 1.427142e-20, 
    1.379164e-21, 2.234457e-21, 1.578488e-20, -2.373157e-20, 1.914031e-20, 
    1.168046e-20, -2.177507e-20, 6.081003e-20, -1.407178e-20, -7.836745e-21, 
    -2.892049e-21, 2.506418e-21, 2.347373e-20, 2.793551e-20, 6.339475e-20, 
    -3.274164e-20, 3.527718e-20, -2.015675e-20, -3.068177e-21, -4.075e-21, 
    -2.525436e-20, -1.567489e-20, -5.7595e-21, 1.02658e-21, -2.900309e-20, 
    -4.914413e-21, -1.519366e-20, 1.046697e-20, -1.137286e-20, 1.877529e-20, 
    1.87097e-20, -9.287427e-21, -7.608282e-21, -7.451658e-21, -3.248692e-20, 
    -3.329607e-20, 1.895703e-21, -1.896265e-21, 8.275518e-21, -1.503648e-20, 
    -2.36097e-20, -2.885183e-20, 4.498247e-21, -2.132046e-20, 2.120365e-20, 
    -8.594188e-21, -4.349524e-21, -1.653128e-20, 1.604102e-20, 3.939797e-20, 
    1.415689e-20, -9.217304e-21, -3.596141e-20, -4.407151e-20, -3.488935e-22, 
    -3.735185e-20, 2.378584e-20, 1.195782e-20, -3.217478e-20, 5.806669e-20, 
    1.200843e-20, -4.149613e-20, 5.661599e-20, 2.321701e-20, 2.078186e-20, 
    -2.220679e-20, 8.440078e-21, 9.472878e-21, 4.531034e-21, -2.397161e-20, 
    -1.949486e-20, -1.300166e-20, 1.634721e-20, -4.278267e-21, 2.055171e-20, 
    1.959033e-21, -1.475317e-20, 1.779902e-20, -1.690647e-20, -2.11313e-20, 
    -5.603733e-21, 9.022772e-21, -3.770471e-20, 2.267134e-20, 4.239561e-21, 
    9.220128e-21, 6.351689e-20, 5.054916e-20, 1.77634e-20, -2.637201e-20, 
    -1.401761e-21, -9.401359e-21, -2.013552e-20, -2.322576e-20, 
    -3.475693e-20, 1.640602e-20, 5.974645e-21, 3.213602e-20, 1.861243e-20, 
    -6.235921e-21, 1.148594e-20, -2.507251e-21, 4.546762e-20, -2.584414e-20, 
    -6.56641e-21, 3.03534e-20, 4.160366e-21, 7.007906e-20, 2.62442e-20, 
    3.814885e-20, 5.899747e-21, 3.878527e-21, 4.191211e-21, -1.159961e-20, 
    -2.486165e-20, -4.15357e-20, 1.986551e-20, -1.933369e-20, -2.199365e-21, 
    -1.23248e-20, -8.739151e-22, -1.467925e-21, -6.295283e-21, 1.605966e-20, 
    -4.280969e-20, 1.844788e-20, 1.875182e-20, -2.613851e-21, 1.842698e-20, 
    1.798505e-20, 2.317375e-20, 1.761677e-21, -1.804529e-20, -3.216485e-20, 
    -2.509545e-20, 1.114328e-20, 2.654784e-20, -2.760857e-21, -8.717435e-21, 
    2.281524e-20, -6.70326e-21, 1.086111e-20, -1.093151e-20, -2.282495e-21, 
    2.008492e-20, -3.093063e-21, -2.863724e-20, 1.350917e-20, 4.465425e-21, 
    -3.816043e-23, -5.811246e-21, 1.21956e-20, -9.299012e-21, -8.639402e-21, 
    -2.559505e-20, -2.201201e-20, 2.222544e-21, -5.4072e-20, 2.078411e-20, 
    4.965041e-21, 9.591368e-21, 2.338748e-20, -1.518805e-21, 3.139755e-20, 
    1.500934e-20, -1.077317e-20, 1.196543e-20, -1.752083e-21, -2.336968e-20, 
    1.011696e-20, -3.898022e-21, -3.354855e-20, -2.468154e-20, -3.398255e-20, 
    4.602301e-21, 1.771674e-20, -3.498792e-20, -2.13179e-20, -2.833726e-20, 
    -1.456572e-20, 3.22993e-21, -2.532676e-20, -1.490868e-20, 5.12803e-20, 
    2.242367e-20, 9.004967e-21, 3.269386e-20, 1.941087e-20, -2.165434e-21, 
    6.268145e-21, 2.852727e-20, 1.404661e-20, -9.166414e-21, -9.490138e-21, 
    -3.258472e-20, 2.464395e-20, -2.074567e-20, 3.180608e-20, 2.809638e-20, 
    2.98869e-20, 2.464875e-20, -2.791008e-20, 3.180408e-20, 6.844959e-22, 
    4.408341e-21, -1.509671e-20, 4.940381e-20, -5.703534e-21, -1.07206e-20, 
    -4.742253e-21, -1.427479e-20, -1.04503e-20, -4.287584e-20, 3.175151e-20, 
    2.246748e-20, -3.532736e-21, 1.100812e-20, 2.020961e-20, -1.123035e-20, 
    -3.401544e-21, -1.863167e-22, -1.079239e-20, 4.433138e-22, -3.902616e-20, 
    4.96278e-21, -2.361706e-20, 1.716686e-20, 1.286396e-20, 1.253542e-20, 
    1.888924e-20, -3.236619e-20, -2.164502e-20, -1.956355e-20, -1.74032e-20, 
    -1.638057e-20, 2.246976e-20, -6.790905e-21, 1.171099e-20, -3.115976e-20, 
    1.155183e-20, 2.302474e-20, -7.100503e-21, 2.237786e-20, -1.816037e-20, 
    5.49165e-20, 2.35676e-20, -4.165613e-20, 3.372666e-20, -4.779253e-20, 
    -1.630962e-20, -1.6647e-21, 3.966407e-21, -1.18761e-20, -4.822255e-21, 
    -8.736663e-21, 4.61671e-21, -1.465082e-20, 2.116495e-20, -5.856199e-21, 
    -1.953048e-20, -1.983468e-20, -2.238577e-20, -3.931031e-20, 
    -1.628616e-20, -3.832302e-20, -1.813294e-20, 2.242628e-21, -1.575037e-20, 
    2.010498e-20, 1.492903e-20, -3.331672e-20, -3.061973e-21, 1.624063e-20, 
    2.692162e-21, 4.118568e-20, 6.618156e-21, -2.268098e-20, 1.929694e-20, 
    1.799887e-21, -4.682319e-21, -2.778536e-20, 9.986054e-21, 1.444528e-20, 
    4.814066e-21, 2.866879e-21, 6.044446e-20, -5.139453e-21, 4.420219e-21, 
    1.753072e-20, -2.666135e-22, 1.729492e-20, -8.208246e-21, 1.556941e-20, 
    -6.184747e-21, -1.276106e-20, -8.895549e-21, -2.502225e-20, 3.675388e-20, 
    2.307309e-20, 1.613009e-20, 1.387616e-20, -2.931549e-20, 1.60543e-20, 
    -3.814885e-21, 3.291835e-20, 1.216789e-20, 2.758095e-20, -2.980406e-20, 
    2.643137e-20, -1.044679e-21, -1.455785e-21, -2.384438e-20, -4.90171e-21, 
    1.117747e-20, -2.170798e-21, -1.823611e-21, -1.441557e-20, -4.59523e-21 ;

 NBP =
  -6.358388e-08, -6.386347e-08, -6.380911e-08, -6.403462e-08, -6.390952e-08, 
    -6.405718e-08, -6.364056e-08, -6.387457e-08, -6.372518e-08, 
    -6.360905e-08, -6.447225e-08, -6.404468e-08, -6.491634e-08, 
    -6.464366e-08, -6.532863e-08, -6.487392e-08, -6.542031e-08, -6.53155e-08, 
    -6.563094e-08, -6.554057e-08, -6.594404e-08, -6.567264e-08, 
    -6.615318e-08, -6.587923e-08, -6.592209e-08, -6.566369e-08, 
    -6.413072e-08, -6.441902e-08, -6.411364e-08, -6.415475e-08, -6.41363e-08, 
    -6.391211e-08, -6.379913e-08, -6.356251e-08, -6.360547e-08, 
    -6.377926e-08, -6.417324e-08, -6.403949e-08, -6.437654e-08, 
    -6.436893e-08, -6.474416e-08, -6.457498e-08, -6.520563e-08, 
    -6.502638e-08, -6.554434e-08, -6.541408e-08, -6.553822e-08, 
    -6.550058e-08, -6.553871e-08, -6.534768e-08, -6.542952e-08, 
    -6.526142e-08, -6.460666e-08, -6.47991e-08, -6.422516e-08, -6.388007e-08, 
    -6.365083e-08, -6.348817e-08, -6.351116e-08, -6.3555e-08, -6.378028e-08, 
    -6.399208e-08, -6.415348e-08, -6.426145e-08, -6.436783e-08, 
    -6.468986e-08, -6.486028e-08, -6.524188e-08, -6.5173e-08, -6.528968e-08, 
    -6.540112e-08, -6.558825e-08, -6.555744e-08, -6.563989e-08, 
    -6.528659e-08, -6.55214e-08, -6.513378e-08, -6.52398e-08, -6.439678e-08, 
    -6.407557e-08, -6.393907e-08, -6.381956e-08, -6.352884e-08, 
    -6.372961e-08, -6.365047e-08, -6.383875e-08, -6.395839e-08, 
    -6.389921e-08, -6.426441e-08, -6.412242e-08, -6.487038e-08, 
    -6.454822e-08, -6.538812e-08, -6.518714e-08, -6.54363e-08, -6.530916e-08, 
    -6.5527e-08, -6.533094e-08, -6.567057e-08, -6.574452e-08, -6.569399e-08, 
    -6.588811e-08, -6.532007e-08, -6.553822e-08, -6.389756e-08, 
    -6.390721e-08, -6.395216e-08, -6.375454e-08, -6.374245e-08, 
    -6.356133e-08, -6.372249e-08, -6.379111e-08, -6.396532e-08, 
    -6.406837e-08, -6.416632e-08, -6.438169e-08, -6.462222e-08, 
    -6.495855e-08, -6.520017e-08, -6.536213e-08, -6.526282e-08, -6.53505e-08, 
    -6.525248e-08, -6.520654e-08, -6.571682e-08, -6.543029e-08, 
    -6.586019e-08, -6.58364e-08, -6.564185e-08, -6.583908e-08, -6.391399e-08, 
    -6.385844e-08, -6.366564e-08, -6.381653e-08, -6.354161e-08, -6.36955e-08, 
    -6.378399e-08, -6.41254e-08, -6.420041e-08, -6.426996e-08, -6.440733e-08, 
    -6.458363e-08, -6.489289e-08, -6.516198e-08, -6.54076e-08, -6.538961e-08, 
    -6.539594e-08, -6.545082e-08, -6.531489e-08, -6.547314e-08, -6.54997e-08, 
    -6.543026e-08, -6.583321e-08, -6.571809e-08, -6.58359e-08, -6.576094e-08, 
    -6.38765e-08, -6.396994e-08, -6.391945e-08, -6.40144e-08, -6.394751e-08, 
    -6.424496e-08, -6.433414e-08, -6.475143e-08, -6.458016e-08, 
    -6.485271e-08, -6.460785e-08, -6.465124e-08, -6.486162e-08, 
    -6.462108e-08, -6.514714e-08, -6.47905e-08, -6.545295e-08, -6.509682e-08, 
    -6.547527e-08, -6.540655e-08, -6.552033e-08, -6.562224e-08, 
    -6.575045e-08, -6.598701e-08, -6.593223e-08, -6.613006e-08, 
    -6.410925e-08, -6.423046e-08, -6.421978e-08, -6.434662e-08, 
    -6.444042e-08, -6.464373e-08, -6.496981e-08, -6.484719e-08, 
    -6.507229e-08, -6.511748e-08, -6.477549e-08, -6.498548e-08, 
    -6.431157e-08, -6.442045e-08, -6.435562e-08, -6.411882e-08, 
    -6.487545e-08, -6.448715e-08, -6.520416e-08, -6.499381e-08, 
    -6.560771e-08, -6.530242e-08, -6.590207e-08, -6.615844e-08, 
    -6.639969e-08, -6.668164e-08, -6.42966e-08, -6.421424e-08, -6.43617e-08, 
    -6.456572e-08, -6.4755e-08, -6.500665e-08, -6.503239e-08, -6.507953e-08, 
    -6.520164e-08, -6.530431e-08, -6.509445e-08, -6.533005e-08, 
    -6.444572e-08, -6.490915e-08, -6.418311e-08, -6.440175e-08, 
    -6.455369e-08, -6.448703e-08, -6.483317e-08, -6.491475e-08, 
    -6.524627e-08, -6.507489e-08, -6.609517e-08, -6.564377e-08, 
    -6.689631e-08, -6.654629e-08, -6.418547e-08, -6.429631e-08, 
    -6.468208e-08, -6.449854e-08, -6.502344e-08, -6.515264e-08, 
    -6.525767e-08, -6.539194e-08, -6.540643e-08, -6.548598e-08, 
    -6.535562e-08, -6.548083e-08, -6.500718e-08, -6.521884e-08, 
    -6.463799e-08, -6.477936e-08, -6.471433e-08, -6.464298e-08, 
    -6.486317e-08, -6.509775e-08, -6.510275e-08, -6.517797e-08, 
    -6.538995e-08, -6.502557e-08, -6.615345e-08, -6.545692e-08, 
    -6.441718e-08, -6.463069e-08, -6.466117e-08, -6.457847e-08, 
    -6.513969e-08, -6.493634e-08, -6.548404e-08, -6.533602e-08, 
    -6.557855e-08, -6.545803e-08, -6.54403e-08, -6.528551e-08, -6.518914e-08, 
    -6.494567e-08, -6.474756e-08, -6.459047e-08, -6.4627e-08, -6.479956e-08, 
    -6.51121e-08, -6.540775e-08, -6.534299e-08, -6.556012e-08, -6.498538e-08, 
    -6.522639e-08, -6.513324e-08, -6.537611e-08, -6.484393e-08, 
    -6.529714e-08, -6.472809e-08, -6.477798e-08, -6.493231e-08, 
    -6.524274e-08, -6.53114e-08, -6.538474e-08, -6.533948e-08, -6.512003e-08, 
    -6.508407e-08, -6.492856e-08, -6.488562e-08, -6.476711e-08, 
    -6.466901e-08, -6.475865e-08, -6.485278e-08, -6.512012e-08, 
    -6.536104e-08, -6.562369e-08, -6.568797e-08, -6.599488e-08, 
    -6.574506e-08, -6.615733e-08, -6.580684e-08, -6.641355e-08, 
    -6.532339e-08, -6.579651e-08, -6.493933e-08, -6.503167e-08, 
    -6.519871e-08, -6.558179e-08, -6.537497e-08, -6.561685e-08, 
    -6.508266e-08, -6.480552e-08, -6.47338e-08, -6.460002e-08, -6.473686e-08, 
    -6.472573e-08, -6.485668e-08, -6.48146e-08, -6.512899e-08, -6.496011e-08, 
    -6.543986e-08, -6.561493e-08, -6.610933e-08, -6.641241e-08, 
    -6.672092e-08, -6.685712e-08, -6.689857e-08, -6.69159e-08 ;

 NDEPLOY =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NDEP_TO_SMINN =
  3.989144e-10, 3.989147e-10, 3.989121e-10, 3.989123e-10, 3.989108e-10, 
    3.989089e-10, 3.989084e-10, 3.989066e-10, 3.98906e-10, 3.989042e-10, 
    3.989026e-10, 3.989029e-10, 3.989014e-10, 3.988995e-10, 3.988979e-10, 
    3.988982e-10, 3.988966e-10, 3.988948e-10, 3.988943e-10, 3.988924e-10, 
    3.988909e-10, 3.988911e-10, 3.988885e-10, 3.988888e-10, 3.988872e-10, 
    3.988854e-10, 3.989112e-10, 3.989115e-10, 3.989089e-10, 3.989092e-10, 
    3.989076e-10, 3.989057e-10, 3.989052e-10, 3.989034e-10, 3.989018e-10, 
    3.989021e-10, 3.989005e-10, 3.988987e-10, 3.988971e-10, 3.988974e-10, 
    3.988947e-10, 3.98895e-10, 3.988934e-10, 3.988916e-10, 3.988911e-10, 
    3.988892e-10, 3.988887e-10, 3.988869e-10, 3.988853e-10, 3.988856e-10, 
    3.98883e-10, 3.988832e-10, 3.989091e-10, 3.989072e-10, 3.989067e-10, 
    3.989049e-10, 3.989033e-10, 3.989036e-10, 3.98901e-10, 3.989012e-10, 
    3.988997e-10, 3.988978e-10, 3.988973e-10, 3.988955e-10, 3.988939e-10, 
    3.988942e-10, 3.988926e-10, 3.988908e-10, 3.988903e-10, 3.988884e-10, 
    3.988879e-10, 3.98886e-10, 3.988855e-10, 3.988837e-10, 3.988821e-10, 
    3.988824e-10, 3.988798e-10, 3.9888e-10, 3.989059e-10, 3.98904e-10, 
    3.989035e-10, 3.989017e-10, 3.989001e-10, 3.989004e-10, 3.988988e-10, 
    3.98897e-10, 3.988965e-10, 3.988946e-10, 3.988941e-10, 3.988923e-10, 
    3.988907e-10, 3.98891e-10, 3.988894e-10, 3.988876e-10, 3.98886e-10, 
    3.988863e-10, 3.988836e-10, 3.988839e-10, 3.988813e-10, 3.988816e-10, 
    3.988789e-10, 3.988792e-10, 3.988766e-10, 3.988768e-10, 3.989017e-10, 
    3.989019e-10, 3.989004e-10, 3.988985e-10, 3.98898e-10, 3.988962e-10, 
    3.988946e-10, 3.988949e-10, 3.988933e-10, 3.988914e-10, 3.988899e-10, 
    3.988901e-10, 3.988886e-10, 3.988867e-10, 3.988862e-10, 3.988844e-10, 
    3.988839e-10, 3.98882e-10, 3.988815e-10, 3.988797e-10, 3.988781e-10, 
    3.988784e-10, 3.988757e-10, 3.98876e-10, 3.988744e-10, 3.988726e-10, 
    3.988995e-10, 3.988977e-10, 3.988972e-10, 3.988953e-10, 3.988938e-10, 
    3.98894e-10, 3.988924e-10, 3.988906e-10, 3.98889e-10, 3.988893e-10, 
    3.988878e-10, 3.988859e-10, 3.988854e-10, 3.988835e-10, 3.98883e-10, 
    3.988812e-10, 3.988807e-10, 3.988788e-10, 3.988783e-10, 3.988765e-10, 
    3.988749e-10, 3.988752e-10, 3.988725e-10, 3.988728e-10, 3.988712e-10, 
    3.988694e-10, 3.988963e-10, 3.988945e-10, 3.988929e-10, 3.988932e-10, 
    3.988906e-10, 3.988908e-10, 3.988893e-10, 3.988874e-10, 3.988858e-10, 
    3.988861e-10, 3.988835e-10, 3.988838e-10, 3.988822e-10, 3.988803e-10, 
    3.988798e-10, 3.98878e-10, 3.988775e-10, 3.988756e-10, 3.988751e-10, 
    3.988733e-10, 3.988717e-10, 3.98872e-10, 3.988694e-10, 3.988696e-10, 
    3.98867e-10, 3.988673e-10, 3.988931e-10, 3.988913e-10, 3.988908e-10, 
    3.988889e-10, 3.988874e-10, 3.988876e-10, 3.988861e-10, 3.988842e-10, 
    3.988826e-10, 3.988829e-10, 3.988803e-10, 3.988806e-10, 3.98879e-10, 
    3.988772e-10, 3.988767e-10, 3.988748e-10, 3.988743e-10, 3.988724e-10, 
    3.988719e-10, 3.988701e-10, 3.988685e-10, 3.988688e-10, 3.988662e-10, 
    3.988664e-10, 3.988649e-10, 3.98863e-10, 3.988899e-10, 3.988881e-10, 
    3.988865e-10, 3.988868e-10, 3.988842e-10, 3.988845e-10, 3.988829e-10, 
    3.98881e-10, 3.988795e-10, 3.988797e-10, 3.988782e-10, 3.988763e-10, 
    3.988758e-10, 3.98874e-10, 3.988724e-10, 3.988727e-10, 3.9887e-10, 
    3.988703e-10, 3.988687e-10, 3.988669e-10, 3.988653e-10, 3.988656e-10, 
    3.98863e-10, 3.988632e-10, 3.988606e-10, 3.988609e-10, 3.988868e-10, 
    3.988849e-10, 3.988833e-10, 3.988836e-10, 3.98881e-10, 3.988813e-10, 
    3.988786e-10, 3.988789e-10, 3.988763e-10, 3.988765e-10, 3.988739e-10, 
    3.988742e-10, 3.988716e-10, 3.988719e-10, 3.988703e-10, 3.988684e-10, 
    3.988679e-10, 3.988661e-10, 3.988645e-10, 3.988648e-10, 3.988632e-10, 
    3.988614e-10, 3.988609e-10, 3.98859e-10, 3.988585e-10, 3.988566e-10, 
    3.988836e-10, 3.988817e-10, 3.988802e-10, 3.988804e-10, 3.988778e-10, 
    3.988781e-10, 3.988765e-10, 3.988747e-10, 3.988731e-10, 3.988734e-10, 
    3.988707e-10, 3.98871e-10, 3.988684e-10, 3.988687e-10, 3.98866e-10, 
    3.988663e-10, 3.988637e-10, 3.988639e-10, 3.988613e-10, 3.988616e-10, 
    3.9886e-10, 3.988582e-10, 3.988566e-10, 3.988569e-10, 3.988542e-10, 
    3.988545e-10, 3.988793e-10, 3.988796e-10, 3.98878e-10, 3.988762e-10, 
    3.988746e-10, 3.988749e-10, 3.988722e-10, 3.988725e-10, 3.988699e-10, 
    3.988702e-10, 3.988686e-10, 3.988667e-10, 3.988652e-10, 3.988655e-10, 
    3.988628e-10, 3.988631e-10, 3.988605e-10, 3.988607e-10, 3.988592e-10, 
    3.988573e-10, 3.988568e-10, 3.98855e-10, 3.988545e-10, 3.988526e-10, 
    3.988521e-10, 3.988503e-10, 3.988761e-10, 3.988764e-10, 3.988748e-10, 
    3.98873e-10, 3.988725e-10, 3.988706e-10, 3.98869e-10, 3.988693e-10, 
    3.988678e-10, 3.988659e-10, 3.988644e-10, 3.988646e-10, 3.98862e-10, 
    3.988623e-10, 3.988607e-10, 3.988589e-10, 3.988573e-10, 3.988576e-10, 
    3.988549e-10, 3.988552e-10, 3.988536e-10, 3.988518e-10, 3.988513e-10, 
    3.988494e-10, 3.988489e-10, 3.988476e-10 ;

 NEE =
  6.358388e-08, 6.386347e-08, 6.380911e-08, 6.403462e-08, 6.390952e-08, 
    6.405718e-08, 6.364056e-08, 6.387457e-08, 6.372518e-08, 6.360905e-08, 
    6.447225e-08, 6.404468e-08, 6.491634e-08, 6.464366e-08, 6.532863e-08, 
    6.487392e-08, 6.542031e-08, 6.53155e-08, 6.563094e-08, 6.554057e-08, 
    6.594404e-08, 6.567264e-08, 6.615318e-08, 6.587923e-08, 6.592209e-08, 
    6.566369e-08, 6.413072e-08, 6.441902e-08, 6.411364e-08, 6.415475e-08, 
    6.41363e-08, 6.391211e-08, 6.379913e-08, 6.356251e-08, 6.360547e-08, 
    6.377926e-08, 6.417324e-08, 6.403949e-08, 6.437654e-08, 6.436893e-08, 
    6.474416e-08, 6.457498e-08, 6.520563e-08, 6.502638e-08, 6.554434e-08, 
    6.541408e-08, 6.553822e-08, 6.550058e-08, 6.553871e-08, 6.534768e-08, 
    6.542952e-08, 6.526142e-08, 6.460666e-08, 6.47991e-08, 6.422516e-08, 
    6.388007e-08, 6.365083e-08, 6.348817e-08, 6.351116e-08, 6.3555e-08, 
    6.378028e-08, 6.399208e-08, 6.415348e-08, 6.426145e-08, 6.436783e-08, 
    6.468986e-08, 6.486028e-08, 6.524188e-08, 6.5173e-08, 6.528968e-08, 
    6.540112e-08, 6.558825e-08, 6.555744e-08, 6.563989e-08, 6.528659e-08, 
    6.55214e-08, 6.513378e-08, 6.52398e-08, 6.439678e-08, 6.407557e-08, 
    6.393907e-08, 6.381956e-08, 6.352884e-08, 6.372961e-08, 6.365047e-08, 
    6.383875e-08, 6.395839e-08, 6.389921e-08, 6.426441e-08, 6.412242e-08, 
    6.487038e-08, 6.454822e-08, 6.538812e-08, 6.518714e-08, 6.54363e-08, 
    6.530916e-08, 6.5527e-08, 6.533094e-08, 6.567057e-08, 6.574452e-08, 
    6.569399e-08, 6.588811e-08, 6.532007e-08, 6.553822e-08, 6.389756e-08, 
    6.390721e-08, 6.395216e-08, 6.375454e-08, 6.374245e-08, 6.356133e-08, 
    6.372249e-08, 6.379111e-08, 6.396532e-08, 6.406837e-08, 6.416632e-08, 
    6.438169e-08, 6.462222e-08, 6.495855e-08, 6.520017e-08, 6.536213e-08, 
    6.526282e-08, 6.53505e-08, 6.525248e-08, 6.520654e-08, 6.571682e-08, 
    6.543029e-08, 6.586019e-08, 6.58364e-08, 6.564185e-08, 6.583908e-08, 
    6.391399e-08, 6.385844e-08, 6.366564e-08, 6.381653e-08, 6.354161e-08, 
    6.36955e-08, 6.378399e-08, 6.41254e-08, 6.420041e-08, 6.426996e-08, 
    6.440733e-08, 6.458363e-08, 6.489289e-08, 6.516198e-08, 6.54076e-08, 
    6.538961e-08, 6.539594e-08, 6.545082e-08, 6.531489e-08, 6.547314e-08, 
    6.54997e-08, 6.543026e-08, 6.583321e-08, 6.571809e-08, 6.58359e-08, 
    6.576094e-08, 6.38765e-08, 6.396994e-08, 6.391945e-08, 6.40144e-08, 
    6.394751e-08, 6.424496e-08, 6.433414e-08, 6.475143e-08, 6.458016e-08, 
    6.485271e-08, 6.460785e-08, 6.465124e-08, 6.486162e-08, 6.462108e-08, 
    6.514714e-08, 6.47905e-08, 6.545295e-08, 6.509682e-08, 6.547527e-08, 
    6.540655e-08, 6.552033e-08, 6.562224e-08, 6.575045e-08, 6.598701e-08, 
    6.593223e-08, 6.613006e-08, 6.410925e-08, 6.423046e-08, 6.421978e-08, 
    6.434662e-08, 6.444042e-08, 6.464373e-08, 6.496981e-08, 6.484719e-08, 
    6.507229e-08, 6.511748e-08, 6.477549e-08, 6.498548e-08, 6.431157e-08, 
    6.442045e-08, 6.435562e-08, 6.411882e-08, 6.487545e-08, 6.448715e-08, 
    6.520416e-08, 6.499381e-08, 6.560771e-08, 6.530242e-08, 6.590207e-08, 
    6.615844e-08, 6.639969e-08, 6.668164e-08, 6.42966e-08, 6.421424e-08, 
    6.43617e-08, 6.456572e-08, 6.4755e-08, 6.500665e-08, 6.503239e-08, 
    6.507953e-08, 6.520164e-08, 6.530431e-08, 6.509445e-08, 6.533005e-08, 
    6.444572e-08, 6.490915e-08, 6.418311e-08, 6.440175e-08, 6.455369e-08, 
    6.448703e-08, 6.483317e-08, 6.491475e-08, 6.524627e-08, 6.507489e-08, 
    6.609517e-08, 6.564377e-08, 6.689631e-08, 6.654629e-08, 6.418547e-08, 
    6.429631e-08, 6.468208e-08, 6.449854e-08, 6.502344e-08, 6.515264e-08, 
    6.525767e-08, 6.539194e-08, 6.540643e-08, 6.548598e-08, 6.535562e-08, 
    6.548083e-08, 6.500718e-08, 6.521884e-08, 6.463799e-08, 6.477936e-08, 
    6.471433e-08, 6.464298e-08, 6.486317e-08, 6.509775e-08, 6.510275e-08, 
    6.517797e-08, 6.538995e-08, 6.502557e-08, 6.615345e-08, 6.545692e-08, 
    6.441718e-08, 6.463069e-08, 6.466117e-08, 6.457847e-08, 6.513969e-08, 
    6.493634e-08, 6.548404e-08, 6.533602e-08, 6.557855e-08, 6.545803e-08, 
    6.54403e-08, 6.528551e-08, 6.518914e-08, 6.494567e-08, 6.474756e-08, 
    6.459047e-08, 6.4627e-08, 6.479956e-08, 6.51121e-08, 6.540775e-08, 
    6.534299e-08, 6.556012e-08, 6.498538e-08, 6.522639e-08, 6.513324e-08, 
    6.537611e-08, 6.484393e-08, 6.529714e-08, 6.472809e-08, 6.477798e-08, 
    6.493231e-08, 6.524274e-08, 6.53114e-08, 6.538474e-08, 6.533948e-08, 
    6.512003e-08, 6.508407e-08, 6.492856e-08, 6.488562e-08, 6.476711e-08, 
    6.466901e-08, 6.475865e-08, 6.485278e-08, 6.512012e-08, 6.536104e-08, 
    6.562369e-08, 6.568797e-08, 6.599488e-08, 6.574506e-08, 6.615733e-08, 
    6.580684e-08, 6.641355e-08, 6.532339e-08, 6.579651e-08, 6.493933e-08, 
    6.503167e-08, 6.519871e-08, 6.558179e-08, 6.537497e-08, 6.561685e-08, 
    6.508266e-08, 6.480552e-08, 6.47338e-08, 6.460002e-08, 6.473686e-08, 
    6.472573e-08, 6.485668e-08, 6.48146e-08, 6.512899e-08, 6.496011e-08, 
    6.543986e-08, 6.561493e-08, 6.610933e-08, 6.641241e-08, 6.672092e-08, 
    6.685712e-08, 6.689857e-08, 6.69159e-08 ;

 NEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NEP =
  -6.358388e-08, -6.386347e-08, -6.380911e-08, -6.403462e-08, -6.390952e-08, 
    -6.405718e-08, -6.364056e-08, -6.387457e-08, -6.372518e-08, 
    -6.360905e-08, -6.447225e-08, -6.404468e-08, -6.491634e-08, 
    -6.464366e-08, -6.532863e-08, -6.487392e-08, -6.542031e-08, -6.53155e-08, 
    -6.563094e-08, -6.554057e-08, -6.594404e-08, -6.567264e-08, 
    -6.615318e-08, -6.587923e-08, -6.592209e-08, -6.566369e-08, 
    -6.413072e-08, -6.441902e-08, -6.411364e-08, -6.415475e-08, -6.41363e-08, 
    -6.391211e-08, -6.379913e-08, -6.356251e-08, -6.360547e-08, 
    -6.377926e-08, -6.417324e-08, -6.403949e-08, -6.437654e-08, 
    -6.436893e-08, -6.474416e-08, -6.457498e-08, -6.520563e-08, 
    -6.502638e-08, -6.554434e-08, -6.541408e-08, -6.553822e-08, 
    -6.550058e-08, -6.553871e-08, -6.534768e-08, -6.542952e-08, 
    -6.526142e-08, -6.460666e-08, -6.47991e-08, -6.422516e-08, -6.388007e-08, 
    -6.365083e-08, -6.348817e-08, -6.351116e-08, -6.3555e-08, -6.378028e-08, 
    -6.399208e-08, -6.415348e-08, -6.426145e-08, -6.436783e-08, 
    -6.468986e-08, -6.486028e-08, -6.524188e-08, -6.5173e-08, -6.528968e-08, 
    -6.540112e-08, -6.558825e-08, -6.555744e-08, -6.563989e-08, 
    -6.528659e-08, -6.55214e-08, -6.513378e-08, -6.52398e-08, -6.439678e-08, 
    -6.407557e-08, -6.393907e-08, -6.381956e-08, -6.352884e-08, 
    -6.372961e-08, -6.365047e-08, -6.383875e-08, -6.395839e-08, 
    -6.389921e-08, -6.426441e-08, -6.412242e-08, -6.487038e-08, 
    -6.454822e-08, -6.538812e-08, -6.518714e-08, -6.54363e-08, -6.530916e-08, 
    -6.5527e-08, -6.533094e-08, -6.567057e-08, -6.574452e-08, -6.569399e-08, 
    -6.588811e-08, -6.532007e-08, -6.553822e-08, -6.389756e-08, 
    -6.390721e-08, -6.395216e-08, -6.375454e-08, -6.374245e-08, 
    -6.356133e-08, -6.372249e-08, -6.379111e-08, -6.396532e-08, 
    -6.406837e-08, -6.416632e-08, -6.438169e-08, -6.462222e-08, 
    -6.495855e-08, -6.520017e-08, -6.536213e-08, -6.526282e-08, -6.53505e-08, 
    -6.525248e-08, -6.520654e-08, -6.571682e-08, -6.543029e-08, 
    -6.586019e-08, -6.58364e-08, -6.564185e-08, -6.583908e-08, -6.391399e-08, 
    -6.385844e-08, -6.366564e-08, -6.381653e-08, -6.354161e-08, -6.36955e-08, 
    -6.378399e-08, -6.41254e-08, -6.420041e-08, -6.426996e-08, -6.440733e-08, 
    -6.458363e-08, -6.489289e-08, -6.516198e-08, -6.54076e-08, -6.538961e-08, 
    -6.539594e-08, -6.545082e-08, -6.531489e-08, -6.547314e-08, -6.54997e-08, 
    -6.543026e-08, -6.583321e-08, -6.571809e-08, -6.58359e-08, -6.576094e-08, 
    -6.38765e-08, -6.396994e-08, -6.391945e-08, -6.40144e-08, -6.394751e-08, 
    -6.424496e-08, -6.433414e-08, -6.475143e-08, -6.458016e-08, 
    -6.485271e-08, -6.460785e-08, -6.465124e-08, -6.486162e-08, 
    -6.462108e-08, -6.514714e-08, -6.47905e-08, -6.545295e-08, -6.509682e-08, 
    -6.547527e-08, -6.540655e-08, -6.552033e-08, -6.562224e-08, 
    -6.575045e-08, -6.598701e-08, -6.593223e-08, -6.613006e-08, 
    -6.410925e-08, -6.423046e-08, -6.421978e-08, -6.434662e-08, 
    -6.444042e-08, -6.464373e-08, -6.496981e-08, -6.484719e-08, 
    -6.507229e-08, -6.511748e-08, -6.477549e-08, -6.498548e-08, 
    -6.431157e-08, -6.442045e-08, -6.435562e-08, -6.411882e-08, 
    -6.487545e-08, -6.448715e-08, -6.520416e-08, -6.499381e-08, 
    -6.560771e-08, -6.530242e-08, -6.590207e-08, -6.615844e-08, 
    -6.639969e-08, -6.668164e-08, -6.42966e-08, -6.421424e-08, -6.43617e-08, 
    -6.456572e-08, -6.4755e-08, -6.500665e-08, -6.503239e-08, -6.507953e-08, 
    -6.520164e-08, -6.530431e-08, -6.509445e-08, -6.533005e-08, 
    -6.444572e-08, -6.490915e-08, -6.418311e-08, -6.440175e-08, 
    -6.455369e-08, -6.448703e-08, -6.483317e-08, -6.491475e-08, 
    -6.524627e-08, -6.507489e-08, -6.609517e-08, -6.564377e-08, 
    -6.689631e-08, -6.654629e-08, -6.418547e-08, -6.429631e-08, 
    -6.468208e-08, -6.449854e-08, -6.502344e-08, -6.515264e-08, 
    -6.525767e-08, -6.539194e-08, -6.540643e-08, -6.548598e-08, 
    -6.535562e-08, -6.548083e-08, -6.500718e-08, -6.521884e-08, 
    -6.463799e-08, -6.477936e-08, -6.471433e-08, -6.464298e-08, 
    -6.486317e-08, -6.509775e-08, -6.510275e-08, -6.517797e-08, 
    -6.538995e-08, -6.502557e-08, -6.615345e-08, -6.545692e-08, 
    -6.441718e-08, -6.463069e-08, -6.466117e-08, -6.457847e-08, 
    -6.513969e-08, -6.493634e-08, -6.548404e-08, -6.533602e-08, 
    -6.557855e-08, -6.545803e-08, -6.54403e-08, -6.528551e-08, -6.518914e-08, 
    -6.494567e-08, -6.474756e-08, -6.459047e-08, -6.4627e-08, -6.479956e-08, 
    -6.51121e-08, -6.540775e-08, -6.534299e-08, -6.556012e-08, -6.498538e-08, 
    -6.522639e-08, -6.513324e-08, -6.537611e-08, -6.484393e-08, 
    -6.529714e-08, -6.472809e-08, -6.477798e-08, -6.493231e-08, 
    -6.524274e-08, -6.53114e-08, -6.538474e-08, -6.533948e-08, -6.512003e-08, 
    -6.508407e-08, -6.492856e-08, -6.488562e-08, -6.476711e-08, 
    -6.466901e-08, -6.475865e-08, -6.485278e-08, -6.512012e-08, 
    -6.536104e-08, -6.562369e-08, -6.568797e-08, -6.599488e-08, 
    -6.574506e-08, -6.615733e-08, -6.580684e-08, -6.641355e-08, 
    -6.532339e-08, -6.579651e-08, -6.493933e-08, -6.503167e-08, 
    -6.519871e-08, -6.558179e-08, -6.537497e-08, -6.561685e-08, 
    -6.508266e-08, -6.480552e-08, -6.47338e-08, -6.460002e-08, -6.473686e-08, 
    -6.472573e-08, -6.485668e-08, -6.48146e-08, -6.512899e-08, -6.496011e-08, 
    -6.543986e-08, -6.561493e-08, -6.610933e-08, -6.641241e-08, 
    -6.672092e-08, -6.685712e-08, -6.689857e-08, -6.69159e-08 ;

 NET_NMIN =
  8.957549e-09, 8.996934e-09, 8.989277e-09, 9.021043e-09, 9.003422e-09, 
    9.024222e-09, 8.965534e-09, 8.998498e-09, 8.977454e-09, 8.961094e-09, 
    9.082692e-09, 9.022461e-09, 9.14525e-09, 9.106839e-09, 9.203327e-09, 
    9.139273e-09, 9.216242e-09, 9.201478e-09, 9.245912e-09, 9.233182e-09, 
    9.290019e-09, 9.251787e-09, 9.319479e-09, 9.280888e-09, 9.286926e-09, 
    9.250527e-09, 9.034581e-09, 9.075193e-09, 9.032175e-09, 9.037966e-09, 
    9.035367e-09, 9.003786e-09, 8.987872e-09, 8.954538e-09, 8.96059e-09, 
    8.985072e-09, 9.04057e-09, 9.02173e-09, 9.069208e-09, 9.068136e-09, 
    9.120994e-09, 9.097162e-09, 9.186e-09, 9.160751e-09, 9.233714e-09, 
    9.215364e-09, 9.232852e-09, 9.227549e-09, 9.232921e-09, 9.20601e-09, 
    9.217541e-09, 9.19386e-09, 9.101626e-09, 9.128733e-09, 9.047885e-09, 
    8.999272e-09, 8.96698e-09, 8.944066e-09, 8.947305e-09, 8.953481e-09, 
    8.985215e-09, 9.015051e-09, 9.037787e-09, 9.052997e-09, 9.067983e-09, 
    9.113346e-09, 9.137352e-09, 9.191107e-09, 9.181405e-09, 9.19784e-09, 
    9.213539e-09, 9.239899e-09, 9.23556e-09, 9.247173e-09, 9.197406e-09, 
    9.230481e-09, 9.175879e-09, 9.190813e-09, 9.07206e-09, 9.026813e-09, 
    9.007584e-09, 8.990749e-09, 8.949796e-09, 8.978078e-09, 8.966929e-09, 
    8.993451e-09, 9.010305e-09, 9.00197e-09, 9.053413e-09, 9.033413e-09, 
    9.138775e-09, 9.093393e-09, 9.211708e-09, 9.183396e-09, 9.218494e-09, 
    9.200584e-09, 9.231272e-09, 9.203653e-09, 9.251495e-09, 9.261913e-09, 
    9.254793e-09, 9.28214e-09, 9.202123e-09, 9.232853e-09, 9.001736e-09, 
    9.003095e-09, 9.009429e-09, 8.98159e-09, 8.979886e-09, 8.954373e-09, 
    8.977074e-09, 8.986742e-09, 9.011281e-09, 9.025798e-09, 9.039596e-09, 
    9.069935e-09, 9.103817e-09, 9.151195e-09, 9.185231e-09, 9.208047e-09, 
    9.194056e-09, 9.206408e-09, 9.1926e-09, 9.186129e-09, 9.258009e-09, 
    9.217648e-09, 9.278207e-09, 9.274856e-09, 9.247449e-09, 9.275233e-09, 
    9.00405e-09, 8.996227e-09, 8.969066e-09, 8.990322e-09, 8.951594e-09, 
    8.973273e-09, 8.985737e-09, 9.033832e-09, 9.044398e-09, 9.054197e-09, 
    9.073547e-09, 9.098382e-09, 9.141948e-09, 9.179852e-09, 9.214452e-09, 
    9.211917e-09, 9.21281e-09, 9.22054e-09, 9.201393e-09, 9.223683e-09, 
    9.227425e-09, 9.217643e-09, 9.274406e-09, 9.25819e-09, 9.274784e-09, 
    9.264225e-09, 8.99877e-09, 9.011933e-09, 9.00482e-09, 9.018196e-09, 
    9.008773e-09, 9.050674e-09, 9.063236e-09, 9.122018e-09, 9.097893e-09, 
    9.136287e-09, 9.101793e-09, 9.107906e-09, 9.137541e-09, 9.103656e-09, 
    9.177763e-09, 9.127523e-09, 9.22084e-09, 9.170673e-09, 9.223984e-09, 
    9.214303e-09, 9.230331e-09, 9.244688e-09, 9.262747e-09, 9.296071e-09, 
    9.288354e-09, 9.316222e-09, 9.031557e-09, 9.048631e-09, 9.047127e-09, 
    9.064994e-09, 9.078208e-09, 9.106848e-09, 9.152782e-09, 9.135508e-09, 
    9.167218e-09, 9.173585e-09, 9.125409e-09, 9.154989e-09, 9.060057e-09, 
    9.075396e-09, 9.066262e-09, 9.032904e-09, 9.13949e-09, 9.084791e-09, 
    9.185794e-09, 9.156163e-09, 9.24264e-09, 9.199635e-09, 9.284106e-09, 
    9.320219e-09, 9.354203e-09, 9.393921e-09, 9.057948e-09, 9.046347e-09, 
    9.067119e-09, 9.095858e-09, 9.122522e-09, 9.15797e-09, 9.161597e-09, 
    9.168238e-09, 9.185439e-09, 9.199902e-09, 9.170338e-09, 9.203528e-09, 
    9.078954e-09, 9.144237e-09, 9.041962e-09, 9.07276e-09, 9.094165e-09, 
    9.084775e-09, 9.133534e-09, 9.145026e-09, 9.191726e-09, 9.167585e-09, 
    9.311307e-09, 9.247721e-09, 9.42416e-09, 9.374854e-09, 9.042294e-09, 
    9.057908e-09, 9.112251e-09, 9.086395e-09, 9.160336e-09, 9.178537e-09, 
    9.193331e-09, 9.212246e-09, 9.214287e-09, 9.225493e-09, 9.20713e-09, 
    9.224768e-09, 9.158046e-09, 9.187862e-09, 9.106039e-09, 9.125954e-09, 
    9.116792e-09, 9.106743e-09, 9.137759e-09, 9.170805e-09, 9.171509e-09, 
    9.182105e-09, 9.211966e-09, 9.160636e-09, 9.319516e-09, 9.221399e-09, 
    9.074935e-09, 9.105011e-09, 9.109305e-09, 9.097655e-09, 9.176712e-09, 
    9.148067e-09, 9.22522e-09, 9.204368e-09, 9.238533e-09, 9.221556e-09, 
    9.219058e-09, 9.197254e-09, 9.183678e-09, 9.149381e-09, 9.121474e-09, 
    9.099344e-09, 9.10449e-09, 9.128799e-09, 9.172825e-09, 9.214473e-09, 
    9.205349e-09, 9.235936e-09, 9.154975e-09, 9.188924e-09, 9.175803e-09, 
    9.210016e-09, 9.135049e-09, 9.198891e-09, 9.118732e-09, 9.125759e-09, 
    9.147499e-09, 9.191228e-09, 9.2009e-09, 9.211231e-09, 9.204856e-09, 
    9.173942e-09, 9.168877e-09, 9.14697e-09, 9.140922e-09, 9.124229e-09, 
    9.110409e-09, 9.123036e-09, 9.136297e-09, 9.173955e-09, 9.207892e-09, 
    9.244892e-09, 9.253946e-09, 9.29718e-09, 9.261988e-09, 9.320063e-09, 
    9.270691e-09, 9.356155e-09, 9.202589e-09, 9.269236e-09, 9.148487e-09, 
    9.161496e-09, 9.185025e-09, 9.23899e-09, 9.209855e-09, 9.243927e-09, 
    9.168679e-09, 9.129638e-09, 9.119536e-09, 9.10069e-09, 9.119967e-09, 
    9.118399e-09, 9.136845e-09, 9.130917e-09, 9.175205e-09, 9.151416e-09, 
    9.218996e-09, 9.243657e-09, 9.313301e-09, 9.355995e-09, 9.399453e-09, 
    9.418638e-09, 9.424478e-09, 9.42692e-09 ;

 NFIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NFIX_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 OCDEP =
  3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 3.347111e-14, 
    3.347111e-14, 3.347111e-14, 3.347111e-14 ;

 O_SCALAR =
  0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 0.9666666, 
    0.9666666, 0.9666666,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 PARVEGLN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PBOT =
  102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 102587.8, 
    102587.8, 102587.8 ;

 PCH4 =
  0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 0.1743993, 
    0.1743993, 0.1743993 ;

 PCO2 =
  29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 29.20676, 
    29.20676, 29.20676 ;

 PFT_CTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_NTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PLANT_NDEMAND =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 POTENTIAL_IMMOB =
  4.718843e-14, 4.731617e-14, 4.729135e-14, 4.739429e-14, 4.733722e-14, 
    4.740459e-14, 4.721436e-14, 4.732122e-14, 4.725302e-14, 4.719996e-14, 
    4.759375e-14, 4.739888e-14, 4.779601e-14, 4.767194e-14, 4.798338e-14, 
    4.777668e-14, 4.802502e-14, 4.797746e-14, 4.812065e-14, 4.807965e-14, 
    4.826253e-14, 4.813958e-14, 4.835728e-14, 4.82332e-14, 4.82526e-14, 
    4.813551e-14, 4.743816e-14, 4.75695e-14, 4.743037e-14, 4.744911e-14, 
    4.744071e-14, 4.733838e-14, 4.728676e-14, 4.717869e-14, 4.719832e-14, 
    4.727771e-14, 4.745753e-14, 4.739655e-14, 4.755027e-14, 4.754681e-14, 
    4.77177e-14, 4.764068e-14, 4.792754e-14, 4.784611e-14, 4.808136e-14, 
    4.802223e-14, 4.807858e-14, 4.80615e-14, 4.80788e-14, 4.799207e-14, 
    4.802923e-14, 4.79529e-14, 4.76551e-14, 4.774269e-14, 4.748123e-14, 
    4.732369e-14, 4.721904e-14, 4.714469e-14, 4.715521e-14, 4.717524e-14, 
    4.727817e-14, 4.737491e-14, 4.744856e-14, 4.74978e-14, 4.754631e-14, 
    4.76929e-14, 4.77705e-14, 4.794399e-14, 4.791273e-14, 4.796571e-14, 
    4.801635e-14, 4.810127e-14, 4.80873e-14, 4.81247e-14, 4.796434e-14, 
    4.807092e-14, 4.789491e-14, 4.794307e-14, 4.755935e-14, 4.741301e-14, 
    4.735064e-14, 4.729612e-14, 4.716329e-14, 4.725503e-14, 4.721886e-14, 
    4.730491e-14, 4.735953e-14, 4.733252e-14, 4.749915e-14, 4.743439e-14, 
    4.77751e-14, 4.762847e-14, 4.801044e-14, 4.791915e-14, 4.803232e-14, 
    4.797459e-14, 4.807348e-14, 4.798448e-14, 4.813862e-14, 4.817214e-14, 
    4.814923e-14, 4.823726e-14, 4.797954e-14, 4.807857e-14, 4.733176e-14, 
    4.733616e-14, 4.735669e-14, 4.726641e-14, 4.726089e-14, 4.717814e-14, 
    4.725179e-14, 4.728313e-14, 4.73627e-14, 4.740972e-14, 4.745441e-14, 
    4.755261e-14, 4.766216e-14, 4.781523e-14, 4.792507e-14, 4.799865e-14, 
    4.795354e-14, 4.799337e-14, 4.794884e-14, 4.792798e-14, 4.815957e-14, 
    4.802957e-14, 4.82246e-14, 4.821382e-14, 4.812558e-14, 4.821504e-14, 
    4.733926e-14, 4.731391e-14, 4.722581e-14, 4.729476e-14, 4.716913e-14, 
    4.723945e-14, 4.727985e-14, 4.743571e-14, 4.746996e-14, 4.750167e-14, 
    4.756431e-14, 4.764462e-14, 4.778537e-14, 4.79077e-14, 4.80193e-14, 
    4.801113e-14, 4.801401e-14, 4.803891e-14, 4.797719e-14, 4.804904e-14, 
    4.806108e-14, 4.802957e-14, 4.821238e-14, 4.816018e-14, 4.821359e-14, 
    4.817961e-14, 4.732215e-14, 4.736481e-14, 4.734176e-14, 4.738509e-14, 
    4.735455e-14, 4.749024e-14, 4.753089e-14, 4.772097e-14, 4.764303e-14, 
    4.776708e-14, 4.765565e-14, 4.76754e-14, 4.777107e-14, 4.766168e-14, 
    4.790093e-14, 4.773873e-14, 4.803988e-14, 4.787804e-14, 4.805001e-14, 
    4.801882e-14, 4.807047e-14, 4.81167e-14, 4.817485e-14, 4.828204e-14, 
    4.825723e-14, 4.834684e-14, 4.742838e-14, 4.748364e-14, 4.74788e-14, 
    4.753663e-14, 4.757937e-14, 4.767199e-14, 4.782037e-14, 4.77646e-14, 
    4.786698e-14, 4.788749e-14, 4.773198e-14, 4.782748e-14, 4.752063e-14, 
    4.757023e-14, 4.754072e-14, 4.743272e-14, 4.777742e-14, 4.760063e-14, 
    4.792688e-14, 4.783129e-14, 4.81101e-14, 4.797148e-14, 4.824357e-14, 
    4.835962e-14, 4.846886e-14, 4.859624e-14, 4.751382e-14, 4.747628e-14, 
    4.754351e-14, 4.763642e-14, 4.772264e-14, 4.783712e-14, 4.784884e-14, 
    4.787026e-14, 4.792575e-14, 4.797239e-14, 4.787701e-14, 4.798408e-14, 
    4.758168e-14, 4.779276e-14, 4.746206e-14, 4.75617e-14, 4.763096e-14, 
    4.760061e-14, 4.775823e-14, 4.779534e-14, 4.794599e-14, 4.786817e-14, 
    4.833096e-14, 4.812642e-14, 4.869322e-14, 4.853509e-14, 4.746315e-14, 
    4.75137e-14, 4.768943e-14, 4.760585e-14, 4.784477e-14, 4.790347e-14, 
    4.795121e-14, 4.801216e-14, 4.801876e-14, 4.805486e-14, 4.79957e-14, 
    4.805254e-14, 4.783736e-14, 4.793356e-14, 4.766938e-14, 4.773373e-14, 
    4.770414e-14, 4.767166e-14, 4.777188e-14, 4.787851e-14, 4.788083e-14, 
    4.791497e-14, 4.801111e-14, 4.784574e-14, 4.835726e-14, 4.804153e-14, 
    4.75688e-14, 4.7666e-14, 4.767993e-14, 4.764228e-14, 4.789758e-14, 
    4.780515e-14, 4.805399e-14, 4.798679e-14, 4.809689e-14, 4.804219e-14, 
    4.803414e-14, 4.796385e-14, 4.792006e-14, 4.780938e-14, 4.771925e-14, 
    4.764775e-14, 4.766438e-14, 4.774291e-14, 4.788504e-14, 4.801934e-14, 
    4.798992e-14, 4.808852e-14, 4.782746e-14, 4.793696e-14, 4.789463e-14, 
    4.800499e-14, 4.776311e-14, 4.796898e-14, 4.771041e-14, 4.773311e-14, 
    4.780331e-14, 4.794436e-14, 4.797561e-14, 4.800889e-14, 4.798837e-14, 
    4.788862e-14, 4.787232e-14, 4.780162e-14, 4.778207e-14, 4.772817e-14, 
    4.768351e-14, 4.772431e-14, 4.776713e-14, 4.788868e-14, 4.799812e-14, 
    4.811735e-14, 4.814652e-14, 4.828552e-14, 4.817232e-14, 4.8359e-14, 
    4.820022e-14, 4.847499e-14, 4.798096e-14, 4.819564e-14, 4.780652e-14, 
    4.784852e-14, 4.792437e-14, 4.809829e-14, 4.800447e-14, 4.811421e-14, 
    4.787169e-14, 4.77456e-14, 4.771301e-14, 4.765209e-14, 4.77144e-14, 
    4.770933e-14, 4.776893e-14, 4.774978e-14, 4.789272e-14, 4.781598e-14, 
    4.803392e-14, 4.811335e-14, 4.833744e-14, 4.847456e-14, 4.861405e-14, 
    4.867555e-14, 4.869427e-14, 4.870209e-14 ;

 POT_F_DENIT =
  4.591369e-13, 4.602407e-13, 4.600251e-13, 4.609153e-13, 4.604209e-13, 
    4.610031e-13, 4.593583e-13, 4.602817e-13, 4.596915e-13, 4.592323e-13, 
    4.626387e-13, 4.609516e-13, 4.643875e-13, 4.633122e-13, 4.660095e-13, 
    4.642194e-13, 4.663697e-13, 4.659563e-13, 4.67197e-13, 4.668409e-13, 
    4.684274e-13, 4.673598e-13, 4.69248e-13, 4.681715e-13, 4.683395e-13, 
    4.673226e-13, 4.612939e-13, 4.62432e-13, 4.612257e-13, 4.61388e-13, 
    4.613146e-13, 4.604294e-13, 4.599836e-13, 4.590482e-13, 4.592172e-13, 
    4.599038e-13, 4.614579e-13, 4.609293e-13, 4.622581e-13, 4.622282e-13, 
    4.637064e-13, 4.630397e-13, 4.655233e-13, 4.648169e-13, 4.668552e-13, 
    4.663421e-13, 4.668304e-13, 4.666815e-13, 4.668311e-13, 4.660796e-13, 
    4.664007e-13, 4.657392e-13, 4.631699e-13, 4.639276e-13, 4.616649e-13, 
    4.603031e-13, 4.593971e-13, 4.587547e-13, 4.588446e-13, 4.590179e-13, 
    4.599069e-13, 4.607419e-13, 4.613785e-13, 4.618037e-13, 4.622226e-13, 
    4.63493e-13, 4.641635e-13, 4.656653e-13, 4.653937e-13, 4.658525e-13, 
    4.662906e-13, 4.670262e-13, 4.669048e-13, 4.672285e-13, 4.658378e-13, 
    4.66762e-13, 4.652353e-13, 4.656529e-13, 4.623423e-13, 4.610737e-13, 
    4.605354e-13, 4.600627e-13, 4.589141e-13, 4.597071e-13, 4.593941e-13, 
    4.601365e-13, 4.606085e-13, 4.603743e-13, 4.618148e-13, 4.612542e-13, 
    4.642026e-13, 4.62933e-13, 4.662401e-13, 4.654484e-13, 4.664283e-13, 
    4.659281e-13, 4.667845e-13, 4.66013e-13, 4.673482e-13, 4.676392e-13, 
    4.674395e-13, 4.682026e-13, 4.659675e-13, 4.668261e-13, 4.603703e-13, 
    4.604085e-13, 4.605853e-13, 4.598049e-13, 4.597569e-13, 4.59041e-13, 
    4.596767e-13, 4.599478e-13, 4.606346e-13, 4.610407e-13, 4.614265e-13, 
    4.62276e-13, 4.632239e-13, 4.645482e-13, 4.654992e-13, 4.661359e-13, 
    4.657448e-13, 4.660892e-13, 4.657033e-13, 4.655218e-13, 4.67529e-13, 
    4.664021e-13, 4.680917e-13, 4.679982e-13, 4.672328e-13, 4.680075e-13, 
    4.604344e-13, 4.602144e-13, 4.594533e-13, 4.600482e-13, 4.589622e-13, 
    4.595701e-13, 4.59919e-13, 4.612656e-13, 4.615606e-13, 4.618352e-13, 
    4.623762e-13, 4.630706e-13, 4.642891e-13, 4.65348e-13, 4.663143e-13, 
    4.662428e-13, 4.662676e-13, 4.664829e-13, 4.659478e-13, 4.665698e-13, 
    4.666738e-13, 4.664006e-13, 4.679844e-13, 4.675319e-13, 4.679945e-13, 
    4.676991e-13, 4.602852e-13, 4.606534e-13, 4.604535e-13, 4.608284e-13, 
    4.605636e-13, 4.617374e-13, 4.620885e-13, 4.637327e-13, 4.630569e-13, 
    4.641311e-13, 4.631651e-13, 4.633363e-13, 4.641653e-13, 4.63216e-13, 
    4.652885e-13, 4.638834e-13, 4.664908e-13, 4.650891e-13, 4.665777e-13, 
    4.663066e-13, 4.667536e-13, 4.671547e-13, 4.676578e-13, 4.685881e-13, 
    4.683717e-13, 4.691491e-13, 4.612025e-13, 4.616802e-13, 4.616376e-13, 
    4.621372e-13, 4.625066e-13, 4.63308e-13, 4.645922e-13, 4.641084e-13, 
    4.649944e-13, 4.651725e-13, 4.638245e-13, 4.64652e-13, 4.619955e-13, 
    4.624245e-13, 4.621683e-13, 4.612337e-13, 4.642164e-13, 4.626857e-13, 
    4.655097e-13, 4.646808e-13, 4.670963e-13, 4.658956e-13, 4.682529e-13, 
    4.692608e-13, 4.70207e-13, 4.713135e-13, 4.619404e-13, 4.616148e-13, 
    4.621957e-13, 4.630006e-13, 4.637453e-13, 4.647366e-13, 4.648373e-13, 
    4.650223e-13, 4.655024e-13, 4.659067e-13, 4.650803e-13, 4.660067e-13, 
    4.625241e-13, 4.64349e-13, 4.614864e-13, 4.623491e-13, 4.629469e-13, 
    4.626841e-13, 4.640474e-13, 4.643682e-13, 4.656732e-13, 4.649983e-13, 
    4.690111e-13, 4.672365e-13, 4.721543e-13, 4.707815e-13, 4.615008e-13, 
    4.619373e-13, 4.634578e-13, 4.627343e-13, 4.648014e-13, 4.653103e-13, 
    4.657226e-13, 4.662514e-13, 4.663073e-13, 4.666204e-13, 4.661064e-13, 
    4.665992e-13, 4.64734e-13, 4.655674e-13, 4.632789e-13, 4.638355e-13, 
    4.635789e-13, 4.632971e-13, 4.641641e-13, 4.650884e-13, 4.651072e-13, 
    4.654028e-13, 4.662382e-13, 4.648017e-13, 4.692391e-13, 4.664999e-13, 
    4.624134e-13, 4.632549e-13, 4.633741e-13, 4.630481e-13, 4.65258e-13, 
    4.644574e-13, 4.666128e-13, 4.660296e-13, 4.669832e-13, 4.665093e-13, 
    4.664385e-13, 4.658295e-13, 4.654492e-13, 4.644908e-13, 4.637094e-13, 
    4.630902e-13, 4.632332e-13, 4.639135e-13, 4.651436e-13, 4.663072e-13, 
    4.660519e-13, 4.669052e-13, 4.646426e-13, 4.655918e-13, 4.652242e-13, 
    4.6618e-13, 4.640938e-13, 4.658796e-13, 4.636368e-13, 4.638327e-13, 
    4.644402e-13, 4.65663e-13, 4.659318e-13, 4.662207e-13, 4.660414e-13, 
    4.65178e-13, 4.650357e-13, 4.644225e-13, 4.642529e-13, 4.63786e-13, 
    4.633985e-13, 4.637519e-13, 4.64122e-13, 4.651747e-13, 4.661225e-13, 
    4.671551e-13, 4.674075e-13, 4.686142e-13, 4.676318e-13, 4.692523e-13, 
    4.678748e-13, 4.702571e-13, 4.659811e-13, 4.678423e-13, 4.644678e-13, 
    4.648309e-13, 4.654887e-13, 4.669956e-13, 4.661809e-13, 4.671328e-13, 
    4.650298e-13, 4.639379e-13, 4.636544e-13, 4.631273e-13, 4.636656e-13, 
    4.636218e-13, 4.641371e-13, 4.639707e-13, 4.652084e-13, 4.645434e-13, 
    4.664311e-13, 4.6712e-13, 4.690628e-13, 4.702526e-13, 4.714627e-13, 
    4.719963e-13, 4.721587e-13, 4.722262e-13 ;

 POT_F_NIT =
  4.023214e-11, 4.057886e-11, 4.051132e-11, 4.079187e-11, 4.063611e-11, 
    4.081998e-11, 4.030228e-11, 4.059263e-11, 4.040715e-11, 4.026324e-11, 
    4.133912e-11, 4.080437e-11, 4.189836e-11, 4.155451e-11, 4.242101e-11, 
    4.184475e-11, 4.25377e-11, 4.240431e-11, 4.280638e-11, 4.269099e-11, 
    4.320742e-11, 4.285968e-11, 4.347637e-11, 4.312423e-11, 4.317922e-11, 
    4.284821e-11, 4.091171e-11, 4.127238e-11, 4.089039e-11, 4.094171e-11, 
    4.091867e-11, 4.063931e-11, 4.049891e-11, 4.020565e-11, 4.02588e-11, 
    4.047422e-11, 4.096476e-11, 4.079789e-11, 4.121908e-11, 4.120955e-11, 
    4.168104e-11, 4.146811e-11, 4.226472e-11, 4.20375e-11, 4.269579e-11, 
    4.252973e-11, 4.268798e-11, 4.263995e-11, 4.268859e-11, 4.24452e-11, 
    4.254938e-11, 4.233553e-11, 4.1508e-11, 4.175035e-11, 4.102967e-11, 
    4.059946e-11, 4.031498e-11, 4.011375e-11, 4.014215e-11, 4.019636e-11, 
    4.047548e-11, 4.073881e-11, 4.094008e-11, 4.1075e-11, 4.120816e-11, 
    4.161264e-11, 4.182751e-11, 4.231073e-11, 4.22233e-11, 4.237145e-11, 
    4.251323e-11, 4.275182e-11, 4.27125e-11, 4.281778e-11, 4.236751e-11, 
    4.266649e-11, 4.21735e-11, 4.230805e-11, 4.124449e-11, 4.084289e-11, 
    4.067284e-11, 4.052426e-11, 4.016401e-11, 4.041261e-11, 4.031451e-11, 
    4.054808e-11, 4.069686e-11, 4.062323e-11, 4.107869e-11, 4.09013e-11, 
    4.184026e-11, 4.143447e-11, 4.249669e-11, 4.224123e-11, 4.255802e-11, 
    4.239621e-11, 4.267365e-11, 4.24239e-11, 4.285699e-11, 4.29516e-11, 
    4.288693e-11, 4.313559e-11, 4.241006e-11, 4.268794e-11, 4.062119e-11, 
    4.06332e-11, 4.068913e-11, 4.044353e-11, 4.042853e-11, 4.020417e-11, 
    4.040376e-11, 4.048891e-11, 4.070548e-11, 4.083386e-11, 4.095609e-11, 
    4.122551e-11, 4.152749e-11, 4.195166e-11, 4.225776e-11, 4.246358e-11, 
    4.23373e-11, 4.244877e-11, 4.232417e-11, 4.226582e-11, 4.291613e-11, 
    4.255034e-11, 4.309977e-11, 4.306927e-11, 4.282025e-11, 4.307269e-11, 
    4.064162e-11, 4.057256e-11, 4.03333e-11, 4.052047e-11, 4.017977e-11, 
    4.03703e-11, 4.048006e-11, 4.090501e-11, 4.099867e-11, 4.108563e-11, 
    4.125765e-11, 4.147896e-11, 4.186868e-11, 4.220928e-11, 4.252147e-11, 
    4.249854e-11, 4.250661e-11, 4.257649e-11, 4.240348e-11, 4.260492e-11, 
    4.263878e-11, 4.255028e-11, 4.306517e-11, 4.291774e-11, 4.30686e-11, 
    4.297257e-11, 4.059499e-11, 4.071124e-11, 4.064839e-11, 4.076661e-11, 
    4.06833e-11, 4.105436e-11, 4.116595e-11, 4.169017e-11, 4.14746e-11, 
    4.181794e-11, 4.15094e-11, 4.156398e-11, 4.182917e-11, 4.152603e-11, 
    4.219046e-11, 4.17394e-11, 4.257921e-11, 4.212665e-11, 4.260764e-11, 
    4.252007e-11, 4.266509e-11, 4.279519e-11, 4.295914e-11, 4.326253e-11, 
    4.319216e-11, 4.344651e-11, 4.088486e-11, 4.103623e-11, 4.102288e-11, 
    4.118157e-11, 4.129914e-11, 4.155455e-11, 4.196589e-11, 4.181095e-11, 
    4.20956e-11, 4.215286e-11, 4.172048e-11, 4.198569e-11, 4.113765e-11, 
    4.127406e-11, 4.11928e-11, 4.089673e-11, 4.18466e-11, 4.135771e-11, 
    4.226277e-11, 4.19962e-11, 4.277662e-11, 4.238757e-11, 4.315346e-11, 
    4.348306e-11, 4.37944e-11, 4.415975e-11, 4.111896e-11, 4.101595e-11, 
    4.120045e-11, 4.145645e-11, 4.169467e-11, 4.201249e-11, 4.204507e-11, 
    4.210476e-11, 4.22596e-11, 4.239003e-11, 4.212365e-11, 4.242274e-11, 
    4.130574e-11, 4.188917e-11, 4.0977e-11, 4.125059e-11, 4.144127e-11, 
    4.135756e-11, 4.17932e-11, 4.189622e-11, 4.231622e-11, 4.209883e-11, 
    4.340158e-11, 4.282267e-11, 4.443895e-11, 4.398416e-11, 4.098e-11, 
    4.111858e-11, 4.160281e-11, 4.137205e-11, 4.203373e-11, 4.219744e-11, 
    4.233075e-11, 4.25015e-11, 4.251995e-11, 4.262131e-11, 4.245526e-11, 
    4.261473e-11, 4.201312e-11, 4.228141e-11, 4.154726e-11, 4.172533e-11, 
    4.164335e-11, 4.155353e-11, 4.183105e-11, 4.212779e-11, 4.213412e-11, 
    4.22295e-11, 4.249891e-11, 4.203634e-11, 4.34766e-11, 4.258418e-11, 
    4.126998e-11, 4.153812e-11, 4.157647e-11, 4.147245e-11, 4.2181e-11, 
    4.192355e-11, 4.261883e-11, 4.243033e-11, 4.27394e-11, 4.258567e-11, 
    4.256306e-11, 4.23661e-11, 4.22437e-11, 4.19353e-11, 4.168523e-11, 
    4.148747e-11, 4.15334e-11, 4.175078e-11, 4.214596e-11, 4.252157e-11, 
    4.243914e-11, 4.271581e-11, 4.198548e-11, 4.229093e-11, 4.217273e-11, 
    4.248127e-11, 4.180683e-11, 4.238091e-11, 4.166073e-11, 4.172361e-11, 
    4.191843e-11, 4.231177e-11, 4.239901e-11, 4.249231e-11, 4.243472e-11, 
    4.215604e-11, 4.211047e-11, 4.191366e-11, 4.185941e-11, 4.170987e-11, 
    4.158628e-11, 4.169919e-11, 4.181793e-11, 4.215612e-11, 4.246209e-11, 
    4.279699e-11, 4.287915e-11, 4.327258e-11, 4.295218e-11, 4.348158e-11, 
    4.303129e-11, 4.381227e-11, 4.241427e-11, 4.301816e-11, 4.192731e-11, 
    4.204412e-11, 4.225585e-11, 4.274352e-11, 4.247986e-11, 4.278828e-11, 
    4.210868e-11, 4.175831e-11, 4.166788e-11, 4.149948e-11, 4.167173e-11, 
    4.16577e-11, 4.182285e-11, 4.176973e-11, 4.216736e-11, 4.195353e-11, 
    4.256244e-11, 4.278579e-11, 4.341977e-11, 4.381081e-11, 4.421071e-11, 
    4.438786e-11, 4.444185e-11, 4.446443e-11 ;

 PROD100C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHA =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHADE_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Q2M =
  0.001212909, 0.001212836, 0.00121285, 0.001212792, 0.001212823, 
    0.001212786, 0.001212894, 0.001212834, 0.001212872, 0.001212902, 
    0.001212681, 0.001212789, 0.001212563, 0.001212633, 0.001212454, 
    0.001212575, 0.00121243, 0.001212456, 0.001212374, 0.001212398, 
    0.001212296, 0.001212363, 0.001212241, 0.001212311, 0.001212301, 
    0.001212366, 0.001212766, 0.001212695, 0.00121277, 0.00121276, 
    0.001212764, 0.001212823, 0.001212854, 0.001212914, 0.001212902, 
    0.001212858, 0.001212756, 0.001212789, 0.001212701, 0.001212703, 
    0.001212607, 0.00121265, 0.001212485, 0.001212533, 0.001212397, 
    0.001212431, 0.001212399, 0.001212408, 0.001212398, 0.001212448, 
    0.001212427, 0.00121247, 0.001212642, 0.001212593, 0.001212742, 
    0.001212833, 0.001212891, 0.001212933, 0.001212927, 0.001212916, 
    0.001212858, 0.001212802, 0.00121276, 0.001212731, 0.001212704, 
    0.001212623, 0.001212578, 0.001212476, 0.001212493, 0.001212464, 
    0.001212434, 0.001212386, 0.001212394, 0.001212373, 0.001212464, 
    0.001212404, 0.001212503, 0.001212476, 0.001212701, 0.00121278, 
    0.001212818, 0.001212847, 0.001212923, 0.001212871, 0.001212891, 
    0.001212842, 0.001212811, 0.001212826, 0.001212731, 0.001212768, 
    0.001212575, 0.001212658, 0.001212438, 0.00121249, 0.001212425, 
    0.001212458, 0.001212402, 0.001212452, 0.001212364, 0.001212346, 
    0.001212359, 0.001212308, 0.001212455, 0.001212399, 0.001212826, 
    0.001212824, 0.001212812, 0.001212865, 0.001212867, 0.001212914, 
    0.001212872, 0.001212855, 0.001212808, 0.001212782, 0.001212756, 
    0.001212701, 0.001212639, 0.001212551, 0.001212486, 0.001212444, 
    0.00121247, 0.001212447, 0.001212472, 0.001212484, 0.001212353, 
    0.001212427, 0.001212315, 0.001212321, 0.001212372, 0.001212321, 
    0.001212822, 0.001212836, 0.001212887, 0.001212847, 0.001212919, 
    0.00121288, 0.001212857, 0.001212768, 0.001212747, 0.00121273, 
    0.001212694, 0.001212648, 0.001212568, 0.001212497, 0.001212432, 
    0.001212437, 0.001212435, 0.001212421, 0.001212456, 0.001212415, 
    0.001212409, 0.001212426, 0.001212322, 0.001212352, 0.001212321, 
    0.001212341, 0.001212832, 0.001212807, 0.001212821, 0.001212796, 
    0.001212814, 0.001212737, 0.001212714, 0.001212606, 0.001212649, 
    0.001212579, 0.001212642, 0.001212631, 0.001212579, 0.001212638, 
    0.001212501, 0.001212596, 0.001212421, 0.001212517, 0.001212415, 
    0.001212432, 0.001212403, 0.001212377, 0.001212343, 0.001212283, 
    0.001212297, 0.001212246, 0.001212771, 0.00121274, 0.001212742, 
    0.001212709, 0.001212685, 0.001212632, 0.001212548, 0.001212579, 
    0.001212521, 0.001212508, 0.001212598, 0.001212544, 0.001212719, 
    0.001212692, 0.001212707, 0.001212769, 0.001212573, 0.001212674, 
    0.001212485, 0.001212541, 0.001212381, 0.001212461, 0.001212305, 
    0.00121224, 0.001212176, 0.001212105, 0.001212723, 0.001212744, 
    0.001212705, 0.001212654, 0.001212604, 0.001212538, 0.001212531, 
    0.001212519, 0.001212485, 0.001212459, 0.001212516, 0.001212452, 
    0.001212687, 0.001212564, 0.001212752, 0.001212697, 0.001212656, 
    0.001212673, 0.001212583, 0.001212562, 0.001212475, 0.00121252, 
    0.001212257, 0.001212373, 0.001212049, 0.00121214, 0.001212751, 
    0.001212722, 0.001212623, 0.00121267, 0.001212533, 0.001212499, 
    0.001212471, 0.001212437, 0.001212433, 0.001212412, 0.001212446, 
    0.001212413, 0.001212538, 0.001212481, 0.001212633, 0.001212597, 
    0.001212614, 0.001212632, 0.001212575, 0.001212516, 0.001212513, 
    0.001212492, 0.001212442, 0.001212533, 0.001212245, 0.001212424, 
    0.001212691, 0.001212637, 0.001212628, 0.001212649, 0.001212502, 
    0.001212556, 0.001212413, 0.001212451, 0.001212388, 0.001212419, 
    0.001212424, 0.001212464, 0.001212489, 0.001212554, 0.001212606, 
    0.001212646, 0.001212636, 0.001212592, 0.001212512, 0.001212433, 
    0.00121245, 0.001212393, 0.001212543, 0.00121248, 0.001212504, 
    0.001212441, 0.00121258, 0.001212465, 0.00121261, 0.001212597, 
    0.001212557, 0.001212477, 0.001212457, 0.001212439, 0.00121245, 
    0.001212508, 0.001212518, 0.001212558, 0.00121257, 0.0012126, 
    0.001212625, 0.001212602, 0.001212579, 0.001212507, 0.001212445, 
    0.001212377, 0.00121236, 0.001212284, 0.001212347, 0.001212244, 
    0.001212335, 0.001212176, 0.001212457, 0.001212335, 0.001212555, 
    0.001212531, 0.001212488, 0.001212389, 0.001212441, 0.00121238, 
    0.001212518, 0.001212591, 0.001212609, 0.001212643, 0.001212608, 
    0.001212611, 0.001212577, 0.001212587, 0.001212505, 0.00121255, 
    0.001212424, 0.00121238, 0.001212252, 0.001212174, 0.001212093, 
    0.001212058, 0.001212047, 0.001212043 ;

 QBOT =
  0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224, 0.001329224, 0.001329224, 
    0.001329224, 0.001329224, 0.001329224 ;

 QCHARGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_PERCH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_XS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRIP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLOOD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_ICE_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_LIQ_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINFL =
  -1.570073e-07, -1.573053e-07, -1.57247e-07, -1.574879e-07, -1.573538e-07, 
    -1.575118e-07, -1.570671e-07, -1.573176e-07, -1.571574e-07, 
    -1.570333e-07, -1.579554e-07, -1.574984e-07, -1.584228e-07, 
    -1.581334e-07, -1.58861e-07, -1.583786e-07, -1.589571e-07, -1.588458e-07, 
    -1.591774e-07, -1.590824e-07, -1.595086e-07, -1.592212e-07, 
    -1.597269e-07, -1.594393e-07, -1.594848e-07, -1.592119e-07, 
    -1.575892e-07, -1.57899e-07, -1.575712e-07, -1.576153e-07, -1.575952e-07, 
    -1.573571e-07, -1.572378e-07, -1.569835e-07, -1.570295e-07, 
    -1.572157e-07, -1.576351e-07, -1.57492e-07, -1.578496e-07, -1.578415e-07, 
    -1.582395e-07, -1.580602e-07, -1.5873e-07, -1.585373e-07, -1.590863e-07, 
    -1.589494e-07, -1.590801e-07, -1.590403e-07, -1.590806e-07, 
    -1.588798e-07, -1.589659e-07, -1.587886e-07, -1.580941e-07, -1.58298e-07, 
    -1.576898e-07, -1.573248e-07, -1.570784e-07, -1.569043e-07, 
    -1.569289e-07, -1.569761e-07, -1.572168e-07, -1.574416e-07, -1.57613e-07, 
    -1.577277e-07, -1.578404e-07, -1.581847e-07, -1.583635e-07, -1.58769e-07, 
    -1.586953e-07, -1.588192e-07, -1.589357e-07, -1.591329e-07, 
    -1.591003e-07, -1.591873e-07, -1.58815e-07, -1.59063e-07, -1.586536e-07, 
    -1.587658e-07, -1.578757e-07, -1.575305e-07, -1.573873e-07, 
    -1.572584e-07, -1.569479e-07, -1.571627e-07, -1.570782e-07, 
    -1.572782e-07, -1.574058e-07, -1.573425e-07, -1.577308e-07, 
    -1.575802e-07, -1.583742e-07, -1.580326e-07, -1.589222e-07, 
    -1.587103e-07, -1.589727e-07, -1.588386e-07, -1.590687e-07, 
    -1.588616e-07, -1.592193e-07, -1.592976e-07, -1.592442e-07, 
    -1.594477e-07, -1.588503e-07, -1.590806e-07, -1.573409e-07, 
    -1.573513e-07, -1.57399e-07, -1.571893e-07, -1.571762e-07, -1.569825e-07, 
    -1.571545e-07, -1.57228e-07, -1.574128e-07, -1.575229e-07, -1.57627e-07, 
    -1.578556e-07, -1.581112e-07, -1.584667e-07, -1.587241e-07, 
    -1.588945e-07, -1.587897e-07, -1.588823e-07, -1.58779e-07, -1.587304e-07, 
    -1.592686e-07, -1.58967e-07, -1.594185e-07, -1.593934e-07, -1.591896e-07, 
    -1.593962e-07, -1.573585e-07, -1.57299e-07, -1.57094e-07, -1.572545e-07, 
    -1.569613e-07, -1.571261e-07, -1.57221e-07, -1.575844e-07, -1.576629e-07, 
    -1.577371e-07, -1.578825e-07, -1.580695e-07, -1.583972e-07, 
    -1.586843e-07, -1.589423e-07, -1.589234e-07, -1.589301e-07, 
    -1.589882e-07, -1.588449e-07, -1.590116e-07, -1.5904e-07, -1.589664e-07, 
    -1.5939e-07, -1.592691e-07, -1.593928e-07, -1.59314e-07, -1.573182e-07, 
    -1.57418e-07, -1.573642e-07, -1.574656e-07, -1.573945e-07, -1.577116e-07, 
    -1.578065e-07, -1.582484e-07, -1.58066e-07, -1.583549e-07, -1.58095e-07, 
    -1.581414e-07, -1.583663e-07, -1.581088e-07, -1.586696e-07, 
    -1.582903e-07, -1.589904e-07, -1.586142e-07, -1.590139e-07, 
    -1.589412e-07, -1.59061e-07, -1.591686e-07, -1.593031e-07, -1.595524e-07, 
    -1.594945e-07, -1.597019e-07, -1.575662e-07, -1.576956e-07, 
    -1.576834e-07, -1.578181e-07, -1.579179e-07, -1.581328e-07, -1.58478e-07, 
    -1.58348e-07, -1.585856e-07, -1.586369e-07, -1.58272e-07, -1.58495e-07, 
    -1.577815e-07, -1.578979e-07, -1.57828e-07, -1.575769e-07, -1.583792e-07, 
    -1.579685e-07, -1.587285e-07, -1.585031e-07, -1.591534e-07, 
    -1.588329e-07, -1.594628e-07, -1.597336e-07, -1.599839e-07, 
    -1.602806e-07, -1.577653e-07, -1.576774e-07, -1.578339e-07, 
    -1.580517e-07, -1.582509e-07, -1.585169e-07, -1.585436e-07, 
    -1.585936e-07, -1.587253e-07, -1.588336e-07, -1.586102e-07, 
    -1.588607e-07, -1.579267e-07, -1.584144e-07, -1.57645e-07, -1.578783e-07, 
    -1.580384e-07, -1.579673e-07, -1.583329e-07, -1.584193e-07, 
    -1.587733e-07, -1.585883e-07, -1.596676e-07, -1.591926e-07, 
    -1.605032e-07, -1.601387e-07, -1.57647e-07, -1.577646e-07, -1.581744e-07, 
    -1.579794e-07, -1.585341e-07, -1.586741e-07, -1.587843e-07, 
    -1.589266e-07, -1.589412e-07, -1.590253e-07, -1.588876e-07, 
    -1.590196e-07, -1.585174e-07, -1.587437e-07, -1.581265e-07, 
    -1.582767e-07, -1.582073e-07, -1.581319e-07, -1.583647e-07, 
    -1.586139e-07, -1.586178e-07, -1.587012e-07, -1.589291e-07, 
    -1.585363e-07, -1.597314e-07, -1.589989e-07, -1.578928e-07, 
    -1.581208e-07, -1.581516e-07, -1.580636e-07, -1.586604e-07, 
    -1.584425e-07, -1.590231e-07, -1.58867e-07, -1.591223e-07, -1.589956e-07, 
    -1.58977e-07, -1.588138e-07, -1.587125e-07, -1.584526e-07, -1.582432e-07, 
    -1.580762e-07, -1.581149e-07, -1.582983e-07, -1.586288e-07, 
    -1.589432e-07, -1.588753e-07, -1.591029e-07, -1.58494e-07, -1.587523e-07, 
    -1.586542e-07, -1.589095e-07, -1.583449e-07, -1.588306e-07, 
    -1.582218e-07, -1.582747e-07, -1.584382e-07, -1.587705e-07, 
    -1.588411e-07, -1.58919e-07, -1.588706e-07, -1.586402e-07, -1.585986e-07, 
    -1.584339e-07, -1.583891e-07, -1.582631e-07, -1.581594e-07, 
    -1.582545e-07, -1.583547e-07, -1.586398e-07, -1.588941e-07, 
    -1.591704e-07, -1.592374e-07, -1.59563e-07, -1.592999e-07, -1.597357e-07, 
    -1.593682e-07, -1.600023e-07, -1.588564e-07, -1.593546e-07, 
    -1.584452e-07, -1.585427e-07, -1.587237e-07, -1.591277e-07, 
    -1.589082e-07, -1.591641e-07, -1.585969e-07, -1.583053e-07, -1.58228e-07, 
    -1.580866e-07, -1.582312e-07, -1.582194e-07, -1.583578e-07, 
    -1.583133e-07, -1.586491e-07, -1.584672e-07, -1.589769e-07, 
    -1.591618e-07, -1.596807e-07, -1.599988e-07, -1.603197e-07, 
    -1.604618e-07, -1.605049e-07, -1.60523e-07 ;

 QINTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QIRRIG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRGWL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 QRUNOFF_NODYNLNDUSE =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 QRUNOFF_R =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 QRUNOFF_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QSNOMELT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSOIL =
  3.281309e-06, 3.287373e-06, 3.286193e-06, 3.291092e-06, 3.288374e-06, 
    3.291583e-06, 3.282538e-06, 3.287613e-06, 3.284372e-06, 3.281855e-06, 
    3.300584e-06, 3.291311e-06, 3.310249e-06, 3.304315e-06, 3.31989e-06, 
    3.309323e-06, 3.3219e-06, 3.319605e-06, 3.326525e-06, 3.324541e-06, 
    3.333406e-06, 3.327441e-06, 3.338018e-06, 3.331982e-06, 3.332924e-06, 
    3.327244e-06, 3.293179e-06, 3.299427e-06, 3.292809e-06, 3.293699e-06, 
    3.2933e-06, 3.288429e-06, 3.285975e-06, 3.280847e-06, 3.281778e-06, 
    3.285545e-06, 3.2941e-06, 3.2912e-06, 3.298512e-06, 3.298346e-06, 
    3.306501e-06, 3.302822e-06, 3.3172e-06, 3.312652e-06, 3.324624e-06, 
    3.321766e-06, 3.324489e-06, 3.323663e-06, 3.3245e-06, 3.32031e-06, 
    3.322104e-06, 3.318421e-06, 3.30351e-06, 3.307696e-06, 3.295226e-06, 
    3.28773e-06, 3.28276e-06, 3.279238e-06, 3.279735e-06, 3.280684e-06, 
    3.285567e-06, 3.290168e-06, 3.293673e-06, 3.296014e-06, 3.298322e-06, 
    3.305315e-06, 3.309027e-06, 3.317992e-06, 3.316487e-06, 3.319039e-06, 
    3.321482e-06, 3.325587e-06, 3.324911e-06, 3.326721e-06, 3.318973e-06, 
    3.324119e-06, 3.31563e-06, 3.317948e-06, 3.298944e-06, 3.291984e-06, 
    3.289013e-06, 3.28642e-06, 3.280118e-06, 3.284468e-06, 3.282752e-06, 
    3.286837e-06, 3.289436e-06, 3.288151e-06, 3.296078e-06, 3.293e-06, 
    3.309248e-06, 3.302239e-06, 3.321197e-06, 3.316796e-06, 3.322254e-06, 
    3.319467e-06, 3.324242e-06, 3.319944e-06, 3.327395e-06, 3.329019e-06, 
    3.327909e-06, 3.332179e-06, 3.319706e-06, 3.324488e-06, 3.288114e-06, 
    3.288324e-06, 3.289301e-06, 3.285008e-06, 3.284747e-06, 3.280822e-06, 
    3.284314e-06, 3.285802e-06, 3.289587e-06, 3.291827e-06, 3.293951e-06, 
    3.298623e-06, 3.303847e-06, 3.311171e-06, 3.317081e-06, 3.320628e-06, 
    3.318453e-06, 3.320373e-06, 3.318226e-06, 3.317221e-06, 3.32841e-06, 
    3.32212e-06, 3.331565e-06, 3.331041e-06, 3.326763e-06, 3.331101e-06, 
    3.288471e-06, 3.287265e-06, 3.283081e-06, 3.286355e-06, 3.280395e-06, 
    3.283728e-06, 3.285646e-06, 3.293063e-06, 3.29469e-06, 3.296198e-06, 
    3.29918e-06, 3.30301e-06, 3.30974e-06, 3.316245e-06, 3.321625e-06, 
    3.32123e-06, 3.321369e-06, 3.322572e-06, 3.319593e-06, 3.323061e-06, 
    3.323643e-06, 3.322121e-06, 3.330971e-06, 3.32844e-06, 3.33103e-06, 
    3.329382e-06, 3.287657e-06, 3.289687e-06, 3.28859e-06, 3.290653e-06, 
    3.289199e-06, 3.295654e-06, 3.297588e-06, 3.306657e-06, 3.302934e-06, 
    3.308864e-06, 3.303536e-06, 3.304479e-06, 3.309054e-06, 3.303825e-06, 
    3.315919e-06, 3.307506e-06, 3.322619e-06, 3.314185e-06, 3.323108e-06, 
    3.321602e-06, 3.324097e-06, 3.326333e-06, 3.329151e-06, 3.334355e-06, 
    3.333149e-06, 3.337509e-06, 3.292714e-06, 3.29534e-06, 3.29511e-06, 
    3.297862e-06, 3.299898e-06, 3.304317e-06, 3.311417e-06, 3.308745e-06, 
    3.313655e-06, 3.315273e-06, 3.307184e-06, 3.311759e-06, 3.2971e-06, 
    3.299462e-06, 3.298057e-06, 3.292921e-06, 3.309359e-06, 3.300911e-06, 
    3.317168e-06, 3.311941e-06, 3.326014e-06, 3.319317e-06, 3.332485e-06, 
    3.33813e-06, 3.343464e-06, 3.3497e-06, 3.296776e-06, 3.29499e-06, 
    3.298189e-06, 3.302619e-06, 3.306737e-06, 3.312221e-06, 3.312784e-06, 
    3.313812e-06, 3.317114e-06, 3.319361e-06, 3.314136e-06, 3.319925e-06, 
    3.300008e-06, 3.310094e-06, 3.294314e-06, 3.299056e-06, 3.302358e-06, 
    3.300911e-06, 3.30844e-06, 3.310218e-06, 3.318088e-06, 3.313711e-06, 
    3.336734e-06, 3.326803e-06, 3.354465e-06, 3.346703e-06, 3.294366e-06, 
    3.29677e-06, 3.305149e-06, 3.301161e-06, 3.312588e-06, 3.316041e-06, 
    3.31834e-06, 3.32128e-06, 3.321599e-06, 3.323343e-06, 3.320485e-06, 
    3.32323e-06, 3.312233e-06, 3.31749e-06, 3.304192e-06, 3.307267e-06, 
    3.305852e-06, 3.304301e-06, 3.309093e-06, 3.314208e-06, 3.314319e-06, 
    3.316594e-06, 3.321227e-06, 3.312635e-06, 3.338013e-06, 3.322695e-06, 
    3.299394e-06, 3.304031e-06, 3.304696e-06, 3.302898e-06, 3.315758e-06, 
    3.310688e-06, 3.3233e-06, 3.320056e-06, 3.325375e-06, 3.32273e-06, 
    3.322341e-06, 3.318949e-06, 3.31684e-06, 3.310891e-06, 3.306575e-06, 
    3.303159e-06, 3.303953e-06, 3.307707e-06, 3.314521e-06, 3.321627e-06, 
    3.320206e-06, 3.32497e-06, 3.311758e-06, 3.317653e-06, 3.315615e-06, 
    3.320934e-06, 3.308674e-06, 3.319195e-06, 3.306152e-06, 3.307238e-06, 
    3.3106e-06, 3.318009e-06, 3.319517e-06, 3.321122e-06, 3.320132e-06, 
    3.315326e-06, 3.313911e-06, 3.310519e-06, 3.309582e-06, 3.307002e-06, 
    3.304867e-06, 3.306817e-06, 3.308866e-06, 3.31533e-06, 3.320602e-06, 
    3.326365e-06, 3.327778e-06, 3.334523e-06, 3.329026e-06, 3.338098e-06, 
    3.330377e-06, 3.34376e-06, 3.319773e-06, 3.330157e-06, 3.310754e-06, 
    3.312768e-06, 3.317046e-06, 3.325442e-06, 3.320909e-06, 3.326212e-06, 
    3.31388e-06, 3.307835e-06, 3.306276e-06, 3.303366e-06, 3.306343e-06, 
    3.306101e-06, 3.308952e-06, 3.308036e-06, 3.315524e-06, 3.311207e-06, 
    3.32233e-06, 3.326171e-06, 3.337051e-06, 3.343741e-06, 3.350576e-06, 
    3.353596e-06, 3.354517e-06, 3.354901e-06 ;

 QVEGE =
  -7.794841e-07, -7.79042e-07, -7.791259e-07, -7.787729e-07, -7.789655e-07, 
    -7.787367e-07, -7.793906e-07, -7.790279e-07, -7.792572e-07, 
    -7.794388e-07, -7.78096e-07, -7.787561e-07, -7.773739e-07, -7.777994e-07, 
    -7.767172e-07, -7.774458e-07, -7.765674e-07, -7.767291e-07, 
    -7.762188e-07, -7.763647e-07, -7.757282e-07, -7.761512e-07, 
    -7.753808e-07, -7.758244e-07, -7.757587e-07, -7.761666e-07, 
    -7.786148e-07, -7.781815e-07, -7.786426e-07, -7.785804e-07, 
    -7.786062e-07, -7.789647e-07, -7.791508e-07, -7.795115e-07, 
    -7.794445e-07, -7.79176e-07, -7.785522e-07, -7.787584e-07, -7.782199e-07, 
    -7.782319e-07, -7.776392e-07, -7.779057e-07, -7.769053e-07, 
    -7.771869e-07, -7.763584e-07, -7.765695e-07, -7.7637e-07, -7.764294e-07, 
    -7.763692e-07, -7.766781e-07, -7.765464e-07, -7.768146e-07, 
    -7.778575e-07, -7.775543e-07, -7.784668e-07, -7.790281e-07, 
    -7.793763e-07, -7.796294e-07, -7.795937e-07, -7.795274e-07, 
    -7.791747e-07, -7.788337e-07, -7.785758e-07, -7.784044e-07, 
    -7.782338e-07, -7.777424e-07, -7.774631e-07, -7.768522e-07, 
    -7.769553e-07, -7.767745e-07, -7.765901e-07, -7.762903e-07, 
    -7.763385e-07, -7.76208e-07, -7.767736e-07, -7.76401e-07, -7.770158e-07, 
    -7.768492e-07, -7.782187e-07, -7.787013e-07, -7.789326e-07, 
    -7.791109e-07, -7.795669e-07, -7.792539e-07, -7.793782e-07, 
    -7.790758e-07, -7.788876e-07, -7.789794e-07, -7.783996e-07, 
    -7.786267e-07, -7.774465e-07, -7.77953e-07, -7.766116e-07, -7.769335e-07, 
    -7.765331e-07, -7.767362e-07, -7.763905e-07, -7.767015e-07, 
    -7.761569e-07, -7.760414e-07, -7.76121e-07, -7.75804e-07, -7.767196e-07, 
    -7.76373e-07, -7.789835e-07, -7.789687e-07, -7.788961e-07, -7.792152e-07, 
    -7.792329e-07, -7.795149e-07, -7.792612e-07, -7.791555e-07, 
    -7.788742e-07, -7.787132e-07, -7.785578e-07, -7.782148e-07, 
    -7.778372e-07, -7.773019e-07, -7.769131e-07, -7.766513e-07, 
    -7.768098e-07, -7.766702e-07, -7.768275e-07, -7.768998e-07, 
    -7.760867e-07, -7.76547e-07, -7.758497e-07, -7.758874e-07, -7.762062e-07, 
    -7.758831e-07, -7.789578e-07, -7.790438e-07, -7.793519e-07, 
    -7.791108e-07, -7.795451e-07, -7.793062e-07, -7.791709e-07, 
    -7.786287e-07, -7.785017e-07, -7.783935e-07, -7.781721e-07, 
    -7.778922e-07, -7.774054e-07, -7.769772e-07, -7.765781e-07, 
    -7.766068e-07, -7.765969e-07, -7.765108e-07, -7.767284e-07, 
    -7.764747e-07, -7.764351e-07, -7.765433e-07, -7.758926e-07, 
    -7.760787e-07, -7.758882e-07, -7.760086e-07, -7.790151e-07, 
    -7.788687e-07, -7.789483e-07, -7.788003e-07, -7.789071e-07, 
    -7.784403e-07, -7.783e-07, -7.776356e-07, -7.778995e-07, -7.774707e-07, 
    -7.778534e-07, -7.777874e-07, -7.774699e-07, -7.778307e-07, -7.77007e-07, 
    -7.775773e-07, -7.765074e-07, -7.770926e-07, -7.764712e-07, 
    -7.765798e-07, -7.763967e-07, -7.762357e-07, -7.760269e-07, 
    -7.756493e-07, -7.757357e-07, -7.754137e-07, -7.786472e-07, 
    -7.784595e-07, -7.784702e-07, -7.782692e-07, -7.781215e-07, 
    -7.777953e-07, -7.772802e-07, -7.774724e-07, -7.77113e-07, -7.770449e-07, 
    -7.775852e-07, -7.77258e-07, -7.783292e-07, -7.781616e-07, -7.782571e-07, 
    -7.786359e-07, -7.774362e-07, -7.780541e-07, -7.769077e-07, 
    -7.772405e-07, -7.762595e-07, -7.767561e-07, -7.757845e-07, -7.75381e-07, 
    -7.749713e-07, -7.745226e-07, -7.783505e-07, -7.784789e-07, 
    -7.782435e-07, -7.779284e-07, -7.776214e-07, -7.772213e-07, -7.77177e-07, 
    -7.771037e-07, -7.769081e-07, -7.767444e-07, -7.770861e-07, 
    -7.767027e-07, -7.781346e-07, -7.773798e-07, -7.785329e-07, 
    -7.781929e-07, -7.779443e-07, -7.780471e-07, -7.774929e-07, 
    -7.773641e-07, -7.768435e-07, -7.771086e-07, -7.75486e-07, -7.762101e-07, 
    -7.74159e-07, -7.747416e-07, -7.785252e-07, -7.783481e-07, -7.777408e-07, 
    -7.780278e-07, -7.771914e-07, -7.769895e-07, -7.768181e-07, 
    -7.766081e-07, -7.76581e-07, -7.764555e-07, -7.766618e-07, -7.764614e-07, 
    -7.772204e-07, -7.768824e-07, -7.778028e-07, -7.775826e-07, 
    -7.776819e-07, -7.777951e-07, -7.77446e-07, -7.770822e-07, -7.770649e-07, 
    -7.769518e-07, -7.766429e-07, -7.771878e-07, -7.754098e-07, 
    -7.765307e-07, -7.781553e-07, -7.778274e-07, -7.777693e-07, 
    -7.778978e-07, -7.770103e-07, -7.773325e-07, -7.764572e-07, 
    -7.766933e-07, -7.763036e-07, -7.764983e-07, -7.765274e-07, 
    -7.767744e-07, -7.769304e-07, -7.773194e-07, -7.77634e-07, -7.77878e-07, 
    -7.778204e-07, -7.775521e-07, -7.770578e-07, -7.765828e-07, 
    -7.766889e-07, -7.763331e-07, -7.772525e-07, -7.768745e-07, 
    -7.770248e-07, -7.766307e-07, -7.774797e-07, -7.767863e-07, 
    -7.776599e-07, -7.775815e-07, -7.773389e-07, -7.768551e-07, -7.76733e-07, 
    -7.766196e-07, -7.766876e-07, -7.770455e-07, -7.770976e-07, 
    -7.773424e-07, -7.774146e-07, -7.775978e-07, -7.777537e-07, 
    -7.776137e-07, -7.774684e-07, -7.770414e-07, -7.766583e-07, 
    -7.762349e-07, -7.761272e-07, -7.756528e-07, -7.760524e-07, 
    -7.754055e-07, -7.759758e-07, -7.749758e-07, -7.767318e-07, -7.75973e-07, 
    -7.773246e-07, -7.771775e-07, -7.769233e-07, -7.763114e-07, 
    -7.766324e-07, -7.762523e-07, -7.77099e-07, -7.775477e-07, -7.776516e-07, 
    -7.778649e-07, -7.776467e-07, -7.776641e-07, -7.774556e-07, 
    -7.775221e-07, -7.77027e-07, -7.772918e-07, -7.765307e-07, -7.762529e-07, 
    -7.75451e-07, -7.749613e-07, -7.744441e-07, -7.742199e-07, -7.741506e-07, 
    -7.741223e-07 ;

 QVEGT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RETRANSN =
  4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 4.500845e-07, 
    4.500845e-07, 4.500845e-07, 4.500845e-07 ;

 RETRANSN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RH2M =
  84.84133, 84.84093, 84.84101, 84.8407, 84.84087, 84.84067, 84.84125, 
    84.84092, 84.84113, 84.84129, 84.84013, 84.84068, 84.83964, 84.83993, 
    84.83878, 84.83968, 84.83869, 84.8388, 84.83849, 84.83858, 84.8382, 
    84.83846, 84.83801, 84.83826, 84.83823, 84.83846, 84.84057, 84.8402, 
    84.84059, 84.84054, 84.84056, 84.84087, 84.84103, 84.84136, 84.8413, 
    84.84106, 84.84052, 84.84069, 84.84025, 84.84026, 84.83982, 84.84, 
    84.83891, 84.83952, 84.83857, 84.8387, 84.83858, 84.83862, 84.83858, 
    84.83876, 84.83868, 84.83885, 84.83997, 84.83976, 84.84045, 84.84092, 
    84.84124, 84.84147, 84.84144, 84.84138, 84.84105, 84.84075, 84.84054, 
    84.84039, 84.84026, 84.83988, 84.8397, 84.83887, 84.83894, 84.83882, 
    84.83871, 84.83853, 84.83856, 84.83849, 84.83882, 84.83859, 84.83897, 
    84.83887, 84.84023, 84.84064, 84.84084, 84.841, 84.84142, 84.84113, 
    84.84124, 84.84097, 84.8408, 84.84088, 84.84039, 84.84058, 84.83969, 
    84.84004, 84.83872, 84.83892, 84.83868, 84.8388, 84.83859, 84.83878, 
    84.83846, 84.83839, 84.83843, 84.83825, 84.83879, 84.83858, 84.84089, 
    84.84087, 84.84081, 84.84109, 84.8411, 84.84136, 84.84113, 84.84103, 
    84.84079, 84.84064, 84.84052, 84.84024, 84.83996, 84.83959, 84.83891, 
    84.83875, 84.83884, 84.83876, 84.83886, 84.83891, 84.83841, 84.83868, 
    84.83828, 84.8383, 84.83848, 84.83829, 84.84086, 84.84094, 84.84122, 
    84.841, 84.84139, 84.84117, 84.84105, 84.84058, 84.84048, 84.84039, 
    84.84021, 84.84, 84.83966, 84.83894, 84.83871, 84.83872, 84.83871, 
    84.83866, 84.8388, 84.83864, 84.83862, 84.83868, 84.8383, 84.83841, 
    84.8383, 84.83837, 84.84091, 84.84078, 84.84085, 84.84072, 84.84082, 
    84.84042, 84.84031, 84.83981, 84.84, 84.83971, 84.83997, 84.83992, 
    84.8397, 84.83995, 84.83897, 84.83978, 84.83866, 84.83945, 84.83864, 
    84.83871, 84.83859, 84.8385, 84.83838, 84.83817, 84.83821, 84.83804, 
    84.84059, 84.84044, 84.84045, 84.84029, 84.84017, 84.83993, 84.83958, 
    84.83971, 84.83948, 84.83899, 84.83979, 84.83957, 84.84033, 84.84019, 
    84.84028, 84.84058, 84.83968, 84.84011, 84.83891, 84.83956, 84.83852, 
    84.83881, 84.83824, 84.83801, 84.83781, 84.83757, 84.84035, 84.84045, 
    84.84027, 84.84002, 84.83981, 84.83955, 84.83952, 84.83947, 84.83891, 
    84.83881, 84.83945, 84.83878, 84.84017, 84.83965, 84.8405, 84.84022, 
    84.84003, 84.84011, 84.83972, 84.83964, 84.83887, 84.83948, 84.83807, 
    84.83848, 84.83739, 84.83768, 84.84049, 84.84035, 84.83989, 84.8401, 
    84.83953, 84.83896, 84.83885, 84.83872, 84.83871, 84.83863, 84.83875, 
    84.83863, 84.83955, 84.83889, 84.83994, 84.83978, 84.83985, 84.83993, 
    84.83969, 84.83945, 84.83945, 84.83893, 84.83873, 84.83952, 84.83802, 
    84.83866, 84.84019, 84.83994, 84.83991, 84.84, 84.83897, 84.83961, 
    84.83863, 84.83878, 84.83854, 84.83865, 84.83868, 84.83882, 84.83892, 
    84.83961, 84.83982, 84.83999, 84.83995, 84.83976, 84.83944, 84.83871, 
    84.83877, 84.83855, 84.83957, 84.83888, 84.83897, 84.83874, 84.83971, 
    84.83882, 84.83984, 84.83978, 84.83962, 84.83887, 84.8388, 84.83873, 
    84.83877, 84.83899, 84.83947, 84.83962, 84.83967, 84.8398, 84.8399, 
    84.83981, 84.83971, 84.83899, 84.83875, 84.8385, 84.83844, 84.83816, 
    84.83839, 84.83802, 84.83833, 84.83779, 84.83879, 84.83834, 84.83961, 
    84.83952, 84.83891, 84.83854, 84.83874, 84.83851, 84.83947, 84.83976, 
    84.83983, 84.83998, 84.83983, 84.83984, 84.8397, 84.83974, 84.83898, 
    84.83959, 84.83868, 84.83851, 84.83806, 84.83779, 84.83754, 84.83743, 
    84.83739, 84.83738 ;

 RH2M_R =
  84.84133, 84.84093, 84.84101, 84.8407, 84.84087, 84.84067, 84.84125, 
    84.84092, 84.84113, 84.84129, 84.84013, 84.84068, 84.83964, 84.83993, 
    84.83878, 84.83968, 84.83869, 84.8388, 84.83849, 84.83858, 84.8382, 
    84.83846, 84.83801, 84.83826, 84.83823, 84.83846, 84.84057, 84.8402, 
    84.84059, 84.84054, 84.84056, 84.84087, 84.84103, 84.84136, 84.8413, 
    84.84106, 84.84052, 84.84069, 84.84025, 84.84026, 84.83982, 84.84, 
    84.83891, 84.83952, 84.83857, 84.8387, 84.83858, 84.83862, 84.83858, 
    84.83876, 84.83868, 84.83885, 84.83997, 84.83976, 84.84045, 84.84092, 
    84.84124, 84.84147, 84.84144, 84.84138, 84.84105, 84.84075, 84.84054, 
    84.84039, 84.84026, 84.83988, 84.8397, 84.83887, 84.83894, 84.83882, 
    84.83871, 84.83853, 84.83856, 84.83849, 84.83882, 84.83859, 84.83897, 
    84.83887, 84.84023, 84.84064, 84.84084, 84.841, 84.84142, 84.84113, 
    84.84124, 84.84097, 84.8408, 84.84088, 84.84039, 84.84058, 84.83969, 
    84.84004, 84.83872, 84.83892, 84.83868, 84.8388, 84.83859, 84.83878, 
    84.83846, 84.83839, 84.83843, 84.83825, 84.83879, 84.83858, 84.84089, 
    84.84087, 84.84081, 84.84109, 84.8411, 84.84136, 84.84113, 84.84103, 
    84.84079, 84.84064, 84.84052, 84.84024, 84.83996, 84.83959, 84.83891, 
    84.83875, 84.83884, 84.83876, 84.83886, 84.83891, 84.83841, 84.83868, 
    84.83828, 84.8383, 84.83848, 84.83829, 84.84086, 84.84094, 84.84122, 
    84.841, 84.84139, 84.84117, 84.84105, 84.84058, 84.84048, 84.84039, 
    84.84021, 84.84, 84.83966, 84.83894, 84.83871, 84.83872, 84.83871, 
    84.83866, 84.8388, 84.83864, 84.83862, 84.83868, 84.8383, 84.83841, 
    84.8383, 84.83837, 84.84091, 84.84078, 84.84085, 84.84072, 84.84082, 
    84.84042, 84.84031, 84.83981, 84.84, 84.83971, 84.83997, 84.83992, 
    84.8397, 84.83995, 84.83897, 84.83978, 84.83866, 84.83945, 84.83864, 
    84.83871, 84.83859, 84.8385, 84.83838, 84.83817, 84.83821, 84.83804, 
    84.84059, 84.84044, 84.84045, 84.84029, 84.84017, 84.83993, 84.83958, 
    84.83971, 84.83948, 84.83899, 84.83979, 84.83957, 84.84033, 84.84019, 
    84.84028, 84.84058, 84.83968, 84.84011, 84.83891, 84.83956, 84.83852, 
    84.83881, 84.83824, 84.83801, 84.83781, 84.83757, 84.84035, 84.84045, 
    84.84027, 84.84002, 84.83981, 84.83955, 84.83952, 84.83947, 84.83891, 
    84.83881, 84.83945, 84.83878, 84.84017, 84.83965, 84.8405, 84.84022, 
    84.84003, 84.84011, 84.83972, 84.83964, 84.83887, 84.83948, 84.83807, 
    84.83848, 84.83739, 84.83768, 84.84049, 84.84035, 84.83989, 84.8401, 
    84.83953, 84.83896, 84.83885, 84.83872, 84.83871, 84.83863, 84.83875, 
    84.83863, 84.83955, 84.83889, 84.83994, 84.83978, 84.83985, 84.83993, 
    84.83969, 84.83945, 84.83945, 84.83893, 84.83873, 84.83952, 84.83802, 
    84.83866, 84.84019, 84.83994, 84.83991, 84.84, 84.83897, 84.83961, 
    84.83863, 84.83878, 84.83854, 84.83865, 84.83868, 84.83882, 84.83892, 
    84.83961, 84.83982, 84.83999, 84.83995, 84.83976, 84.83944, 84.83871, 
    84.83877, 84.83855, 84.83957, 84.83888, 84.83897, 84.83874, 84.83971, 
    84.83882, 84.83984, 84.83978, 84.83962, 84.83887, 84.8388, 84.83873, 
    84.83877, 84.83899, 84.83947, 84.83962, 84.83967, 84.8398, 84.8399, 
    84.83981, 84.83971, 84.83899, 84.83875, 84.8385, 84.83844, 84.83816, 
    84.83839, 84.83802, 84.83833, 84.83779, 84.83879, 84.83834, 84.83961, 
    84.83952, 84.83891, 84.83854, 84.83874, 84.83851, 84.83947, 84.83976, 
    84.83983, 84.83998, 84.83983, 84.83984, 84.8397, 84.83974, 84.83898, 
    84.83959, 84.83868, 84.83851, 84.83806, 84.83779, 84.83754, 84.83743, 
    84.83739, 84.83738 ;

 RH2M_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 RR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABG_PEN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN =
  0.0004638631, 0.0004658033, 0.000465426, 0.0004669909, 0.0004661227, 
    0.0004671474, 0.0004642561, 0.0004658801, 0.0004648432, 0.0004640371, 
    0.0004700274, 0.0004670603, 0.0004731078, 0.0004712159, 0.0004759673, 
    0.0004728134, 0.0004766031, 0.0004758759, 0.0004780634, 0.0004774367, 
    0.0004802349, 0.0004783525, 0.0004816847, 0.0004797851, 0.0004800823, 
    0.0004782902, 0.0004676576, 0.0004696585, 0.000467539, 0.0004678243, 
    0.0004676961, 0.0004661405, 0.0004653566, 0.0004637141, 0.0004640122, 
    0.0004652184, 0.0004679522, 0.000467024, 0.0004693625, 0.0004693097, 
    0.0004719128, 0.0004707391, 0.0004751138, 0.0004738704, 0.0004774628, 
    0.0004765594, 0.0004774203, 0.0004771591, 0.0004774235, 0.0004760986, 
    0.0004766662, 0.0004755002, 0.0004709597, 0.0004722946, 0.0004683127, 
    0.0004659183, 0.0004643271, 0.0004631982, 0.0004633577, 0.000463662, 
    0.0004652253, 0.0004666949, 0.0004678148, 0.0004685639, 0.0004693019, 
    0.0004715365, 0.0004727185, 0.0004753652, 0.0004748873, 0.0004756966, 
    0.0004764694, 0.0004777671, 0.0004775534, 0.0004781251, 0.0004756748, 
    0.0004773033, 0.0004746147, 0.0004753501, 0.000469504, 0.0004672746, 
    0.0004663276, 0.000465498, 0.0004634803, 0.0004648738, 0.0004643244, 
    0.0004656308, 0.0004664611, 0.0004660503, 0.0004685843, 0.0004675991, 
    0.0004727884, 0.0004705534, 0.0004763794, 0.0004749853, 0.0004767133, 
    0.0004758314, 0.0004773423, 0.0004759825, 0.0004783377, 0.0004788507, 
    0.0004785, 0.0004798461, 0.0004759067, 0.0004774198, 0.0004660392, 
    0.0004661062, 0.0004664181, 0.0004650467, 0.0004649627, 0.0004637056, 
    0.000464824, 0.0004653003, 0.000466509, 0.000467224, 0.0004679036, 
    0.0004693979, 0.0004710667, 0.0004733998, 0.0004750756, 0.0004761988, 
    0.0004755099, 0.000476118, 0.0004754382, 0.0004751194, 0.0004786584, 
    0.0004766713, 0.0004796524, 0.0004794874, 0.0004781383, 0.0004795058, 
    0.0004661531, 0.0004657676, 0.0004644296, 0.0004654766, 0.0004635686, 
    0.0004646367, 0.0004652508, 0.0004676198, 0.00046814, 0.0004686227, 
    0.0004695757, 0.0004707988, 0.0004729443, 0.0004748106, 0.0004765141, 
    0.0004763892, 0.0004764331, 0.0004768136, 0.0004758709, 0.0004769683, 
    0.0004771525, 0.0004766708, 0.0004794651, 0.0004786669, 0.0004794837, 
    0.0004789638, 0.0004658928, 0.0004665412, 0.0004661907, 0.0004668497, 
    0.0004663854, 0.0004684495, 0.0004690682, 0.0004719631, 0.0004707747, 
    0.0004726656, 0.0004709666, 0.0004712677, 0.0004727274, 0.0004710582, 
    0.0004747077, 0.0004722338, 0.0004768284, 0.0004743586, 0.000476983, 
    0.0004765063, 0.0004772953, 0.0004780022, 0.000478891, 0.0004805316, 
    0.0004801515, 0.0004815233, 0.0004675077, 0.0004683487, 0.0004682745, 
    0.0004691545, 0.0004698053, 0.0004712158, 0.0004734778, 0.000472627, 
    0.0004741884, 0.0004745019, 0.0004721294, 0.0004735862, 0.0004689109, 
    0.0004696664, 0.0004692164, 0.0004675733, 0.0004728228, 0.0004701289, 
    0.0004751026, 0.0004736435, 0.0004779013, 0.000475784, 0.0004799424, 
    0.0004817202, 0.0004833924, 0.0004853473, 0.0004688075, 0.000468236, 
    0.000469259, 0.0004706747, 0.0004719875, 0.0004737332, 0.0004739116, 
    0.0004742386, 0.0004750854, 0.0004757976, 0.000474342, 0.0004759759, 
    0.0004698419, 0.0004730565, 0.0004680193, 0.0004695365, 0.0004705904, 
    0.0004701279, 0.000472529, 0.0004730949, 0.0004753944, 0.0004742056, 
    0.0004812815, 0.0004781513, 0.0004868349, 0.0004844088, 0.0004680363, 
    0.0004688053, 0.0004714818, 0.0004702083, 0.0004738494, 0.0004747457, 
    0.000475474, 0.0004764053, 0.0004765057, 0.0004770574, 0.0004761532, 
    0.0004770216, 0.0004737363, 0.0004752044, 0.000471175, 0.0004721558, 
    0.0004717045, 0.0004712095, 0.0004727369, 0.0004743643, 0.0004743988, 
    0.0004749205, 0.0004763914, 0.0004738632, 0.0004816857, 0.0004768555, 
    0.0004696438, 0.0004711252, 0.0004713364, 0.0004707626, 0.0004746557, 
    0.0004732452, 0.0004770439, 0.0004760172, 0.0004776992, 0.0004768634, 
    0.0004767403, 0.0004756667, 0.0004749983, 0.0004733095, 0.0004719351, 
    0.0004708451, 0.0004710985, 0.0004722957, 0.0004744636, 0.0004765142, 
    0.000476065, 0.0004775707, 0.0004735843, 0.0004752561, 0.0004746099, 
    0.0004762943, 0.0004726042, 0.0004757484, 0.0004718005, 0.0004721465, 
    0.000473217, 0.0004753705, 0.0004758464, 0.0004763551, 0.000476041, 
    0.000474519, 0.0004742695, 0.0004731906, 0.0004728928, 0.0004720706, 
    0.0004713899, 0.0004720118, 0.0004726648, 0.0004745191, 0.0004761901, 
    0.0004780116, 0.0004784572, 0.0004805858, 0.0004788533, 0.0004817123, 
    0.0004792821, 0.0004834884, 0.0004759301, 0.0004792112, 0.0004732657, 
    0.0004739062, 0.0004750649, 0.0004777218, 0.0004762871, 0.0004779648, 
    0.0004742597, 0.0004723373, 0.0004718395, 0.0004709114, 0.0004718606, 
    0.0004717834, 0.0004726917, 0.0004723997, 0.0004745805, 0.0004734091, 
    0.0004767365, 0.0004779508, 0.0004813789, 0.0004834803, 0.0004856186, 
    0.0004865626, 0.00048685, 0.00048697 ;

 SMINN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_PLANT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_SOIL1N_L1 =
  3.27577e-14, 3.284635e-14, 3.282913e-14, 3.290056e-14, 3.286095e-14, 
    3.290771e-14, 3.277569e-14, 3.284986e-14, 3.280253e-14, 3.27657e-14, 
    3.303898e-14, 3.290375e-14, 3.317934e-14, 3.309325e-14, 3.330937e-14, 
    3.316593e-14, 3.333827e-14, 3.330526e-14, 3.340464e-14, 3.337618e-14, 
    3.350309e-14, 3.341777e-14, 3.356885e-14, 3.348274e-14, 3.349621e-14, 
    3.341495e-14, 3.293101e-14, 3.302215e-14, 3.29256e-14, 3.29386e-14, 
    3.293278e-14, 3.286176e-14, 3.282594e-14, 3.275094e-14, 3.276457e-14, 
    3.281966e-14, 3.294445e-14, 3.290213e-14, 3.300881e-14, 3.30064e-14, 
    3.3125e-14, 3.307155e-14, 3.327063e-14, 3.321411e-14, 3.337737e-14, 
    3.333634e-14, 3.337544e-14, 3.336359e-14, 3.33756e-14, 3.33154e-14, 
    3.33412e-14, 3.328822e-14, 3.308156e-14, 3.314234e-14, 3.29609e-14, 
    3.285157e-14, 3.277894e-14, 3.272735e-14, 3.273465e-14, 3.274854e-14, 
    3.281998e-14, 3.288711e-14, 3.293822e-14, 3.29724e-14, 3.300606e-14, 
    3.310779e-14, 3.316164e-14, 3.328204e-14, 3.326034e-14, 3.329711e-14, 
    3.333225e-14, 3.339119e-14, 3.338149e-14, 3.340744e-14, 3.329616e-14, 
    3.337013e-14, 3.324798e-14, 3.32814e-14, 3.301511e-14, 3.291355e-14, 
    3.287027e-14, 3.283243e-14, 3.274025e-14, 3.280392e-14, 3.277882e-14, 
    3.283853e-14, 3.287644e-14, 3.28577e-14, 3.297333e-14, 3.292839e-14, 
    3.316483e-14, 3.306307e-14, 3.332815e-14, 3.32648e-14, 3.334334e-14, 
    3.330328e-14, 3.33719e-14, 3.331014e-14, 3.341711e-14, 3.344037e-14, 
    3.342447e-14, 3.348556e-14, 3.330671e-14, 3.337543e-14, 3.285717e-14, 
    3.286022e-14, 3.287447e-14, 3.281182e-14, 3.280799e-14, 3.275056e-14, 
    3.280167e-14, 3.282342e-14, 3.287864e-14, 3.291127e-14, 3.294228e-14, 
    3.301043e-14, 3.308646e-14, 3.319268e-14, 3.326891e-14, 3.331997e-14, 
    3.328867e-14, 3.331631e-14, 3.328541e-14, 3.327093e-14, 3.343165e-14, 
    3.334143e-14, 3.347677e-14, 3.346929e-14, 3.340806e-14, 3.347014e-14, 
    3.286237e-14, 3.284478e-14, 3.278364e-14, 3.283149e-14, 3.274431e-14, 
    3.279311e-14, 3.282115e-14, 3.292931e-14, 3.295308e-14, 3.297508e-14, 
    3.301855e-14, 3.307429e-14, 3.317196e-14, 3.325685e-14, 3.33343e-14, 
    3.332863e-14, 3.333063e-14, 3.334791e-14, 3.330508e-14, 3.335494e-14, 
    3.33633e-14, 3.334143e-14, 3.346829e-14, 3.343207e-14, 3.346913e-14, 
    3.344555e-14, 3.28505e-14, 3.28801e-14, 3.286411e-14, 3.289418e-14, 
    3.287298e-14, 3.296715e-14, 3.299536e-14, 3.312727e-14, 3.307318e-14, 
    3.315927e-14, 3.308194e-14, 3.309564e-14, 3.316203e-14, 3.308613e-14, 
    3.325216e-14, 3.31396e-14, 3.334858e-14, 3.323627e-14, 3.335561e-14, 
    3.333397e-14, 3.336981e-14, 3.340189e-14, 3.344225e-14, 3.351663e-14, 
    3.349942e-14, 3.35616e-14, 3.292422e-14, 3.296257e-14, 3.295921e-14, 
    3.299934e-14, 3.3029e-14, 3.309328e-14, 3.319625e-14, 3.315755e-14, 
    3.32286e-14, 3.324283e-14, 3.313491e-14, 3.320118e-14, 3.298824e-14, 
    3.302266e-14, 3.300218e-14, 3.292723e-14, 3.316644e-14, 3.304375e-14, 
    3.327016e-14, 3.320383e-14, 3.339732e-14, 3.330112e-14, 3.348994e-14, 
    3.357047e-14, 3.364628e-14, 3.373468e-14, 3.298351e-14, 3.295746e-14, 
    3.300412e-14, 3.30686e-14, 3.312842e-14, 3.320787e-14, 3.321601e-14, 
    3.323087e-14, 3.326938e-14, 3.330175e-14, 3.323556e-14, 3.330986e-14, 
    3.303061e-14, 3.317709e-14, 3.294759e-14, 3.301674e-14, 3.306481e-14, 
    3.304374e-14, 3.315313e-14, 3.317888e-14, 3.328343e-14, 3.322942e-14, 
    3.355059e-14, 3.340864e-14, 3.380198e-14, 3.369224e-14, 3.294835e-14, 
    3.298343e-14, 3.310538e-14, 3.304738e-14, 3.321319e-14, 3.325392e-14, 
    3.328705e-14, 3.332935e-14, 3.333393e-14, 3.335898e-14, 3.331792e-14, 
    3.335737e-14, 3.320804e-14, 3.32748e-14, 3.309147e-14, 3.313612e-14, 
    3.311559e-14, 3.309305e-14, 3.31626e-14, 3.32366e-14, 3.323821e-14, 
    3.32619e-14, 3.332862e-14, 3.321386e-14, 3.356883e-14, 3.334973e-14, 
    3.302166e-14, 3.308912e-14, 3.309879e-14, 3.307266e-14, 3.324983e-14, 
    3.318569e-14, 3.335838e-14, 3.331174e-14, 3.338814e-14, 3.335018e-14, 
    3.33446e-14, 3.329582e-14, 3.326543e-14, 3.318862e-14, 3.312608e-14, 
    3.307645e-14, 3.3088e-14, 3.31425e-14, 3.324113e-14, 3.333433e-14, 
    3.331391e-14, 3.338234e-14, 3.320117e-14, 3.327716e-14, 3.324778e-14, 
    3.332437e-14, 3.315651e-14, 3.329938e-14, 3.311994e-14, 3.31357e-14, 
    3.318441e-14, 3.32823e-14, 3.330398e-14, 3.332708e-14, 3.331283e-14, 
    3.324362e-14, 3.32323e-14, 3.318324e-14, 3.316967e-14, 3.313227e-14, 
    3.310128e-14, 3.312959e-14, 3.31593e-14, 3.324366e-14, 3.331961e-14, 
    3.340234e-14, 3.342259e-14, 3.351905e-14, 3.344049e-14, 3.357005e-14, 
    3.345985e-14, 3.365054e-14, 3.33077e-14, 3.345667e-14, 3.318664e-14, 
    3.321578e-14, 3.326842e-14, 3.338912e-14, 3.332401e-14, 3.340017e-14, 
    3.323186e-14, 3.314436e-14, 3.312174e-14, 3.307947e-14, 3.312271e-14, 
    3.311919e-14, 3.316055e-14, 3.314727e-14, 3.324646e-14, 3.31932e-14, 
    3.334445e-14, 3.339957e-14, 3.355508e-14, 3.365024e-14, 3.374704e-14, 
    3.378972e-14, 3.380271e-14, 3.380813e-14 ;

 SMINN_TO_SOIL1N_L2 =
  1.089232e-14, 1.092182e-14, 1.091609e-14, 1.093987e-14, 1.092668e-14, 
    1.094225e-14, 1.089831e-14, 1.092299e-14, 1.090724e-14, 1.089498e-14, 
    1.098594e-14, 1.094093e-14, 1.103266e-14, 1.1004e-14, 1.107594e-14, 
    1.10282e-14, 1.108556e-14, 1.107457e-14, 1.110765e-14, 1.109818e-14, 
    1.114042e-14, 1.111202e-14, 1.116231e-14, 1.113365e-14, 1.113813e-14, 
    1.111108e-14, 1.095e-14, 1.098034e-14, 1.09482e-14, 1.095253e-14, 
    1.095059e-14, 1.092695e-14, 1.091503e-14, 1.089007e-14, 1.08946e-14, 
    1.091294e-14, 1.095448e-14, 1.094039e-14, 1.09759e-14, 1.09751e-14, 
    1.101457e-14, 1.099678e-14, 1.106304e-14, 1.104423e-14, 1.109858e-14, 
    1.108492e-14, 1.109793e-14, 1.109399e-14, 1.109798e-14, 1.107795e-14, 
    1.108653e-14, 1.10689e-14, 1.100011e-14, 1.102034e-14, 1.095995e-14, 
    1.092356e-14, 1.089939e-14, 1.088221e-14, 1.088464e-14, 1.088927e-14, 
    1.091305e-14, 1.093539e-14, 1.09524e-14, 1.096378e-14, 1.097498e-14, 
    1.100884e-14, 1.102677e-14, 1.106684e-14, 1.105962e-14, 1.107186e-14, 
    1.108356e-14, 1.110317e-14, 1.109995e-14, 1.110858e-14, 1.107154e-14, 
    1.109616e-14, 1.105551e-14, 1.106663e-14, 1.0978e-14, 1.094419e-14, 
    1.092978e-14, 1.091719e-14, 1.088651e-14, 1.09077e-14, 1.089935e-14, 
    1.091922e-14, 1.093184e-14, 1.09256e-14, 1.096409e-14, 1.094913e-14, 
    1.102783e-14, 1.099396e-14, 1.108219e-14, 1.106111e-14, 1.108725e-14, 
    1.107391e-14, 1.109675e-14, 1.10762e-14, 1.11118e-14, 1.111954e-14, 
    1.111425e-14, 1.113459e-14, 1.107506e-14, 1.109793e-14, 1.092542e-14, 
    1.092644e-14, 1.093118e-14, 1.091033e-14, 1.090906e-14, 1.088994e-14, 
    1.090695e-14, 1.091419e-14, 1.093257e-14, 1.094343e-14, 1.095375e-14, 
    1.097644e-14, 1.100174e-14, 1.10371e-14, 1.106247e-14, 1.107947e-14, 
    1.106905e-14, 1.107825e-14, 1.106796e-14, 1.106314e-14, 1.111664e-14, 
    1.108661e-14, 1.113166e-14, 1.112917e-14, 1.110879e-14, 1.112945e-14, 
    1.092716e-14, 1.09213e-14, 1.090095e-14, 1.091688e-14, 1.088786e-14, 
    1.09041e-14, 1.091343e-14, 1.094944e-14, 1.095735e-14, 1.096467e-14, 
    1.097914e-14, 1.099769e-14, 1.10302e-14, 1.105846e-14, 1.108424e-14, 
    1.108235e-14, 1.108302e-14, 1.108877e-14, 1.107451e-14, 1.109111e-14, 
    1.109389e-14, 1.108661e-14, 1.112884e-14, 1.111678e-14, 1.112912e-14, 
    1.112127e-14, 1.09232e-14, 1.093306e-14, 1.092773e-14, 1.093774e-14, 
    1.093069e-14, 1.096203e-14, 1.097142e-14, 1.101533e-14, 1.099732e-14, 
    1.102598e-14, 1.100024e-14, 1.10048e-14, 1.10269e-14, 1.100163e-14, 
    1.10569e-14, 1.101943e-14, 1.108899e-14, 1.105161e-14, 1.109133e-14, 
    1.108413e-14, 1.109606e-14, 1.110674e-14, 1.112017e-14, 1.114493e-14, 
    1.11392e-14, 1.11599e-14, 1.094774e-14, 1.096051e-14, 1.095939e-14, 
    1.097275e-14, 1.098262e-14, 1.100401e-14, 1.103829e-14, 1.102541e-14, 
    1.104906e-14, 1.105379e-14, 1.101787e-14, 1.103993e-14, 1.096905e-14, 
    1.098051e-14, 1.097369e-14, 1.094875e-14, 1.102837e-14, 1.098753e-14, 
    1.106289e-14, 1.104081e-14, 1.110521e-14, 1.107319e-14, 1.113604e-14, 
    1.116285e-14, 1.118808e-14, 1.121751e-14, 1.096748e-14, 1.095881e-14, 
    1.097434e-14, 1.09958e-14, 1.101571e-14, 1.104216e-14, 1.104486e-14, 
    1.104981e-14, 1.106263e-14, 1.10734e-14, 1.105137e-14, 1.10761e-14, 
    1.098315e-14, 1.103191e-14, 1.095552e-14, 1.097854e-14, 1.099454e-14, 
    1.098753e-14, 1.102393e-14, 1.103251e-14, 1.106731e-14, 1.104933e-14, 
    1.115623e-14, 1.110898e-14, 1.123991e-14, 1.120338e-14, 1.095577e-14, 
    1.096745e-14, 1.100804e-14, 1.098874e-14, 1.104392e-14, 1.105748e-14, 
    1.106851e-14, 1.108259e-14, 1.108411e-14, 1.109245e-14, 1.107879e-14, 
    1.109192e-14, 1.104221e-14, 1.106443e-14, 1.100341e-14, 1.101827e-14, 
    1.101144e-14, 1.100394e-14, 1.102709e-14, 1.105172e-14, 1.105225e-14, 
    1.106014e-14, 1.108235e-14, 1.104415e-14, 1.116231e-14, 1.108937e-14, 
    1.098018e-14, 1.100263e-14, 1.100585e-14, 1.099715e-14, 1.105612e-14, 
    1.103477e-14, 1.109225e-14, 1.107673e-14, 1.110216e-14, 1.108953e-14, 
    1.108767e-14, 1.107143e-14, 1.106132e-14, 1.103575e-14, 1.101493e-14, 
    1.099841e-14, 1.100226e-14, 1.10204e-14, 1.105323e-14, 1.108425e-14, 
    1.107745e-14, 1.110023e-14, 1.103993e-14, 1.106522e-14, 1.105544e-14, 
    1.108093e-14, 1.102506e-14, 1.107262e-14, 1.101289e-14, 1.101813e-14, 
    1.103435e-14, 1.106693e-14, 1.107415e-14, 1.108183e-14, 1.107709e-14, 
    1.105405e-14, 1.105029e-14, 1.103396e-14, 1.102944e-14, 1.101699e-14, 
    1.100667e-14, 1.10161e-14, 1.102599e-14, 1.105407e-14, 1.107935e-14, 
    1.110689e-14, 1.111363e-14, 1.114573e-14, 1.111959e-14, 1.116271e-14, 
    1.112603e-14, 1.11895e-14, 1.107538e-14, 1.112497e-14, 1.103509e-14, 
    1.104479e-14, 1.106231e-14, 1.110249e-14, 1.108081e-14, 1.110616e-14, 
    1.105014e-14, 1.102102e-14, 1.101349e-14, 1.099942e-14, 1.101381e-14, 
    1.101264e-14, 1.10264e-14, 1.102198e-14, 1.1055e-14, 1.103727e-14, 
    1.108762e-14, 1.110596e-14, 1.115773e-14, 1.11894e-14, 1.122162e-14, 
    1.123583e-14, 1.124015e-14, 1.124196e-14 ;

 SMINN_TO_SOIL1N_S2 =
  -8.366578e-11, -8.403394e-11, -8.396236e-11, -8.425931e-11, -8.409459e-11, 
    -8.428903e-11, -8.374042e-11, -8.404856e-11, -8.385185e-11, 
    -8.369892e-11, -8.483559e-11, -8.427255e-11, -8.542037e-11, 
    -8.506131e-11, -8.596328e-11, -8.536451e-11, -8.608401e-11, 
    -8.594599e-11, -8.636136e-11, -8.624237e-11, -8.677367e-11, 
    -8.641628e-11, -8.704908e-11, -8.668832e-11, -8.674476e-11, 
    -8.640449e-11, -8.438585e-11, -8.476549e-11, -8.436336e-11, -8.44175e-11, 
    -8.439321e-11, -8.409799e-11, -8.394923e-11, -8.363764e-11, -8.36942e-11, 
    -8.392306e-11, -8.444184e-11, -8.426573e-11, -8.470955e-11, 
    -8.469953e-11, -8.519363e-11, -8.497086e-11, -8.580131e-11, 
    -8.556528e-11, -8.624734e-11, -8.607581e-11, -8.623928e-11, 
    -8.618971e-11, -8.623992e-11, -8.598836e-11, -8.609614e-11, 
    -8.587477e-11, -8.501258e-11, -8.526598e-11, -8.451022e-11, -8.40558e-11, 
    -8.375393e-11, -8.353974e-11, -8.357002e-11, -8.362775e-11, -8.39244e-11, 
    -8.420329e-11, -8.441583e-11, -8.455801e-11, -8.469809e-11, 
    -8.512214e-11, -8.534655e-11, -8.584904e-11, -8.575835e-11, 
    -8.591199e-11, -8.605874e-11, -8.630515e-11, -8.626459e-11, 
    -8.637315e-11, -8.590792e-11, -8.621712e-11, -8.570669e-11, -8.58463e-11, 
    -8.473621e-11, -8.431324e-11, -8.413349e-11, -8.397612e-11, 
    -8.359331e-11, -8.385768e-11, -8.375346e-11, -8.400139e-11, 
    -8.415893e-11, -8.408101e-11, -8.456189e-11, -8.437494e-11, 
    -8.535985e-11, -8.493562e-11, -8.604163e-11, -8.577696e-11, 
    -8.610506e-11, -8.593764e-11, -8.622451e-11, -8.596632e-11, 
    -8.641355e-11, -8.651094e-11, -8.644439e-11, -8.670002e-11, 
    -8.595202e-11, -8.623928e-11, -8.407883e-11, -8.409154e-11, 
    -8.415073e-11, -8.389051e-11, -8.387458e-11, -8.363609e-11, -8.38483e-11, 
    -8.393867e-11, -8.416806e-11, -8.430375e-11, -8.443274e-11, 
    -8.471634e-11, -8.503307e-11, -8.547595e-11, -8.579412e-11, -8.60074e-11, 
    -8.587662e-11, -8.599208e-11, -8.5863e-11, -8.580251e-11, -8.647445e-11, 
    -8.609715e-11, -8.666325e-11, -8.663192e-11, -8.637573e-11, 
    -8.663546e-11, -8.410046e-11, -8.402733e-11, -8.377344e-11, 
    -8.397213e-11, -8.361012e-11, -8.381276e-11, -8.392928e-11, 
    -8.437886e-11, -8.447762e-11, -8.456921e-11, -8.475011e-11, 
    -8.498226e-11, -8.53895e-11, -8.574383e-11, -8.606728e-11, -8.604358e-11, 
    -8.605192e-11, -8.612418e-11, -8.59452e-11, -8.615357e-11, -8.618854e-11, 
    -8.60971e-11, -8.662773e-11, -8.647613e-11, -8.663126e-11, -8.653255e-11, 
    -8.40511e-11, -8.417415e-11, -8.410766e-11, -8.423269e-11, -8.414461e-11, 
    -8.453629e-11, -8.465372e-11, -8.520321e-11, -8.497769e-11, 
    -8.533659e-11, -8.501414e-11, -8.507128e-11, -8.534831e-11, 
    -8.503157e-11, -8.57243e-11, -8.525466e-11, -8.612699e-11, -8.565803e-11, 
    -8.615638e-11, -8.606588e-11, -8.621572e-11, -8.634991e-11, 
    -8.651874e-11, -8.683025e-11, -8.675811e-11, -8.701862e-11, 
    -8.435758e-11, -8.451719e-11, -8.450313e-11, -8.467015e-11, 
    -8.479368e-11, -8.50614e-11, -8.549078e-11, -8.532931e-11, -8.562574e-11, 
    -8.568524e-11, -8.52349e-11, -8.551141e-11, -8.4624e-11, -8.476739e-11, 
    -8.468201e-11, -8.437018e-11, -8.536653e-11, -8.485521e-11, 
    -8.579938e-11, -8.552239e-11, -8.633078e-11, -8.592876e-11, -8.67184e-11, 
    -8.705599e-11, -8.737367e-11, -8.774496e-11, -8.460429e-11, 
    -8.449584e-11, -8.469001e-11, -8.495867e-11, -8.520792e-11, 
    -8.553928e-11, -8.557319e-11, -8.563526e-11, -8.579606e-11, 
    -8.593126e-11, -8.56549e-11, -8.596515e-11, -8.480065e-11, -8.541091e-11, 
    -8.445485e-11, -8.474275e-11, -8.494283e-11, -8.485505e-11, 
    -8.531086e-11, -8.541828e-11, -8.585483e-11, -8.562916e-11, 
    -8.697268e-11, -8.637827e-11, -8.802765e-11, -8.756672e-11, 
    -8.445795e-11, -8.460391e-11, -8.51119e-11, -8.48702e-11, -8.556141e-11, 
    -8.573154e-11, -8.586984e-11, -8.604665e-11, -8.606573e-11, 
    -8.617049e-11, -8.599883e-11, -8.616371e-11, -8.553999e-11, 
    -8.581871e-11, -8.505383e-11, -8.524e-11, -8.515436e-11, -8.506041e-11, 
    -8.535035e-11, -8.565926e-11, -8.566584e-11, -8.57649e-11, -8.604404e-11, 
    -8.55642e-11, -8.704942e-11, -8.613221e-11, -8.476307e-11, -8.504422e-11, 
    -8.508437e-11, -8.497546e-11, -8.571448e-11, -8.544671e-11, 
    -8.616793e-11, -8.597301e-11, -8.629238e-11, -8.613368e-11, 
    -8.611033e-11, -8.59065e-11, -8.57796e-11, -8.545899e-11, -8.519813e-11, 
    -8.499126e-11, -8.503936e-11, -8.52666e-11, -8.567815e-11, -8.606747e-11, 
    -8.598219e-11, -8.626811e-11, -8.551129e-11, -8.582864e-11, 
    -8.570598e-11, -8.60258e-11, -8.532502e-11, -8.592182e-11, -8.517248e-11, 
    -8.523818e-11, -8.54414e-11, -8.585017e-11, -8.594059e-11, -8.603716e-11, 
    -8.597757e-11, -8.568859e-11, -8.564124e-11, -8.543646e-11, 
    -8.537992e-11, -8.522387e-11, -8.509469e-11, -8.521272e-11, 
    -8.533668e-11, -8.568871e-11, -8.600595e-11, -8.635183e-11, 
    -8.643646e-11, -8.684062e-11, -8.651164e-11, -8.705453e-11, -8.6593e-11, 
    -8.739193e-11, -8.595638e-11, -8.65794e-11, -8.545064e-11, -8.557224e-11, 
    -8.579219e-11, -8.629665e-11, -8.60243e-11, -8.634281e-11, -8.563938e-11, 
    -8.527444e-11, -8.518e-11, -8.500383e-11, -8.518403e-11, -8.516938e-11, 
    -8.534181e-11, -8.52864e-11, -8.570039e-11, -8.547801e-11, -8.610975e-11, 
    -8.634029e-11, -8.699132e-11, -8.739044e-11, -8.779668e-11, 
    -8.797604e-11, -8.803062e-11, -8.805345e-11 ;

 SMINN_TO_SOIL1N_S3 =
  -2.016494e-12, -2.025365e-12, -2.02364e-12, -2.030796e-12, -2.026826e-12, 
    -2.031512e-12, -2.018292e-12, -2.025717e-12, -2.020977e-12, 
    -2.017292e-12, -2.044682e-12, -2.031115e-12, -2.058773e-12, 
    -2.050121e-12, -2.071855e-12, -2.057427e-12, -2.074764e-12, 
    -2.071439e-12, -2.081448e-12, -2.07858e-12, -2.091383e-12, -2.082771e-12, 
    -2.098019e-12, -2.089326e-12, -2.090686e-12, -2.082487e-12, 
    -2.033845e-12, -2.042993e-12, -2.033303e-12, -2.034608e-12, 
    -2.034022e-12, -2.026909e-12, -2.023324e-12, -2.015816e-12, 
    -2.017179e-12, -2.022693e-12, -2.035194e-12, -2.03095e-12, -2.041645e-12, 
    -2.041404e-12, -2.05331e-12, -2.047941e-12, -2.067952e-12, -2.062265e-12, 
    -2.0787e-12, -2.074567e-12, -2.078506e-12, -2.077311e-12, -2.078521e-12, 
    -2.07246e-12, -2.075057e-12, -2.069723e-12, -2.048947e-12, -2.055053e-12, 
    -2.036842e-12, -2.025892e-12, -2.018618e-12, -2.013457e-12, 
    -2.014186e-12, -2.015577e-12, -2.022726e-12, -2.029446e-12, 
    -2.034567e-12, -2.037993e-12, -2.041369e-12, -2.051587e-12, 
    -2.056994e-12, -2.069102e-12, -2.066917e-12, -2.070619e-12, 
    -2.074156e-12, -2.080093e-12, -2.079116e-12, -2.081731e-12, 
    -2.070521e-12, -2.077972e-12, -2.065673e-12, -2.069036e-12, 
    -2.042287e-12, -2.032095e-12, -2.027764e-12, -2.023972e-12, 
    -2.014747e-12, -2.021118e-12, -2.018607e-12, -2.024581e-12, 
    -2.028377e-12, -2.026499e-12, -2.038087e-12, -2.033582e-12, 
    -2.057315e-12, -2.047093e-12, -2.073743e-12, -2.067366e-12, 
    -2.075272e-12, -2.071237e-12, -2.07815e-12, -2.071929e-12, -2.082705e-12, 
    -2.085052e-12, -2.083448e-12, -2.089608e-12, -2.071584e-12, 
    -2.078506e-12, -2.026447e-12, -2.026753e-12, -2.028179e-12, 
    -2.021909e-12, -2.021525e-12, -2.015778e-12, -2.020892e-12, 
    -2.023069e-12, -2.028597e-12, -2.031867e-12, -2.034975e-12, 
    -2.041809e-12, -2.049441e-12, -2.060112e-12, -2.067779e-12, 
    -2.072918e-12, -2.069767e-12, -2.072549e-12, -2.069439e-12, 
    -2.067981e-12, -2.084172e-12, -2.075081e-12, -2.088722e-12, 
    -2.087967e-12, -2.081794e-12, -2.088052e-12, -2.026968e-12, 
    -2.025206e-12, -2.019088e-12, -2.023876e-12, -2.015153e-12, 
    -2.020035e-12, -2.022843e-12, -2.033676e-12, -2.036056e-12, 
    -2.038263e-12, -2.042622e-12, -2.048216e-12, -2.058029e-12, 
    -2.066567e-12, -2.074361e-12, -2.07379e-12, -2.073991e-12, -2.075732e-12, 
    -2.071419e-12, -2.07644e-12, -2.077283e-12, -2.07508e-12, -2.087866e-12, 
    -2.084213e-12, -2.087951e-12, -2.085573e-12, -2.025779e-12, 
    -2.028744e-12, -2.027141e-12, -2.030154e-12, -2.028032e-12, -2.03747e-12, 
    -2.0403e-12, -2.05354e-12, -2.048106e-12, -2.056754e-12, -2.048984e-12, 
    -2.050361e-12, -2.057037e-12, -2.049404e-12, -2.066097e-12, -2.05478e-12, 
    -2.0758e-12, -2.0645e-12, -2.076508e-12, -2.074327e-12, -2.077938e-12, 
    -2.081172e-12, -2.08524e-12, -2.092746e-12, -2.091008e-12, -2.097285e-12, 
    -2.033164e-12, -2.03701e-12, -2.036671e-12, -2.040696e-12, -2.043672e-12, 
    -2.050123e-12, -2.06047e-12, -2.056579e-12, -2.063722e-12, -2.065156e-12, 
    -2.054304e-12, -2.060967e-12, -2.039584e-12, -2.043038e-12, 
    -2.040981e-12, -2.033467e-12, -2.057476e-12, -2.045155e-12, 
    -2.067906e-12, -2.061231e-12, -2.080711e-12, -2.071023e-12, 
    -2.090051e-12, -2.098185e-12, -2.10584e-12, -2.114787e-12, -2.039108e-12, 
    -2.036495e-12, -2.041174e-12, -2.047648e-12, -2.053654e-12, 
    -2.061639e-12, -2.062455e-12, -2.063951e-12, -2.067826e-12, 
    -2.071084e-12, -2.064425e-12, -2.0719e-12, -2.04384e-12, -2.058545e-12, 
    -2.035508e-12, -2.042445e-12, -2.047266e-12, -2.045151e-12, 
    -2.056134e-12, -2.058723e-12, -2.069242e-12, -2.063804e-12, 
    -2.096178e-12, -2.081855e-12, -2.121598e-12, -2.110492e-12, 
    -2.035582e-12, -2.039099e-12, -2.05134e-12, -2.045516e-12, -2.062171e-12, 
    -2.066271e-12, -2.069604e-12, -2.073864e-12, -2.074324e-12, 
    -2.076848e-12, -2.072712e-12, -2.076685e-12, -2.061656e-12, 
    -2.068372e-12, -2.049941e-12, -2.054427e-12, -2.052363e-12, 
    -2.050099e-12, -2.057086e-12, -2.064529e-12, -2.064688e-12, 
    -2.067075e-12, -2.073801e-12, -2.062239e-12, -2.098027e-12, 
    -2.075926e-12, -2.042935e-12, -2.049709e-12, -2.050677e-12, 
    -2.048052e-12, -2.06586e-12, -2.059408e-12, -2.076787e-12, -2.07209e-12, 
    -2.079785e-12, -2.075961e-12, -2.075399e-12, -2.070487e-12, 
    -2.067429e-12, -2.059704e-12, -2.053418e-12, -2.048433e-12, 
    -2.049592e-12, -2.055068e-12, -2.064985e-12, -2.074366e-12, 
    -2.072311e-12, -2.079201e-12, -2.060964e-12, -2.068611e-12, 
    -2.065655e-12, -2.073362e-12, -2.056476e-12, -2.070856e-12, -2.0528e-12, 
    -2.054383e-12, -2.05928e-12, -2.06913e-12, -2.071309e-12, -2.073636e-12, 
    -2.0722e-12, -2.065236e-12, -2.064095e-12, -2.059161e-12, -2.057798e-12, 
    -2.054038e-12, -2.050925e-12, -2.053769e-12, -2.056756e-12, 
    -2.065239e-12, -2.072884e-12, -2.081218e-12, -2.083257e-12, 
    -2.092996e-12, -2.085068e-12, -2.09815e-12, -2.087029e-12, -2.10628e-12, 
    -2.071689e-12, -2.086701e-12, -2.059503e-12, -2.062433e-12, 
    -2.067733e-12, -2.079888e-12, -2.073326e-12, -2.081001e-12, 
    -2.064051e-12, -2.055257e-12, -2.052981e-12, -2.048736e-12, 
    -2.053078e-12, -2.052725e-12, -2.05688e-12, -2.055545e-12, -2.065521e-12, 
    -2.060162e-12, -2.075385e-12, -2.08094e-12, -2.096627e-12, -2.106244e-12, 
    -2.116033e-12, -2.120355e-12, -2.12167e-12, -2.12222e-12 ;

 SMINN_TO_SOIL2N_L3 =
  3.538413e-15, 3.547998e-15, 3.546136e-15, 3.55386e-15, 3.549577e-15, 
    3.554633e-15, 3.540358e-15, 3.548377e-15, 3.543259e-15, 3.539278e-15, 
    3.568827e-15, 3.554204e-15, 3.584003e-15, 3.574694e-15, 3.598063e-15, 
    3.582553e-15, 3.601189e-15, 3.59762e-15, 3.608365e-15, 3.605288e-15, 
    3.619011e-15, 3.609785e-15, 3.626121e-15, 3.61681e-15, 3.618266e-15, 
    3.609479e-15, 3.557152e-15, 3.567007e-15, 3.556567e-15, 3.557973e-15, 
    3.557343e-15, 3.549664e-15, 3.54579e-15, 3.537682e-15, 3.539155e-15, 
    3.545112e-15, 3.558606e-15, 3.554029e-15, 3.565564e-15, 3.565304e-15, 
    3.578127e-15, 3.572348e-15, 3.593874e-15, 3.587763e-15, 3.605416e-15, 
    3.600979e-15, 3.605208e-15, 3.603926e-15, 3.605224e-15, 3.598716e-15, 
    3.601505e-15, 3.595776e-15, 3.57343e-15, 3.580003e-15, 3.560384e-15, 
    3.548562e-15, 3.540709e-15, 3.535131e-15, 3.53592e-15, 3.537423e-15, 
    3.545146e-15, 3.552405e-15, 3.557932e-15, 3.561627e-15, 3.565267e-15, 
    3.576267e-15, 3.58209e-15, 3.595108e-15, 3.592762e-15, 3.596738e-15, 
    3.600538e-15, 3.60691e-15, 3.605862e-15, 3.608668e-15, 3.596635e-15, 
    3.604633e-15, 3.591425e-15, 3.595039e-15, 3.566245e-15, 3.555265e-15, 
    3.550584e-15, 3.546493e-15, 3.536526e-15, 3.54341e-15, 3.540696e-15, 
    3.547152e-15, 3.551251e-15, 3.549225e-15, 3.561728e-15, 3.556869e-15, 
    3.582435e-15, 3.571432e-15, 3.600095e-15, 3.593244e-15, 3.601736e-15, 
    3.597404e-15, 3.604824e-15, 3.598147e-15, 3.609713e-15, 3.612228e-15, 
    3.610509e-15, 3.617114e-15, 3.597776e-15, 3.605206e-15, 3.549167e-15, 
    3.549498e-15, 3.551038e-15, 3.544264e-15, 3.54385e-15, 3.537641e-15, 
    3.543167e-15, 3.545519e-15, 3.551489e-15, 3.555018e-15, 3.558371e-15, 
    3.565739e-15, 3.57396e-15, 3.585446e-15, 3.593688e-15, 3.59921e-15, 
    3.595825e-15, 3.598813e-15, 3.595472e-15, 3.593907e-15, 3.611285e-15, 
    3.60153e-15, 3.616165e-15, 3.615356e-15, 3.608734e-15, 3.615447e-15, 
    3.54973e-15, 3.547828e-15, 3.541218e-15, 3.546391e-15, 3.536964e-15, 
    3.542241e-15, 3.545273e-15, 3.556968e-15, 3.559538e-15, 3.561917e-15, 
    3.566617e-15, 3.572644e-15, 3.583205e-15, 3.592384e-15, 3.600759e-15, 
    3.600146e-15, 3.600362e-15, 3.602231e-15, 3.597599e-15, 3.602991e-15, 
    3.603894e-15, 3.60153e-15, 3.615248e-15, 3.611331e-15, 3.615339e-15, 
    3.612789e-15, 3.548447e-15, 3.551647e-15, 3.549918e-15, 3.553169e-15, 
    3.550878e-15, 3.561059e-15, 3.56411e-15, 3.578373e-15, 3.572525e-15, 
    3.581833e-15, 3.573471e-15, 3.574953e-15, 3.582132e-15, 3.573924e-15, 
    3.591877e-15, 3.579706e-15, 3.602303e-15, 3.590159e-15, 3.603063e-15, 
    3.600723e-15, 3.604599e-15, 3.608068e-15, 3.612432e-15, 3.620475e-15, 
    3.618613e-15, 3.625337e-15, 3.556418e-15, 3.560564e-15, 3.560201e-15, 
    3.56454e-15, 3.567748e-15, 3.574698e-15, 3.585831e-15, 3.581647e-15, 
    3.58933e-15, 3.590869e-15, 3.579199e-15, 3.586365e-15, 3.56334e-15, 
    3.567062e-15, 3.564847e-15, 3.556743e-15, 3.582609e-15, 3.569343e-15, 
    3.593824e-15, 3.586651e-15, 3.607573e-15, 3.597171e-15, 3.617588e-15, 
    3.626297e-15, 3.634494e-15, 3.644052e-15, 3.562829e-15, 3.560012e-15, 
    3.565057e-15, 3.572029e-15, 3.578498e-15, 3.587088e-15, 3.587968e-15, 
    3.589576e-15, 3.593739e-15, 3.597239e-15, 3.590082e-15, 3.598116e-15, 
    3.567921e-15, 3.58376e-15, 3.558945e-15, 3.566422e-15, 3.571619e-15, 
    3.569341e-15, 3.581169e-15, 3.583954e-15, 3.595258e-15, 3.589419e-15, 
    3.624146e-15, 3.608797e-15, 3.65133e-15, 3.639464e-15, 3.559027e-15, 
    3.56282e-15, 3.576006e-15, 3.569735e-15, 3.587663e-15, 3.592067e-15, 
    3.59565e-15, 3.600224e-15, 3.600719e-15, 3.603428e-15, 3.598988e-15, 
    3.603253e-15, 3.587107e-15, 3.594325e-15, 3.574502e-15, 3.57933e-15, 
    3.57711e-15, 3.574673e-15, 3.582193e-15, 3.590194e-15, 3.590369e-15, 
    3.59293e-15, 3.600145e-15, 3.587736e-15, 3.626119e-15, 3.602427e-15, 
    3.566954e-15, 3.574248e-15, 3.575293e-15, 3.572468e-15, 3.591626e-15, 
    3.58469e-15, 3.603362e-15, 3.59832e-15, 3.606581e-15, 3.602476e-15, 
    3.601873e-15, 3.596598e-15, 3.593312e-15, 3.585007e-15, 3.578244e-15, 
    3.572879e-15, 3.574127e-15, 3.580019e-15, 3.590684e-15, 3.600762e-15, 
    3.598555e-15, 3.605954e-15, 3.586364e-15, 3.594581e-15, 3.591404e-15, 
    3.599685e-15, 3.581535e-15, 3.596983e-15, 3.57758e-15, 3.579284e-15, 
    3.584552e-15, 3.595136e-15, 3.597481e-15, 3.599978e-15, 3.598438e-15, 
    3.590953e-15, 3.58973e-15, 3.584425e-15, 3.582958e-15, 3.578913e-15, 
    3.575562e-15, 3.578624e-15, 3.581836e-15, 3.590958e-15, 3.59917e-15, 
    3.608116e-15, 3.610306e-15, 3.620736e-15, 3.612242e-15, 3.626251e-15, 
    3.614335e-15, 3.634954e-15, 3.597883e-15, 3.613991e-15, 3.584793e-15, 
    3.587944e-15, 3.593636e-15, 3.606687e-15, 3.599647e-15, 3.607881e-15, 
    3.589682e-15, 3.580221e-15, 3.577775e-15, 3.573204e-15, 3.57788e-15, 
    3.5775e-15, 3.581971e-15, 3.580535e-15, 3.591261e-15, 3.585502e-15, 
    3.601856e-15, 3.607817e-15, 3.624632e-15, 3.634922e-15, 3.645389e-15, 
    3.650004e-15, 3.651408e-15, 3.651995e-15 ;

 SMINN_TO_SOIL2N_S1 =
  -8.759354e-09, -8.797866e-09, -8.790379e-09, -8.821442e-09, -8.804211e-09, 
    -8.824551e-09, -8.767161e-09, -8.799396e-09, -8.778818e-09, -8.76282e-09, 
    -8.881726e-09, -8.822828e-09, -8.942898e-09, -8.905337e-09, 
    -8.999689e-09, -8.937054e-09, -9.012319e-09, -8.997882e-09, 
    -9.041331e-09, -9.028883e-09, -9.084461e-09, -9.047077e-09, 
    -9.113269e-09, -9.075533e-09, -9.081437e-09, -9.045843e-09, -8.83468e-09, 
    -8.874393e-09, -8.832327e-09, -8.83799e-09, -8.835449e-09, -8.804567e-09, 
    -8.789005e-09, -8.75641e-09, -8.762327e-09, -8.786267e-09, -8.840536e-09, 
    -8.822114e-09, -8.868541e-09, -8.867493e-09, -8.919179e-09, 
    -8.895875e-09, -8.982747e-09, -8.958057e-09, -9.029403e-09, 
    -9.011461e-09, -9.028561e-09, -9.023376e-09, -9.028629e-09, 
    -9.002313e-09, -9.013588e-09, -8.990432e-09, -8.90024e-09, -8.926747e-09, 
    -8.847689e-09, -8.800153e-09, -8.768575e-09, -8.746168e-09, 
    -8.749336e-09, -8.755375e-09, -8.786407e-09, -8.815582e-09, 
    -8.837815e-09, -8.852687e-09, -8.867342e-09, -8.911701e-09, 
    -8.935175e-09, -8.987739e-09, -8.978253e-09, -8.994324e-09, 
    -9.009676e-09, -9.035451e-09, -9.031209e-09, -9.042565e-09, 
    -8.993899e-09, -9.026243e-09, -8.972849e-09, -8.987453e-09, 
    -8.871329e-09, -8.827083e-09, -8.80828e-09, -8.791818e-09, -8.751772e-09, 
    -8.779428e-09, -8.768525e-09, -8.794461e-09, -8.810941e-09, -8.80279e-09, 
    -8.853094e-09, -8.833537e-09, -8.936567e-09, -8.892189e-09, 
    -9.007885e-09, -8.9802e-09, -9.014521e-09, -8.997008e-09, -9.027016e-09, 
    -9.000009e-09, -9.046791e-09, -9.056978e-09, -9.050017e-09, 
    -9.076757e-09, -8.998511e-09, -9.028561e-09, -8.802562e-09, 
    -8.803891e-09, -8.810084e-09, -8.782862e-09, -8.781196e-09, 
    -8.756247e-09, -8.778446e-09, -8.7879e-09, -8.811896e-09, -8.826091e-09, 
    -8.839584e-09, -8.86925e-09, -8.902384e-09, -8.948712e-09, -8.981995e-09, 
    -9.004305e-09, -8.990624e-09, -9.002703e-09, -8.9892e-09, -8.982872e-09, 
    -9.053161e-09, -9.013693e-09, -9.07291e-09, -9.069634e-09, -9.042835e-09, 
    -9.070003e-09, -8.804824e-09, -8.797175e-09, -8.770615e-09, -8.7914e-09, 
    -8.75353e-09, -8.774728e-09, -8.786918e-09, -8.833948e-09, -8.844279e-09, 
    -8.853861e-09, -8.872783e-09, -8.897068e-09, -8.939669e-09, 
    -8.976733e-09, -9.010568e-09, -9.008089e-09, -9.008962e-09, 
    -9.016521e-09, -8.997798e-09, -9.019595e-09, -9.023253e-09, 
    -9.013688e-09, -9.069195e-09, -9.053337e-09, -9.069564e-09, 
    -9.059239e-09, -8.799661e-09, -8.812534e-09, -8.805578e-09, 
    -8.818658e-09, -8.809443e-09, -8.850416e-09, -8.862701e-09, 
    -8.920181e-09, -8.89659e-09, -8.934133e-09, -8.900404e-09, -8.906381e-09, 
    -8.93536e-09, -8.902227e-09, -8.97469e-09, -8.925563e-09, -9.016815e-09, 
    -8.967759e-09, -9.019889e-09, -9.010422e-09, -9.026096e-09, 
    -9.040134e-09, -9.057794e-09, -9.09038e-09, -9.082834e-09, -9.110084e-09, 
    -8.831722e-09, -8.848418e-09, -8.846948e-09, -8.864419e-09, 
    -8.877341e-09, -8.905346e-09, -8.950263e-09, -8.933372e-09, -8.96438e-09, 
    -8.970605e-09, -8.923496e-09, -8.952421e-09, -8.859591e-09, 
    -8.874591e-09, -8.865659e-09, -8.83304e-09, -8.937266e-09, -8.883778e-09, 
    -8.982544e-09, -8.953569e-09, -9.038133e-09, -8.996079e-09, -9.07868e-09, 
    -9.113993e-09, -9.147224e-09, -9.186063e-09, -8.85753e-09, -8.846185e-09, 
    -8.866497e-09, -8.894601e-09, -8.920673e-09, -8.955337e-09, 
    -8.958883e-09, -8.965377e-09, -8.982197e-09, -8.99634e-09, -8.967431e-09, 
    -8.999885e-09, -8.878071e-09, -8.941908e-09, -8.841897e-09, 
    -8.872014e-09, -8.892943e-09, -8.883761e-09, -8.931441e-09, 
    -8.942679e-09, -8.988345e-09, -8.964738e-09, -9.105278e-09, -9.0431e-09, 
    -9.215633e-09, -9.167418e-09, -8.842222e-09, -8.85749e-09, -8.91063e-09, 
    -8.885346e-09, -8.957651e-09, -8.975448e-09, -8.989915e-09, 
    -9.008411e-09, -9.010407e-09, -9.021365e-09, -9.003408e-09, 
    -9.020655e-09, -8.955411e-09, -8.984567e-09, -8.904555e-09, -8.92403e-09, 
    -8.91507e-09, -8.905244e-09, -8.935573e-09, -8.967887e-09, -8.968576e-09, 
    -8.978937e-09, -9.008137e-09, -8.957944e-09, -9.113306e-09, 
    -9.017361e-09, -8.87414e-09, -8.90355e-09, -8.907749e-09, -8.896357e-09, 
    -8.973664e-09, -8.945653e-09, -9.021098e-09, -9.000708e-09, 
    -9.034116e-09, -9.017515e-09, -9.015072e-09, -8.993751e-09, 
    -8.980476e-09, -8.946938e-09, -8.919649e-09, -8.898009e-09, 
    -8.903041e-09, -8.926812e-09, -8.969863e-09, -9.010588e-09, 
    -9.001667e-09, -9.031577e-09, -8.952408e-09, -8.985606e-09, 
    -8.972775e-09, -9.00623e-09, -8.932924e-09, -8.995352e-09, -8.916967e-09, 
    -8.923839e-09, -8.945097e-09, -8.987858e-09, -8.997317e-09, 
    -9.007419e-09, -9.001185e-09, -8.970956e-09, -8.966002e-09, -8.94458e-09, 
    -8.938666e-09, -8.922343e-09, -8.908829e-09, -8.921177e-09, 
    -8.934143e-09, -8.970967e-09, -9.004153e-09, -9.040334e-09, 
    -9.049187e-09, -9.091464e-09, -9.057051e-09, -9.11384e-09, -9.065562e-09, 
    -9.149133e-09, -8.998968e-09, -9.064139e-09, -8.946064e-09, 
    -8.958785e-09, -8.981793e-09, -9.034562e-09, -9.006073e-09, 
    -9.039391e-09, -8.965809e-09, -8.927633e-09, -8.917754e-09, 
    -8.899325e-09, -8.918176e-09, -8.916642e-09, -8.93468e-09, -8.928883e-09, 
    -8.97219e-09, -8.948928e-09, -9.015012e-09, -9.039127e-09, -9.107229e-09, 
    -9.148978e-09, -9.191472e-09, -9.210233e-09, -9.215944e-09, -9.218331e-09 ;

 SMINN_TO_SOIL3N_S1 =
  -1.039394e-10, -1.043966e-10, -1.043077e-10, -1.046764e-10, -1.044719e-10, 
    -1.047133e-10, -1.040321e-10, -1.044147e-10, -1.041705e-10, 
    -1.039806e-10, -1.053921e-10, -1.046929e-10, -1.061182e-10, 
    -1.056724e-10, -1.067924e-10, -1.060489e-10, -1.069424e-10, -1.06771e-10, 
    -1.072868e-10, -1.07139e-10, -1.077988e-10, -1.07355e-10, -1.081408e-10, 
    -1.076928e-10, -1.077629e-10, -1.073403e-10, -1.048336e-10, -1.05305e-10, 
    -1.048057e-10, -1.048729e-10, -1.048427e-10, -1.044761e-10, 
    -1.042914e-10, -1.039045e-10, -1.039747e-10, -1.042589e-10, 
    -1.049031e-10, -1.046844e-10, -1.052355e-10, -1.052231e-10, 
    -1.058367e-10, -1.0556e-10, -1.065913e-10, -1.062982e-10, -1.071452e-10, 
    -1.069322e-10, -1.071352e-10, -1.070736e-10, -1.07136e-10, -1.068236e-10, 
    -1.069574e-10, -1.066825e-10, -1.056118e-10, -1.059265e-10, -1.04988e-10, 
    -1.044237e-10, -1.040489e-10, -1.037829e-10, -1.038205e-10, 
    -1.038922e-10, -1.042606e-10, -1.046069e-10, -1.048708e-10, 
    -1.050474e-10, -1.052213e-10, -1.057479e-10, -1.060266e-10, 
    -1.066506e-10, -1.065379e-10, -1.067287e-10, -1.06911e-10, -1.07217e-10, 
    -1.071666e-10, -1.073014e-10, -1.067237e-10, -1.071077e-10, 
    -1.064738e-10, -1.066472e-10, -1.052687e-10, -1.047434e-10, 
    -1.045202e-10, -1.043248e-10, -1.038494e-10, -1.041777e-10, 
    -1.040483e-10, -1.043562e-10, -1.045518e-10, -1.04455e-10, -1.050522e-10, 
    -1.0482e-10, -1.060431e-10, -1.055163e-10, -1.068897e-10, -1.065611e-10, 
    -1.069685e-10, -1.067606e-10, -1.071168e-10, -1.067962e-10, 
    -1.073516e-10, -1.074725e-10, -1.073899e-10, -1.077073e-10, 
    -1.067784e-10, -1.071352e-10, -1.044523e-10, -1.044681e-10, 
    -1.045416e-10, -1.042185e-10, -1.041987e-10, -1.039025e-10, 
    -1.041661e-10, -1.042783e-10, -1.045631e-10, -1.047316e-10, 
    -1.048918e-10, -1.05244e-10, -1.056373e-10, -1.061873e-10, -1.065824e-10, 
    -1.068472e-10, -1.066848e-10, -1.068282e-10, -1.066679e-10, 
    -1.065928e-10, -1.074272e-10, -1.069587e-10, -1.076617e-10, 
    -1.076228e-10, -1.073046e-10, -1.076272e-10, -1.044792e-10, 
    -1.043884e-10, -1.040731e-10, -1.043198e-10, -1.038703e-10, 
    -1.041219e-10, -1.042666e-10, -1.048249e-10, -1.049475e-10, 
    -1.050613e-10, -1.052859e-10, -1.055742e-10, -1.060799e-10, 
    -1.065199e-10, -1.069216e-10, -1.068921e-10, -1.069025e-10, 
    -1.069922e-10, -1.0677e-10, -1.070287e-10, -1.070722e-10, -1.069586e-10, 
    -1.076176e-10, -1.074293e-10, -1.076219e-10, -1.074994e-10, 
    -1.044179e-10, -1.045707e-10, -1.044881e-10, -1.046434e-10, -1.04534e-10, 
    -1.050204e-10, -1.051662e-10, -1.058486e-10, -1.055685e-10, 
    -1.060142e-10, -1.056138e-10, -1.056847e-10, -1.060288e-10, 
    -1.056354e-10, -1.064957e-10, -1.059125e-10, -1.069957e-10, 
    -1.064134e-10, -1.070322e-10, -1.069198e-10, -1.071059e-10, 
    -1.072726e-10, -1.074822e-10, -1.078691e-10, -1.077795e-10, -1.08103e-10, 
    -1.047985e-10, -1.049967e-10, -1.049792e-10, -1.051866e-10, -1.0534e-10, 
    -1.056725e-10, -1.062057e-10, -1.060052e-10, -1.063733e-10, 
    -1.064472e-10, -1.058879e-10, -1.062313e-10, -1.051293e-10, 
    -1.053074e-10, -1.052013e-10, -1.048141e-10, -1.060514e-10, 
    -1.054164e-10, -1.065889e-10, -1.062449e-10, -1.072488e-10, 
    -1.067496e-10, -1.077302e-10, -1.081494e-10, -1.085439e-10, -1.09005e-10, 
    -1.051048e-10, -1.049702e-10, -1.052113e-10, -1.055449e-10, 
    -1.058544e-10, -1.062659e-10, -1.06308e-10, -1.063851e-10, -1.065848e-10, 
    -1.067527e-10, -1.064095e-10, -1.067948e-10, -1.053487e-10, 
    -1.061065e-10, -1.049193e-10, -1.052768e-10, -1.055252e-10, 
    -1.054162e-10, -1.059822e-10, -1.061156e-10, -1.066578e-10, 
    -1.063775e-10, -1.080459e-10, -1.073078e-10, -1.093561e-10, 
    -1.087836e-10, -1.049231e-10, -1.051044e-10, -1.057352e-10, -1.05435e-10, 
    -1.062934e-10, -1.065047e-10, -1.066764e-10, -1.06896e-10, -1.069197e-10, 
    -1.070497e-10, -1.068366e-10, -1.070413e-10, -1.062668e-10, 
    -1.066129e-10, -1.056631e-10, -1.058943e-10, -1.057879e-10, 
    -1.056712e-10, -1.060313e-10, -1.064149e-10, -1.064231e-10, 
    -1.065461e-10, -1.068927e-10, -1.062969e-10, -1.081412e-10, 
    -1.070022e-10, -1.05302e-10, -1.056511e-10, -1.05701e-10, -1.055658e-10, 
    -1.064835e-10, -1.061509e-10, -1.070466e-10, -1.068045e-10, 
    -1.072011e-10, -1.07004e-10, -1.06975e-10, -1.067219e-10, -1.065643e-10, 
    -1.061662e-10, -1.058423e-10, -1.055854e-10, -1.056451e-10, 
    -1.059273e-10, -1.064384e-10, -1.069218e-10, -1.068159e-10, -1.07171e-10, 
    -1.062311e-10, -1.066252e-10, -1.064729e-10, -1.068701e-10, 
    -1.059998e-10, -1.067409e-10, -1.058104e-10, -1.05892e-10, -1.061444e-10, 
    -1.06652e-10, -1.067643e-10, -1.068842e-10, -1.068102e-10, -1.064513e-10, 
    -1.063925e-10, -1.061382e-10, -1.06068e-10, -1.058742e-10, -1.057138e-10, 
    -1.058604e-10, -1.060143e-10, -1.064515e-10, -1.068454e-10, 
    -1.072749e-10, -1.0738e-10, -1.078819e-10, -1.074734e-10, -1.081476e-10, 
    -1.075744e-10, -1.085666e-10, -1.067839e-10, -1.075575e-10, 
    -1.061558e-10, -1.063068e-10, -1.0658e-10, -1.072064e-10, -1.068682e-10, 
    -1.072637e-10, -1.063902e-10, -1.05937e-10, -1.058198e-10, -1.05601e-10, 
    -1.058248e-10, -1.058066e-10, -1.060207e-10, -1.059519e-10, -1.06466e-10, 
    -1.061898e-10, -1.069743e-10, -1.072606e-10, -1.080691e-10, 
    -1.085647e-10, -1.090692e-10, -1.09292e-10, -1.093598e-10, -1.093881e-10 ;

 SMINN_TO_SOIL3N_S2 =
  -8.621298e-12, -8.659235e-12, -8.65186e-12, -8.682458e-12, -8.665484e-12, 
    -8.68552e-12, -8.628989e-12, -8.660741e-12, -8.640471e-12, -8.624713e-12, 
    -8.741841e-12, -8.683824e-12, -8.8021e-12, -8.7651e-12, -8.858043e-12, 
    -8.796342e-12, -8.870483e-12, -8.856261e-12, -8.899063e-12, 
    -8.886801e-12, -8.94155e-12, -8.904722e-12, -8.969928e-12, -8.932754e-12, 
    -8.93857e-12, -8.903508e-12, -8.695497e-12, -8.734617e-12, -8.69318e-12, 
    -8.698759e-12, -8.696256e-12, -8.665835e-12, -8.650506e-12, 
    -8.618399e-12, -8.624227e-12, -8.647809e-12, -8.701267e-12, 
    -8.683119e-12, -8.728853e-12, -8.727821e-12, -8.778735e-12, 
    -8.755779e-12, -8.841353e-12, -8.817031e-12, -8.887313e-12, 
    -8.869639e-12, -8.886483e-12, -8.881375e-12, -8.886549e-12, 
    -8.860628e-12, -8.871734e-12, -8.848923e-12, -8.760079e-12, -8.78619e-12, 
    -8.708313e-12, -8.661487e-12, -8.630382e-12, -8.60831e-12, -8.611431e-12, 
    -8.617379e-12, -8.647947e-12, -8.676685e-12, -8.698587e-12, 
    -8.713237e-12, -8.727671e-12, -8.771368e-12, -8.794492e-12, 
    -8.846272e-12, -8.836926e-12, -8.852757e-12, -8.86788e-12, -8.893271e-12, 
    -8.889091e-12, -8.900278e-12, -8.852339e-12, -8.8842e-12, -8.831603e-12, 
    -8.845989e-12, -8.731601e-12, -8.688016e-12, -8.669493e-12, 
    -8.653278e-12, -8.61383e-12, -8.641072e-12, -8.630333e-12, -8.655881e-12, 
    -8.672114e-12, -8.664085e-12, -8.713637e-12, -8.694373e-12, 
    -8.795862e-12, -8.752148e-12, -8.866116e-12, -8.838844e-12, 
    -8.872653e-12, -8.855401e-12, -8.88496e-12, -8.858357e-12, -8.904441e-12, 
    -8.914476e-12, -8.907619e-12, -8.933959e-12, -8.856882e-12, 
    -8.886484e-12, -8.66386e-12, -8.66517e-12, -8.67127e-12, -8.644455e-12, 
    -8.642814e-12, -8.618239e-12, -8.640105e-12, -8.649418e-12, 
    -8.673055e-12, -8.687037e-12, -8.700329e-12, -8.729552e-12, -8.76219e-12, 
    -8.807827e-12, -8.840612e-12, -8.862589e-12, -8.849112e-12, -8.86101e-12, 
    -8.84771e-12, -8.841476e-12, -8.910716e-12, -8.871837e-12, -8.930171e-12, 
    -8.926943e-12, -8.900544e-12, -8.927307e-12, -8.66609e-12, -8.658554e-12, 
    -8.632392e-12, -8.652866e-12, -8.615562e-12, -8.636444e-12, -8.64845e-12, 
    -8.694777e-12, -8.704954e-12, -8.714392e-12, -8.733032e-12, 
    -8.756953e-12, -8.798918e-12, -8.83543e-12, -8.868759e-12, -8.866317e-12, 
    -8.867177e-12, -8.874623e-12, -8.856179e-12, -8.877651e-12, 
    -8.881255e-12, -8.871832e-12, -8.926511e-12, -8.910889e-12, 
    -8.926875e-12, -8.916703e-12, -8.661003e-12, -8.673682e-12, 
    -8.666831e-12, -8.679716e-12, -8.670639e-12, -8.711e-12, -8.7231e-12, 
    -8.779722e-12, -8.756483e-12, -8.793466e-12, -8.76024e-12, -8.766128e-12, 
    -8.794674e-12, -8.762035e-12, -8.833417e-12, -8.785024e-12, 
    -8.874912e-12, -8.826589e-12, -8.877941e-12, -8.868615e-12, 
    -8.884055e-12, -8.897883e-12, -8.91528e-12, -8.947379e-12, -8.939946e-12, 
    -8.96679e-12, -8.692585e-12, -8.709032e-12, -8.707582e-12, -8.724793e-12, 
    -8.737522e-12, -8.765108e-12, -8.809354e-12, -8.792716e-12, 
    -8.823261e-12, -8.829393e-12, -8.782987e-12, -8.81148e-12, -8.720038e-12, 
    -8.734812e-12, -8.726015e-12, -8.693882e-12, -8.796551e-12, 
    -8.743862e-12, -8.841154e-12, -8.812611e-12, -8.895912e-12, 
    -8.854486e-12, -8.935855e-12, -8.970641e-12, -9.003376e-12, 
    -9.041635e-12, -8.718006e-12, -8.706831e-12, -8.72684e-12, -8.754523e-12, 
    -8.780207e-12, -8.814353e-12, -8.817846e-12, -8.824243e-12, 
    -8.840812e-12, -8.854743e-12, -8.826266e-12, -8.858235e-12, -8.73824e-12, 
    -8.801124e-12, -8.702607e-12, -8.732274e-12, -8.752891e-12, 
    -8.743847e-12, -8.790814e-12, -8.801884e-12, -8.846868e-12, 
    -8.823614e-12, -8.962056e-12, -8.900805e-12, -9.070764e-12, 
    -9.023269e-12, -8.702927e-12, -8.717967e-12, -8.770313e-12, 
    -8.745407e-12, -8.816631e-12, -8.834163e-12, -8.848415e-12, 
    -8.866634e-12, -8.8686e-12, -8.879395e-12, -8.861706e-12, -8.878696e-12, 
    -8.814425e-12, -8.843146e-12, -8.764329e-12, -8.783513e-12, 
    -8.774688e-12, -8.765007e-12, -8.794884e-12, -8.826715e-12, 
    -8.827394e-12, -8.8376e-12, -8.866364e-12, -8.81692e-12, -8.969964e-12, 
    -8.87545e-12, -8.734368e-12, -8.763339e-12, -8.767475e-12, -8.756254e-12, 
    -8.832405e-12, -8.804814e-12, -8.879131e-12, -8.859045e-12, 
    -8.891956e-12, -8.875602e-12, -8.873196e-12, -8.852192e-12, 
    -8.839116e-12, -8.806079e-12, -8.779198e-12, -8.757881e-12, 
    -8.762838e-12, -8.786254e-12, -8.828662e-12, -8.868779e-12, 
    -8.859991e-12, -8.889454e-12, -8.811467e-12, -8.844169e-12, -8.83153e-12, 
    -8.864486e-12, -8.792274e-12, -8.85377e-12, -8.776555e-12, -8.783325e-12, 
    -8.804265e-12, -8.846388e-12, -8.855705e-12, -8.865656e-12, 
    -8.859516e-12, -8.829737e-12, -8.824858e-12, -8.803756e-12, 
    -8.797931e-12, -8.781851e-12, -8.768539e-12, -8.780702e-12, 
    -8.793475e-12, -8.829749e-12, -8.86244e-12, -8.89808e-12, -8.906802e-12, 
    -8.948447e-12, -8.914548e-12, -8.97049e-12, -8.922932e-12, -9.005257e-12, 
    -8.857332e-12, -8.92153e-12, -8.805218e-12, -8.817749e-12, -8.840414e-12, 
    -8.892396e-12, -8.864331e-12, -8.897151e-12, -8.824668e-12, 
    -8.787062e-12, -8.77733e-12, -8.759177e-12, -8.777746e-12, -8.776236e-12, 
    -8.794004e-12, -8.788294e-12, -8.830954e-12, -8.808039e-12, 
    -8.873136e-12, -8.896892e-12, -8.963977e-12, -9.005103e-12, 
    -9.046965e-12, -9.065446e-12, -9.071071e-12, -9.073423e-12 ;

 SMIN_NH4 =
  0.0004625078, 0.0004644365, 0.0004640614, 0.000465617, 0.0004647539, 
    0.0004657724, 0.0004628984, 0.0004645127, 0.0004634821, 0.0004626808, 
    0.0004686351, 0.0004656859, 0.0004716969, 0.0004698165, 0.000474539, 
    0.0004714043, 0.0004751708, 0.0004744481, 0.0004766223, 0.0004759994, 
    0.0004787803, 0.0004769096, 0.0004802212, 0.0004783333, 0.0004786287, 
    0.0004768476, 0.0004662796, 0.0004682685, 0.0004661617, 0.0004664453, 
    0.000466318, 0.0004647716, 0.0004639924, 0.0004623597, 0.000462656, 
    0.000463855, 0.0004665724, 0.0004656498, 0.0004679742, 0.0004679217, 
    0.0004705092, 0.0004693426, 0.0004736907, 0.0004724548, 0.0004760253, 
    0.0004751274, 0.000475983, 0.0004757235, 0.0004759863, 0.0004746695, 
    0.0004752336, 0.0004740748, 0.0004695618, 0.0004708887, 0.0004669308, 
    0.0004645507, 0.0004629691, 0.0004618468, 0.0004620054, 0.0004623079, 
    0.0004638619, 0.0004653227, 0.0004664359, 0.0004671804, 0.000467914, 
    0.0004701351, 0.0004713099, 0.0004739406, 0.0004734656, 0.0004742699, 
    0.000475038, 0.0004763277, 0.0004761154, 0.0004766835, 0.0004742482, 
    0.0004758668, 0.0004731946, 0.0004739256, 0.0004681149, 0.0004658989, 
    0.0004649576, 0.000464133, 0.0004621273, 0.0004635124, 0.0004629664, 
    0.000464265, 0.0004650903, 0.000464682, 0.0004672008, 0.0004662215, 
    0.0004713795, 0.000469158, 0.0004749485, 0.0004735629, 0.0004752804, 
    0.000474404, 0.0004759055, 0.000474554, 0.0004768949, 0.0004774047, 
    0.0004770562, 0.000478394, 0.0004744788, 0.0004759826, 0.0004646709, 
    0.0004647375, 0.0004650475, 0.0004636843, 0.0004636009, 0.0004623513, 
    0.000463463, 0.0004639364, 0.0004651379, 0.0004658486, 0.0004665241, 
    0.0004680095, 0.0004696682, 0.0004719871, 0.0004736527, 0.000474769, 
    0.0004740844, 0.0004746887, 0.0004740131, 0.0004736962, 0.0004772135, 
    0.0004752387, 0.0004782014, 0.0004780375, 0.0004766966, 0.0004780558, 
    0.0004647841, 0.0004644009, 0.0004630709, 0.0004641117, 0.0004622151, 
    0.0004632768, 0.0004638872, 0.0004662421, 0.0004667591, 0.0004672389, 
    0.0004681862, 0.0004694019, 0.0004715344, 0.0004733893, 0.0004750824, 
    0.0004749583, 0.0004750019, 0.0004753801, 0.0004744432, 0.0004755338, 
    0.0004757169, 0.0004752382, 0.0004780153, 0.000477222, 0.0004780338, 
    0.0004775171, 0.0004645254, 0.0004651699, 0.0004648215, 0.0004654765, 
    0.000465015, 0.0004670667, 0.0004676817, 0.0004705591, 0.000469378, 
    0.0004712574, 0.0004695687, 0.000469868, 0.0004713188, 0.0004696598, 
    0.000473287, 0.0004708282, 0.0004753948, 0.0004729401, 0.0004755485, 
    0.0004750746, 0.0004758589, 0.0004765614, 0.0004774448, 0.0004790752, 
    0.0004786975, 0.0004800607, 0.0004661306, 0.0004669666, 0.0004668928, 
    0.0004677675, 0.0004684144, 0.0004698163, 0.0004720646, 0.000471219, 
    0.0004727709, 0.0004730825, 0.0004707245, 0.0004721724, 0.0004675254, 
    0.0004682764, 0.0004678291, 0.0004661958, 0.0004714136, 0.0004687361, 
    0.0004736796, 0.0004722293, 0.000476461, 0.0004743568, 0.0004784896, 
    0.0004802565, 0.0004819183, 0.000483861, 0.0004674227, 0.0004668545, 
    0.0004678714, 0.0004692785, 0.0004705834, 0.0004723185, 0.0004724958, 
    0.0004728208, 0.0004736625, 0.0004743703, 0.0004729236, 0.0004745475, 
    0.0004684508, 0.0004716459, 0.0004666391, 0.0004681472, 0.0004691947, 
    0.000468735, 0.0004711216, 0.000471684, 0.0004739696, 0.000472788, 
    0.0004798204, 0.0004767095, 0.0004853393, 0.0004829283, 0.000466656, 
    0.0004674204, 0.0004700807, 0.0004688149, 0.000472434, 0.0004733248, 
    0.0004740487, 0.0004749743, 0.000475074, 0.0004756224, 0.0004747237, 
    0.0004755868, 0.0004723216, 0.0004737808, 0.0004697758, 0.0004707507, 
    0.0004703021, 0.0004698101, 0.0004713282, 0.0004729458, 0.00047298, 
    0.0004734986, 0.0004749605, 0.0004724477, 0.0004802222, 0.0004754217, 
    0.0004682539, 0.0004697264, 0.0004699363, 0.000469366, 0.0004732354, 
    0.0004718335, 0.000475609, 0.0004745886, 0.0004762602, 0.0004754296, 
    0.0004753073, 0.0004742403, 0.0004735758, 0.0004718974, 0.0004705313, 
    0.000469448, 0.0004696997, 0.0004708898, 0.0004730445, 0.0004750825, 
    0.000474636, 0.0004761325, 0.0004721705, 0.0004738321, 0.0004731899, 
    0.000474864, 0.0004711964, 0.0004743215, 0.0004703975, 0.0004707414, 
    0.0004718055, 0.0004739458, 0.0004744188, 0.0004749244, 0.0004746123, 
    0.0004730996, 0.0004728515, 0.0004717792, 0.0004714832, 0.000470666, 
    0.0004699894, 0.0004706076, 0.0004712566, 0.0004730996, 0.0004747604, 
    0.0004765707, 0.0004770136, 0.0004791291, 0.0004774072, 0.0004802487, 
    0.0004778334, 0.0004820137, 0.000474502, 0.000477763, 0.0004718538, 
    0.0004724904, 0.0004736421, 0.0004762827, 0.0004748568, 0.0004765242, 
    0.0004728418, 0.0004709311, 0.0004704363, 0.0004695138, 0.0004704573, 
    0.0004703805, 0.0004712833, 0.0004709931, 0.0004731606, 0.0004719963, 
    0.0004753035, 0.0004765103, 0.0004799173, 0.0004820056, 0.0004841306, 
    0.0004850687, 0.0004853542, 0.0004854736 ;

 SMIN_NH4_vr =
  0.003059624, 0.003064774, 0.003063766, 0.003067918, 0.003065611, 
    0.003068323, 0.003060652, 0.003064957, 0.003062204, 0.003060059, 
    0.003075937, 0.003068077, 0.003084073, 0.003079068, 0.003091607, 
    0.003083288, 0.003093279, 0.003091357, 0.003097117, 0.003095462, 
    0.003102822, 0.00309787, 0.003106624, 0.003101633, 0.003102411, 
    0.003097691, 0.003069681, 0.003074984, 0.00306936, 0.003070117, 
    0.003069773, 0.003065645, 0.003063566, 0.003059199, 0.003059987, 
    0.00306319, 0.003070434, 0.003067969, 0.003074158, 0.003074019, 
    0.003080897, 0.003077795, 0.003089344, 0.003086059, 0.003095528, 
    0.003093143, 0.00309541, 0.003094717, 0.003095409, 0.00309192, 
    0.003093409, 0.003090336, 0.003078415, 0.003081939, 0.003071405, 
    0.003065056, 0.003060827, 0.003057829, 0.003058246, 0.003059056, 
    0.003063202, 0.003067094, 0.003070061, 0.00307204, 0.00307399, 
    0.003079904, 0.003083022, 0.003090001, 0.003088738, 0.003090868, 
    0.003092903, 0.003096316, 0.003095752, 0.003097253, 0.003090793, 
    0.003095086, 0.003087991, 0.003089932, 0.003074561, 0.003068647, 
    0.003066138, 0.003063931, 0.00305857, 0.003062271, 0.003060809, 
    0.00306427, 0.003066471, 0.003065377, 0.003072091, 0.003069476, 
    0.003083202, 0.003077294, 0.00309267, 0.00308899, 0.00309354, 
    0.003091217, 0.003095192, 0.003091609, 0.003097806, 0.003099157, 
    0.003098227, 0.003101768, 0.00309139, 0.003095378, 0.003065365, 
    0.003065544, 0.003066367, 0.003062725, 0.003062501, 0.003059158, 
    0.003062123, 0.003063388, 0.003066589, 0.00306848, 0.003070277, 
    0.003074235, 0.003078646, 0.003084805, 0.003089224, 0.00309218, 
    0.003090363, 0.003091961, 0.003090168, 0.003089322, 0.003098642, 
    0.003093411, 0.00310125, 0.003100816, 0.003097264, 0.003100856, 
    0.003065662, 0.003064635, 0.003061083, 0.003063857, 0.003058788, 
    0.003061625, 0.003063251, 0.003069528, 0.003070901, 0.00307218, 
    0.003074699, 0.00307793, 0.003083598, 0.003088519, 0.003093008, 
    0.003092674, 0.003092788, 0.003093786, 0.003091301, 0.003094188, 
    0.003094669, 0.003093401, 0.003100749, 0.00309865, 0.003100794, 
    0.003099422, 0.003064963, 0.003066678, 0.003065745, 0.003067493, 
    0.003066255, 0.003071727, 0.003073361, 0.003081013, 0.003077866, 
    0.003082865, 0.003078367, 0.003079164, 0.00308302, 0.003078601, 
    0.003088239, 0.003081704, 0.003093822, 0.003087308, 0.003094223, 
    0.003092962, 0.003095036, 0.003096899, 0.003099231, 0.003103546, 
    0.00310254, 0.003106145, 0.003069236, 0.00307146, 0.003071261, 
    0.003073587, 0.003075306, 0.003079036, 0.003085008, 0.003082757, 
    0.003086874, 0.003087703, 0.003081432, 0.003085281, 0.003072917, 
    0.003074913, 0.003073719, 0.003069363, 0.00308325, 0.003076124, 
    0.003089259, 0.003085404, 0.003096624, 0.003091048, 0.003101988, 
    0.003106662, 0.003111044, 0.003116166, 0.003072671, 0.003071152, 
    0.003073857, 0.003077605, 0.003081067, 0.003085678, 0.003086145, 
    0.003087003, 0.003089232, 0.003091111, 0.00308727, 0.003091572, 
    0.003075376, 0.003083865, 0.003070538, 0.003074558, 0.003077338, 
    0.003076115, 0.003082457, 0.003083947, 0.003090012, 0.003086876, 
    0.003105501, 0.00309727, 0.003120054, 0.003113701, 0.00307062, 
    0.003072652, 0.003079729, 0.003076362, 0.003085976, 0.003088342, 
    0.003090255, 0.003092711, 0.003092968, 0.003094423, 0.003092033, 
    0.003094322, 0.003085653, 0.003089527, 0.003078883, 0.003081471, 
    0.003080277, 0.003078964, 0.003082996, 0.003087294, 0.003087379, 
    0.003088752, 0.003092633, 0.003085955, 0.003106554, 0.003093844, 
    0.003074868, 0.003078784, 0.003079336, 0.003077819, 0.003088095, 
    0.003084374, 0.003094387, 0.003091677, 0.003096103, 0.003093903, 
    0.003093572, 0.003090743, 0.003088974, 0.003084519, 0.003080882, 
    0.003078001, 0.003078664, 0.00308183, 0.003087547, 0.003092953, 
    0.003091766, 0.003095726, 0.003085213, 0.003089625, 0.003087914, 
    0.003092355, 0.003082684, 0.003090986, 0.003080557, 0.003081466, 
    0.00308429, 0.003089974, 0.00309122, 0.003092562, 0.003091727, 
    0.003087715, 0.003087053, 0.0030842, 0.00308341, 0.003081238, 
    0.003079432, 0.003081077, 0.003082796, 0.003087691, 0.003092093, 
    0.003096886, 0.003098056, 0.003103653, 0.003099095, 0.003106609, 
    0.003100221, 0.003111262, 0.003091454, 0.003100095, 0.003084419, 
    0.003086105, 0.003089162, 0.003096159, 0.003092374, 0.003096795, 
    0.003087024, 0.003081945, 0.003080624, 0.003078172, 0.003080674, 
    0.003080471, 0.003082866, 0.00308209, 0.003087844, 0.003084752, 
    0.003093522, 0.003096721, 0.003105731, 0.003111242, 0.003116844, 
    0.003119311, 0.003120062, 0.003120373,
  0.001810791, 0.001817542, 0.00181623, 0.001821671, 0.001818652, 
    0.001822215, 0.00181216, 0.00181781, 0.001814203, 0.001811399, 
    0.001832217, 0.001821913, 0.001842897, 0.00183634, 0.001852796, 
    0.001841878, 0.001854995, 0.00185248, 0.001860043, 0.001857877, 
    0.001867542, 0.001861042, 0.001872543, 0.00186599, 0.001867016, 
    0.001860828, 0.001823987, 0.001830936, 0.001823575, 0.001824567, 
    0.001824122, 0.001818715, 0.00181599, 0.001810274, 0.001811312, 
    0.001815509, 0.001825012, 0.001821787, 0.00182991, 0.001829727, 
    0.001838757, 0.001834687, 0.001849844, 0.00184554, 0.001857968, 
    0.001854845, 0.001857821, 0.001856919, 0.001857833, 0.001853252, 
    0.001855216, 0.001851183, 0.00183545, 0.001840078, 0.001826264, 
    0.001817943, 0.001812408, 0.001808478, 0.001809034, 0.001810093, 
    0.001815534, 0.001820644, 0.001824536, 0.001827138, 0.0018297, 
    0.001837453, 0.00184155, 0.001850714, 0.001849061, 0.001851861, 
    0.001854534, 0.00185902, 0.001858282, 0.001860258, 0.001851787, 
    0.001857418, 0.001848119, 0.001850664, 0.0018304, 0.001822658, 
    0.001819367, 0.001816482, 0.001809461, 0.001814311, 0.001812399, 
    0.001816945, 0.001819831, 0.001818404, 0.001827209, 0.001823787, 
    0.001841792, 0.001834044, 0.001854223, 0.0018494, 0.001855378, 
    0.001852328, 0.001857553, 0.001852851, 0.001860993, 0.001862765, 
    0.001861554, 0.001866202, 0.00185259, 0.001857822, 0.001818364, 
    0.001818597, 0.001819681, 0.001814913, 0.001814621, 0.001810246, 
    0.001814138, 0.001815795, 0.001819998, 0.001822484, 0.001824845, 
    0.001830034, 0.001835825, 0.001843911, 0.001849713, 0.001853599, 
    0.001851216, 0.00185332, 0.001850968, 0.001849865, 0.001862101, 
    0.001855234, 0.001865534, 0.001864964, 0.001860305, 0.001865028, 
    0.00181876, 0.00181742, 0.001812766, 0.001816408, 0.001809769, 
    0.001813487, 0.001815624, 0.00182386, 0.001825667, 0.001827343, 
    0.001830652, 0.001834895, 0.001842333, 0.001848796, 0.00185469, 
    0.001854258, 0.00185441, 0.001855726, 0.001852466, 0.001856261, 
    0.001856898, 0.001855233, 0.001864888, 0.001862131, 0.001864952, 
    0.001863157, 0.001817856, 0.00182011, 0.001818892, 0.001821183, 
    0.001819569, 0.001826741, 0.00182889, 0.001838933, 0.001834812, 
    0.001841368, 0.001835478, 0.001836522, 0.001841583, 0.001835796, 
    0.001848441, 0.001839873, 0.001855777, 0.001847233, 0.001856312, 
    0.001854664, 0.001857392, 0.001859835, 0.001862906, 0.001868569, 
    0.001867258, 0.00187199, 0.001823469, 0.001826391, 0.001826133, 
    0.001829189, 0.001831449, 0.001836341, 0.001844181, 0.001841234, 
    0.001846642, 0.001847728, 0.00183951, 0.001844558, 0.001828345, 
    0.001830969, 0.001829406, 0.0018237, 0.001841914, 0.001832574, 
    0.001849809, 0.001844758, 0.001859487, 0.001852167, 0.001866536, 
    0.00187267, 0.001878433, 0.001885164, 0.001827985, 0.001826, 0.001829552, 
    0.001834465, 0.001839018, 0.001845066, 0.001845684, 0.001846816, 
    0.001849748, 0.001852212, 0.001847175, 0.001852829, 0.001831578, 
    0.001842724, 0.00182525, 0.001830518, 0.001834175, 0.001832571, 
    0.001840897, 0.001842858, 0.00185082, 0.001846705, 0.001871157, 
    0.001860352, 0.001890281, 0.001881934, 0.001825307, 0.001827977, 
    0.001837265, 0.001832847, 0.001845469, 0.001848572, 0.001851093, 
    0.001854314, 0.001854662, 0.001856569, 0.001853443, 0.001856446, 
    0.001845079, 0.001850161, 0.001836203, 0.001839604, 0.001838039, 
    0.001836323, 0.001841618, 0.001847255, 0.001847374, 0.00184918, 
    0.00185427, 0.00184552, 0.001872553, 0.001855875, 0.001830889, 
    0.001836029, 0.001836761, 0.001834771, 0.001848261, 0.001843377, 
    0.001856523, 0.001852972, 0.001858788, 0.001855899, 0.001855474, 
    0.001851761, 0.001849448, 0.001843601, 0.001838839, 0.001835059, 
    0.001835939, 0.001840089, 0.001847599, 0.001854693, 0.00185314, 
    0.001858346, 0.001844555, 0.001850342, 0.001848107, 0.001853934, 
    0.001841156, 0.001852043, 0.00183837, 0.00183957, 0.00184328, 
    0.001850736, 0.001852382, 0.001854142, 0.001853056, 0.001847789, 
    0.001846926, 0.001843189, 0.001842158, 0.001839309, 0.001836949, 
    0.001839105, 0.001841369, 0.001847791, 0.001853573, 0.00185987, 
    0.001861409, 0.001868759, 0.001862778, 0.001872646, 0.00186426, 
    0.001878766, 0.001852671, 0.001864011, 0.001843448, 0.001845667, 
    0.001849678, 0.001858867, 0.001853907, 0.001859706, 0.001846892, 
    0.001840233, 0.001838508, 0.00183529, 0.001838581, 0.001838314, 
    0.001841462, 0.00184045, 0.001848004, 0.001843948, 0.001855463, 
    0.00185966, 0.001871495, 0.001878738, 0.001886099, 0.001889347, 
    0.001890334, 0.001890747,
  0.00164664, 0.001653845, 0.001652445, 0.001658253, 0.001655031, 
    0.001658834, 0.001648101, 0.001654131, 0.001650282, 0.001647289, 
    0.001669515, 0.001658512, 0.001680927, 0.001673921, 0.00169151, 
    0.001679838, 0.001693861, 0.001691172, 0.00169926, 0.001696944, 
    0.001707282, 0.001700329, 0.001712635, 0.001705622, 0.00170672, 
    0.0017001, 0.001660727, 0.001668146, 0.001660287, 0.001661345, 
    0.00166087, 0.001655098, 0.001652188, 0.001646089, 0.001647196, 
    0.001651676, 0.001661821, 0.001658378, 0.001667052, 0.001666856, 
    0.001676503, 0.001672155, 0.001688353, 0.001683752, 0.001697041, 
    0.001693701, 0.001696884, 0.001695919, 0.001696897, 0.001691998, 
    0.001694097, 0.001689785, 0.00167297, 0.001677915, 0.001663157, 
    0.001654273, 0.001648366, 0.001644172, 0.001644765, 0.001645896, 
    0.001651702, 0.001657157, 0.001661312, 0.001664091, 0.001666828, 
    0.001675109, 0.001679487, 0.001689284, 0.001687516, 0.00169051, 
    0.001693368, 0.001698166, 0.001697377, 0.00169949, 0.001690431, 
    0.001696453, 0.001686509, 0.00168923, 0.001667574, 0.001659307, 
    0.001655793, 0.001652714, 0.001645221, 0.001650396, 0.001648357, 
    0.001653208, 0.00165629, 0.001654765, 0.001664167, 0.001660513, 
    0.001679747, 0.001671467, 0.001693035, 0.001687879, 0.001694271, 
    0.001691009, 0.001696597, 0.001691568, 0.001700276, 0.001702171, 
    0.001700876, 0.001705849, 0.00169129, 0.001696884, 0.001654723, 
    0.001654972, 0.001656129, 0.001651039, 0.001650727, 0.001646059, 
    0.001650213, 0.001651981, 0.001656468, 0.001659121, 0.001661643, 
    0.001667185, 0.00167337, 0.001682011, 0.001688213, 0.001692368, 
    0.001689821, 0.00169207, 0.001689555, 0.001688376, 0.001701462, 
    0.001694117, 0.001705134, 0.001704525, 0.00169954, 0.001704593, 
    0.001655146, 0.001653715, 0.001648747, 0.001652636, 0.00164555, 
    0.001649517, 0.001651798, 0.00166059, 0.00166252, 0.00166431, 
    0.001667844, 0.001672377, 0.001680325, 0.001687233, 0.001693535, 
    0.001693073, 0.001693236, 0.001694643, 0.001691157, 0.001695215, 
    0.001695896, 0.001694116, 0.001704443, 0.001701494, 0.001704512, 
    0.001702591, 0.00165418, 0.001656587, 0.001655287, 0.001657732, 
    0.00165601, 0.001663667, 0.001665962, 0.001676691, 0.001672288, 
    0.001679293, 0.001673, 0.001674115, 0.001679522, 0.00167334, 0.001686853, 
    0.001677695, 0.001694698, 0.001685562, 0.00169527, 0.001693507, 
    0.001696425, 0.001699038, 0.001702323, 0.001708382, 0.001706979, 
    0.001712043, 0.001660174, 0.001663294, 0.001663019, 0.001666282, 
    0.001668695, 0.001673922, 0.0016823, 0.00167915, 0.001684931, 
    0.001686091, 0.001677308, 0.001682702, 0.001665381, 0.001668182, 
    0.001666514, 0.00166042, 0.001679877, 0.001669897, 0.001688316, 
    0.001682916, 0.001698665, 0.001690837, 0.001706207, 0.00171277, 
    0.00171894, 0.001726147, 0.001664995, 0.001662876, 0.00166667, 
    0.001671917, 0.001676782, 0.001683246, 0.001683906, 0.001685117, 
    0.001688251, 0.001690885, 0.0016855, 0.001691545, 0.001668833, 
    0.001680742, 0.001662075, 0.001667701, 0.001671608, 0.001669894, 
    0.00167879, 0.001680886, 0.001689396, 0.001684998, 0.001711151, 
    0.00169959, 0.001731629, 0.001722688, 0.001662136, 0.001664988, 
    0.001674908, 0.00167019, 0.001683677, 0.001686994, 0.001689689, 
    0.001693133, 0.001693505, 0.001695545, 0.001692201, 0.001695412, 
    0.001683259, 0.001688692, 0.001673774, 0.001677408, 0.001675736, 
    0.001673903, 0.001679561, 0.001685585, 0.001685713, 0.001687644, 
    0.001693084, 0.001683731, 0.001712644, 0.001694801, 0.001668097, 
    0.001673588, 0.001674371, 0.001672245, 0.001686661, 0.00168144, 
    0.001695495, 0.001691699, 0.001697918, 0.001694828, 0.001694373, 
    0.001690403, 0.00168793, 0.00168168, 0.001676591, 0.001672553, 
    0.001673492, 0.001677927, 0.001685953, 0.001693539, 0.001691878, 
    0.001697445, 0.001682699, 0.001688886, 0.001686496, 0.001692727, 
    0.001679067, 0.001690703, 0.00167609, 0.001677372, 0.001681337, 
    0.001689306, 0.001691067, 0.001692948, 0.001691787, 0.001686157, 
    0.001685233, 0.00168124, 0.001680138, 0.001677093, 0.001674572, 
    0.001676876, 0.001679294, 0.001686159, 0.00169234, 0.001699075, 
    0.001700722, 0.001708584, 0.001702186, 0.001712743, 0.00170377, 
    0.001719296, 0.001691376, 0.001703504, 0.001681517, 0.001683888, 
    0.001688176, 0.001698002, 0.001692698, 0.0016989, 0.001685197, 
    0.00167808, 0.001676237, 0.001672799, 0.001676316, 0.00167603, 
    0.001679394, 0.001678313, 0.001686386, 0.001682051, 0.001694362, 
    0.001698851, 0.001711513, 0.001719266, 0.00172715, 0.001730628, 
    0.001731686, 0.001732129,
  0.001515202, 0.001522334, 0.001520947, 0.001526698, 0.001523508, 
    0.001527274, 0.001516648, 0.001522617, 0.001518806, 0.001515844, 
    0.001537857, 0.001526955, 0.001549173, 0.001542224, 0.001559674, 
    0.001548092, 0.001562009, 0.001559339, 0.001567371, 0.00156507, 
    0.001575341, 0.001568432, 0.001580662, 0.001573691, 0.001574782, 
    0.001568204, 0.001529149, 0.0015365, 0.001528713, 0.001529762, 
    0.001529291, 0.001523574, 0.001520693, 0.001514656, 0.001515752, 
    0.001520186, 0.001530233, 0.001526822, 0.001535415, 0.001535221, 
    0.001544785, 0.001540473, 0.001556541, 0.001551975, 0.001565166, 
    0.00156185, 0.00156501, 0.001564052, 0.001565023, 0.001560159, 
    0.001562243, 0.001557962, 0.001541281, 0.001546185, 0.001531557, 
    0.001522758, 0.00151691, 0.00151276, 0.001513346, 0.001514465, 
    0.001520212, 0.001525613, 0.001529729, 0.001532482, 0.001535194, 
    0.001543402, 0.001547744, 0.001557465, 0.00155571, 0.001558682, 
    0.00156152, 0.001566284, 0.0015655, 0.001567599, 0.001558603, 
    0.001564582, 0.001554711, 0.001557411, 0.001535933, 0.001527742, 
    0.001524262, 0.001521214, 0.001513798, 0.001518919, 0.001516901, 
    0.001521703, 0.001524754, 0.001523245, 0.001532557, 0.001528937, 
    0.001548002, 0.001539792, 0.001561189, 0.00155607, 0.001562415, 
    0.001559178, 0.001564725, 0.001559732, 0.00156838, 0.001570262, 
    0.001568976, 0.001573917, 0.001559456, 0.001565011, 0.001523203, 
    0.001523449, 0.001524595, 0.001519555, 0.001519247, 0.001514627, 
    0.001518738, 0.001520488, 0.001524931, 0.001527559, 0.001530056, 
    0.001535547, 0.001541678, 0.001550248, 0.001556402, 0.001560527, 
    0.001557997, 0.00156023, 0.001557734, 0.001556564, 0.001569557, 
    0.001562263, 0.001573206, 0.001572601, 0.001567649, 0.001572669, 
    0.001523622, 0.001522205, 0.001517287, 0.001521136, 0.001514123, 
    0.001518049, 0.001520307, 0.001529013, 0.001530925, 0.001532699, 
    0.001536201, 0.001540694, 0.001548575, 0.001555429, 0.001561685, 
    0.001561226, 0.001561388, 0.001562785, 0.001559324, 0.001563353, 
    0.00156403, 0.001562261, 0.00157252, 0.001569589, 0.001572588, 
    0.00157068, 0.001522666, 0.001525049, 0.001523761, 0.001526183, 
    0.001524477, 0.001532062, 0.001534335, 0.001544971, 0.001540606, 
    0.001547551, 0.001541311, 0.001542417, 0.001547779, 0.001541648, 
    0.001555052, 0.001545966, 0.001562839, 0.001553771, 0.001563408, 
    0.001561658, 0.001564555, 0.00156715, 0.001570413, 0.001576434, 
    0.00157504, 0.001580074, 0.001528601, 0.001531692, 0.001531419, 
    0.001534653, 0.001537044, 0.001542226, 0.001550534, 0.00154741, 
    0.001553145, 0.001554296, 0.001545583, 0.001550934, 0.00153376, 
    0.001536536, 0.001534882, 0.001528845, 0.001548131, 0.001538236, 
    0.001556504, 0.001551146, 0.00156678, 0.001559006, 0.001574272, 
    0.001580796, 0.001586933, 0.001594104, 0.001533378, 0.001531278, 
    0.001535037, 0.001540238, 0.001545061, 0.001551473, 0.001552128, 
    0.001553329, 0.001556439, 0.001559054, 0.00155371, 0.00155971, 
    0.00153718, 0.001548989, 0.001530485, 0.001536059, 0.001539931, 
    0.001538232, 0.001547053, 0.001549131, 0.001557576, 0.001553211, 
    0.001579187, 0.001567698, 0.001599561, 0.001590662, 0.001530544, 
    0.00153337, 0.001543203, 0.001538525, 0.0015519, 0.001555192, 
    0.001557866, 0.001561286, 0.001561655, 0.00156368, 0.001560361, 
    0.001563549, 0.001551486, 0.001556878, 0.001542079, 0.001545682, 
    0.001544025, 0.001542207, 0.001547817, 0.001553794, 0.001553921, 
    0.001555837, 0.001561237, 0.001551954, 0.001580671, 0.001562942, 
    0.001536452, 0.001541894, 0.00154267, 0.001540562, 0.001554862, 
    0.001549682, 0.001563631, 0.001559862, 0.001566037, 0.001562969, 
    0.001562517, 0.001558575, 0.001556121, 0.001549919, 0.001544872, 
    0.001540868, 0.001541799, 0.001546197, 0.001554159, 0.001561688, 
    0.001560039, 0.001565568, 0.001550931, 0.00155707, 0.001554698, 
    0.001560883, 0.001547327, 0.001558873, 0.001544375, 0.001545647, 
    0.001549579, 0.001557487, 0.001559235, 0.001561103, 0.00155995, 
    0.001554361, 0.001553445, 0.001549483, 0.001548389, 0.00154537, 
    0.00154287, 0.001545154, 0.001547553, 0.001554363, 0.001560499, 
    0.001567187, 0.001568823, 0.001576635, 0.001570277, 0.00158077, 
    0.001571851, 0.001587287, 0.001559541, 0.001571587, 0.001549757, 
    0.00155211, 0.001556365, 0.00156612, 0.001560854, 0.001567013, 
    0.001553409, 0.001546349, 0.001544521, 0.001541112, 0.001544599, 
    0.001544315, 0.001547652, 0.00154658, 0.001554589, 0.001550287, 
    0.001562506, 0.001566964, 0.001579546, 0.001587257, 0.001595102, 
    0.001598565, 0.001599618, 0.001600059,
  0.001379622, 0.001386015, 0.001384772, 0.00138993, 0.001387068, 
    0.001390446, 0.001380918, 0.001386269, 0.001382852, 0.001380197, 
    0.001399948, 0.00139016, 0.001410122, 0.001403873, 0.001419577, 
    0.00140915, 0.001421681, 0.001419276, 0.001426515, 0.001424441, 
    0.001433708, 0.001427473, 0.001438514, 0.001432218, 0.001433203, 
    0.001427268, 0.001392128, 0.001398729, 0.001391737, 0.001392678, 
    0.001392256, 0.001387127, 0.001384544, 0.001379134, 0.001380116, 
    0.001384089, 0.001393102, 0.001390041, 0.001397755, 0.00139758, 
    0.001406175, 0.001402299, 0.001416755, 0.001412644, 0.001424527, 
    0.001421538, 0.001424387, 0.001423523, 0.001424398, 0.001420014, 
    0.001421892, 0.001418035, 0.001403025, 0.001407434, 0.00139429, 
    0.001386395, 0.001381153, 0.001377434, 0.00137796, 0.001378962, 
    0.001384112, 0.001388956, 0.001392649, 0.00139512, 0.001397555, 
    0.001404932, 0.001408837, 0.001417587, 0.001416007, 0.001418683, 
    0.00142124, 0.001425535, 0.001424828, 0.001426721, 0.001418612, 
    0.001424001, 0.001415107, 0.001417539, 0.00139822, 0.001390866, 
    0.001387744, 0.001385011, 0.001378364, 0.001382954, 0.001381144, 
    0.001385449, 0.001388185, 0.001386832, 0.001395188, 0.001391939, 
    0.001409068, 0.001401687, 0.001420942, 0.001416331, 0.001422047, 
    0.00141913, 0.00142413, 0.00141963, 0.001427426, 0.001429124, 
    0.001427963, 0.001432422, 0.001419381, 0.001424387, 0.001386794, 
    0.001387015, 0.001388043, 0.001383524, 0.001383247, 0.001379107, 
    0.001382791, 0.00138436, 0.001388344, 0.001390702, 0.001392943, 
    0.001397873, 0.001403382, 0.001411089, 0.00141663, 0.001420346, 
    0.001418067, 0.001420079, 0.00141783, 0.001416776, 0.001428488, 
    0.00142191, 0.001431781, 0.001431234, 0.001426766, 0.001431296, 
    0.00138717, 0.001385899, 0.001381491, 0.001384941, 0.001378656, 
    0.001382174, 0.001384197, 0.001392007, 0.001393723, 0.001395315, 
    0.00139846, 0.001402498, 0.001409584, 0.001415754, 0.001421389, 
    0.001420976, 0.001421121, 0.001422381, 0.001419262, 0.001422893, 
    0.001423503, 0.001421909, 0.001431161, 0.001428517, 0.001431222, 
    0.001429501, 0.001386312, 0.00138845, 0.001387295, 0.001389467, 
    0.001387937, 0.001394743, 0.001396785, 0.001406342, 0.001402418, 
    0.001408663, 0.001403052, 0.001404046, 0.001408868, 0.001403355, 
    0.001415414, 0.001407238, 0.00142243, 0.00141426, 0.001422942, 
    0.001421365, 0.001423976, 0.001426316, 0.00142926, 0.001434695, 
    0.001433436, 0.001437982, 0.001391637, 0.001394411, 0.001394166, 
    0.00139707, 0.001399218, 0.001403874, 0.001411347, 0.001408536, 
    0.001413697, 0.001414733, 0.001406893, 0.001411707, 0.001396268, 
    0.001398761, 0.001397276, 0.001391856, 0.001409185, 0.001400288, 
    0.001416721, 0.001411898, 0.001425982, 0.001418976, 0.001432743, 
    0.001438635, 0.001444182, 0.001450671, 0.001395925, 0.00139404, 
    0.001397415, 0.001402088, 0.001406424, 0.001412192, 0.001412782, 
    0.001413863, 0.001416663, 0.001419019, 0.001414205, 0.001419609, 
    0.00139934, 0.001409957, 0.001393327, 0.001398333, 0.001401812, 
    0.001400285, 0.001408215, 0.001410085, 0.001417688, 0.001413757, 
    0.001437181, 0.001426811, 0.001455612, 0.001447555, 0.001393381, 
    0.001395918, 0.001404753, 0.001400548, 0.001412577, 0.00141554, 
    0.001417949, 0.00142103, 0.001421362, 0.001423188, 0.001420196, 
    0.00142307, 0.001412204, 0.001417058, 0.001403742, 0.001406982, 
    0.001405491, 0.001403857, 0.001408902, 0.001414281, 0.001414395, 
    0.001416121, 0.001420986, 0.001412625, 0.001438522, 0.001422522, 
    0.001398685, 0.001403576, 0.001404274, 0.001402379, 0.001415243, 
    0.00141058, 0.001423143, 0.001419746, 0.001425313, 0.001422546, 
    0.001422139, 0.001418588, 0.001416377, 0.001410794, 0.001406253, 
    0.001402654, 0.001403491, 0.001407445, 0.00141461, 0.001421393, 
    0.001419907, 0.00142489, 0.001411704, 0.001417231, 0.001415095, 
    0.001420666, 0.001408462, 0.001418856, 0.001405807, 0.00140695, 
    0.001410487, 0.001417607, 0.001419181, 0.001420864, 0.001419826, 
    0.001414792, 0.001413967, 0.001410401, 0.001409417, 0.001406701, 
    0.001404453, 0.001406507, 0.001408665, 0.001414794, 0.001420321, 
    0.001426349, 0.001427825, 0.001434876, 0.001429137, 0.001438611, 
    0.001430557, 0.001444502, 0.001419457, 0.001430319, 0.001410648, 
    0.001412765, 0.001416597, 0.001425388, 0.00142064, 0.001426192, 
    0.001413935, 0.001407582, 0.001405938, 0.001402873, 0.001406008, 
    0.001405753, 0.001408754, 0.001407789, 0.001414997, 0.001411125, 
    0.001422129, 0.001426148, 0.001437506, 0.001444475, 0.001451574, 
    0.00145471, 0.001455664, 0.001456063,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3 =
  1.355297e-06, 1.366868e-06, 1.364614e-06, 1.373977e-06, 1.368779e-06, 
    1.374915e-06, 1.357638e-06, 1.367328e-06, 1.361137e-06, 1.356335e-06, 
    1.392239e-06, 1.374394e-06, 1.410893e-06, 1.399422e-06, 1.428326e-06, 
    1.409105e-06, 1.432217e-06, 1.427767e-06, 1.441176e-06, 1.437328e-06, 
    1.454549e-06, 1.442953e-06, 1.463515e-06, 1.451775e-06, 1.453608e-06, 
    1.44257e-06, 1.377975e-06, 1.390012e-06, 1.377264e-06, 1.378977e-06, 
    1.378208e-06, 1.368886e-06, 1.364201e-06, 1.354412e-06, 1.356186e-06, 
    1.363376e-06, 1.379746e-06, 1.374177e-06, 1.388231e-06, 1.387913e-06, 
    1.403643e-06, 1.396539e-06, 1.423112e-06, 1.415533e-06, 1.437488e-06, 
    1.43195e-06, 1.437227e-06, 1.435626e-06, 1.437248e-06, 1.429131e-06, 
    1.432606e-06, 1.425473e-06, 1.39787e-06, 1.405955e-06, 1.381911e-06, 
    1.367557e-06, 1.358061e-06, 1.351345e-06, 1.352293e-06, 1.354103e-06, 
    1.363418e-06, 1.372205e-06, 1.378922e-06, 1.383424e-06, 1.387866e-06, 
    1.401363e-06, 1.40853e-06, 1.424647e-06, 1.42173e-06, 1.426672e-06, 
    1.4314e-06, 1.439356e-06, 1.438045e-06, 1.441556e-06, 1.42654e-06, 
    1.436511e-06, 1.420069e-06, 1.424557e-06, 1.389081e-06, 1.375679e-06, 
    1.370006e-06, 1.365046e-06, 1.353023e-06, 1.36132e-06, 1.358046e-06, 
    1.36584e-06, 1.370806e-06, 1.368348e-06, 1.383547e-06, 1.377628e-06, 
    1.408955e-06, 1.395417e-06, 1.430848e-06, 1.422328e-06, 1.432893e-06, 
    1.427497e-06, 1.43675e-06, 1.428421e-06, 1.442863e-06, 1.446018e-06, 
    1.443862e-06, 1.452153e-06, 1.427959e-06, 1.437226e-06, 1.368281e-06, 
    1.368681e-06, 1.370548e-06, 1.362352e-06, 1.361851e-06, 1.354363e-06, 
    1.361024e-06, 1.363866e-06, 1.371093e-06, 1.375377e-06, 1.379456e-06, 
    1.388446e-06, 1.398521e-06, 1.41267e-06, 1.42288e-06, 1.429744e-06, 
    1.425532e-06, 1.42925e-06, 1.425094e-06, 1.423148e-06, 1.444836e-06, 
    1.432638e-06, 1.450958e-06, 1.449941e-06, 1.441638e-06, 1.450055e-06, 
    1.368962e-06, 1.366657e-06, 1.358673e-06, 1.364919e-06, 1.353548e-06, 
    1.359908e-06, 1.363571e-06, 1.377752e-06, 1.380876e-06, 1.383778e-06, 
    1.389517e-06, 1.396901e-06, 1.409902e-06, 1.421263e-06, 1.431674e-06, 
    1.43091e-06, 1.431179e-06, 1.43351e-06, 1.427739e-06, 1.434458e-06, 
    1.435587e-06, 1.432635e-06, 1.449805e-06, 1.444889e-06, 1.449919e-06, 
    1.446717e-06, 1.367406e-06, 1.371286e-06, 1.369188e-06, 1.373133e-06, 
    1.370353e-06, 1.382736e-06, 1.386459e-06, 1.403948e-06, 1.396756e-06, 
    1.40821e-06, 1.397917e-06, 1.399738e-06, 1.408586e-06, 1.398471e-06, 
    1.420636e-06, 1.405591e-06, 1.4336e-06, 1.418508e-06, 1.434548e-06, 
    1.431628e-06, 1.436464e-06, 1.440802e-06, 1.446269e-06, 1.456385e-06, 
    1.454039e-06, 1.462519e-06, 1.377079e-06, 1.38213e-06, 1.381684e-06, 
    1.386979e-06, 1.390902e-06, 1.399423e-06, 1.413145e-06, 1.407976e-06, 
    1.417471e-06, 1.419381e-06, 1.404958e-06, 1.413805e-06, 1.385514e-06, 
    1.390066e-06, 1.387354e-06, 1.377475e-06, 1.409166e-06, 1.392857e-06, 
    1.423047e-06, 1.414155e-06, 1.440183e-06, 1.42721e-06, 1.452749e-06, 
    1.463739e-06, 1.474116e-06, 1.486295e-06, 1.38489e-06, 1.381453e-06, 
    1.387609e-06, 1.396151e-06, 1.404097e-06, 1.414699e-06, 1.415785e-06, 
    1.417777e-06, 1.422941e-06, 1.427291e-06, 1.418407e-06, 1.428382e-06, 
    1.391124e-06, 1.410586e-06, 1.380154e-06, 1.389283e-06, 1.395644e-06, 
    1.392851e-06, 1.407384e-06, 1.41082e-06, 1.42483e-06, 1.417578e-06, 
    1.461023e-06, 1.44172e-06, 1.4956e-06, 1.480442e-06, 1.380253e-06, 
    1.384877e-06, 1.401033e-06, 1.393334e-06, 1.415407e-06, 1.420868e-06, 
    1.425314e-06, 1.431009e-06, 1.431624e-06, 1.435004e-06, 1.429466e-06, 
    1.434785e-06, 1.41472e-06, 1.423668e-06, 1.399179e-06, 1.40512e-06, 
    1.402385e-06, 1.399389e-06, 1.408646e-06, 1.418545e-06, 1.418755e-06, 
    1.421937e-06, 1.430925e-06, 1.415494e-06, 1.463525e-06, 1.433768e-06, 
    1.389929e-06, 1.398876e-06, 1.400154e-06, 1.396684e-06, 1.420319e-06, 
    1.411732e-06, 1.434921e-06, 1.428635e-06, 1.438942e-06, 1.433815e-06, 
    1.433062e-06, 1.426493e-06, 1.42241e-06, 1.412124e-06, 1.403782e-06, 
    1.397185e-06, 1.398717e-06, 1.405969e-06, 1.419151e-06, 1.431678e-06, 
    1.428929e-06, 1.438155e-06, 1.413798e-06, 1.423986e-06, 1.420044e-06, 
    1.430334e-06, 1.407839e-06, 1.42699e-06, 1.402965e-06, 1.405062e-06, 
    1.411562e-06, 1.424682e-06, 1.427591e-06, 1.430702e-06, 1.428781e-06, 
    1.419487e-06, 1.417967e-06, 1.411402e-06, 1.409593e-06, 1.404604e-06, 
    1.400481e-06, 1.404248e-06, 1.408209e-06, 1.41949e-06, 1.429695e-06, 
    1.440863e-06, 1.443602e-06, 1.456722e-06, 1.446038e-06, 1.463691e-06, 
    1.448679e-06, 1.474714e-06, 1.428101e-06, 1.448239e-06, 1.411857e-06, 
    1.415754e-06, 1.422817e-06, 1.439081e-06, 1.430287e-06, 1.440573e-06, 
    1.417907e-06, 1.406221e-06, 1.403203e-06, 1.397585e-06, 1.403332e-06, 
    1.402864e-06, 1.408373e-06, 1.406601e-06, 1.419864e-06, 1.412732e-06, 
    1.433041e-06, 1.440489e-06, 1.461628e-06, 1.474664e-06, 1.487992e-06, 
    1.493896e-06, 1.495696e-06, 1.496448e-06 ;

 SMIN_NO3_LEACHED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_RUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_vr =
  8.645419e-06, 8.683197e-06, 8.675828e-06, 8.706324e-06, 8.68939e-06, 
    8.709349e-06, 8.653026e-06, 8.684641e-06, 8.664441e-06, 8.648737e-06, 
    8.765499e-06, 8.707612e-06, 8.82565e-06, 8.788669e-06, 8.881559e-06, 
    8.819878e-06, 8.893993e-06, 8.879743e-06, 8.922573e-06, 8.910284e-06, 
    8.96512e-06, 8.928216e-06, 8.99354e-06, 8.956283e-06, 8.962102e-06, 
    8.926957e-06, 8.719308e-06, 8.758357e-06, 8.716981e-06, 8.722548e-06, 
    8.720037e-06, 8.689705e-06, 8.674439e-06, 8.642445e-06, 8.648236e-06, 
    8.671723e-06, 8.724985e-06, 8.706874e-06, 8.752468e-06, 8.751439e-06, 
    8.80225e-06, 8.779327e-06, 8.864821e-06, 8.840488e-06, 8.910786e-06, 
    8.893084e-06, 8.909939e-06, 8.904811e-06, 8.90998e-06, 8.884042e-06, 
    8.895136e-06, 8.872315e-06, 8.783727e-06, 8.809792e-06, 8.732056e-06, 
    8.68538e-06, 8.654378e-06, 8.632409e-06, 8.635495e-06, 8.641419e-06, 
    8.671843e-06, 8.700455e-06, 8.722282e-06, 8.736878e-06, 8.751264e-06, 
    8.794906e-06, 8.817983e-06, 8.869726e-06, 8.860368e-06, 8.876194e-06, 
    8.891314e-06, 8.916714e-06, 8.912525e-06, 8.923714e-06, 8.875722e-06, 
    8.907609e-06, 8.854964e-06, 8.869356e-06, 8.755305e-06, 8.711794e-06, 
    8.693345e-06, 8.677165e-06, 8.637877e-06, 8.665002e-06, 8.654297e-06, 
    8.679719e-06, 8.69589e-06, 8.687874e-06, 8.737267e-06, 8.718044e-06, 
    8.819338e-06, 8.775678e-06, 8.889561e-06, 8.862267e-06, 8.896075e-06, 
    8.878815e-06, 8.90838e-06, 8.881755e-06, 8.927862e-06, 8.937918e-06, 
    8.931028e-06, 8.957412e-06, 8.880225e-06, 8.909853e-06, 8.687703e-06, 
    8.689011e-06, 8.695077e-06, 8.668356e-06, 8.666718e-06, 8.642234e-06, 
    8.663991e-06, 8.67327e-06, 8.696801e-06, 8.710726e-06, 8.723965e-06, 
    8.753116e-06, 8.785686e-06, 8.831258e-06, 8.864025e-06, 8.885992e-06, 
    8.872506e-06, 8.884395e-06, 8.871088e-06, 8.864838e-06, 8.934127e-06, 
    8.895207e-06, 8.953591e-06, 8.950358e-06, 8.923911e-06, 8.950697e-06, 
    8.689909e-06, 8.682386e-06, 8.656331e-06, 8.676703e-06, 8.639552e-06, 
    8.660344e-06, 8.672293e-06, 8.718441e-06, 8.728569e-06, 8.737987e-06, 
    8.756569e-06, 8.780433e-06, 8.822345e-06, 8.858826e-06, 8.892156e-06, 
    8.889699e-06, 8.890555e-06, 8.897994e-06, 8.879536e-06, 8.901006e-06, 
    8.904605e-06, 8.895174e-06, 8.949899e-06, 8.934255e-06, 8.950254e-06, 
    8.94005e-06, 8.684816e-06, 8.697438e-06, 8.690598e-06, 8.703442e-06, 
    8.694377e-06, 8.734622e-06, 8.746682e-06, 8.803188e-06, 8.779964e-06, 
    8.816904e-06, 8.783694e-06, 8.789578e-06, 8.818096e-06, 8.785461e-06, 
    8.856792e-06, 8.808417e-06, 8.898274e-06, 8.84994e-06, 8.901286e-06, 
    8.891939e-06, 8.907378e-06, 8.921227e-06, 8.938625e-06, 8.970793e-06, 
    8.963321e-06, 8.990228e-06, 8.716268e-06, 8.732658e-06, 8.731203e-06, 
    8.748358e-06, 8.761049e-06, 8.788586e-06, 8.832777e-06, 8.816133e-06, 
    8.846648e-06, 8.852781e-06, 8.806384e-06, 8.834863e-06, 8.743543e-06, 
    8.758277e-06, 8.749487e-06, 8.717428e-06, 8.8199e-06, 8.767272e-06, 
    8.864461e-06, 8.83591e-06, 8.919227e-06, 8.877777e-06, 8.959215e-06, 
    8.994096e-06, 9.026899e-06, 9.065294e-06, 8.741597e-06, 8.730433e-06, 
    8.750379e-06, 8.778021e-06, 8.80364e-06, 8.83776e-06, 8.841236e-06, 
    8.847619e-06, 8.864172e-06, 8.878109e-06, 8.849626e-06, 8.881577e-06, 
    8.761701e-06, 8.824464e-06, 8.726109e-06, 8.755712e-06, 8.776263e-06, 
    8.767233e-06, 8.814116e-06, 8.825164e-06, 8.870129e-06, 8.846871e-06, 
    8.985465e-06, 8.924096e-06, 9.094516e-06, 9.046839e-06, 8.726531e-06, 
    8.741516e-06, 8.793757e-06, 8.76889e-06, 8.840008e-06, 8.85754e-06, 
    8.871769e-06, 8.890003e-06, 8.891947e-06, 8.902754e-06, 8.88503e-06, 
    8.902034e-06, 8.837736e-06, 8.866451e-06, 8.787675e-06, 8.806825e-06, 
    8.798002e-06, 8.788322e-06, 8.81815e-06, 8.849976e-06, 8.850633e-06, 
    8.860829e-06, 8.889629e-06, 8.840131e-06, 8.993377e-06, 8.898684e-06, 
    8.757869e-06, 8.786787e-06, 8.790895e-06, 8.77969e-06, 8.855756e-06, 
    8.828178e-06, 8.902489e-06, 8.882374e-06, 8.915298e-06, 8.898932e-06, 
    8.896505e-06, 8.875491e-06, 8.862395e-06, 8.829373e-06, 8.802497e-06, 
    8.781208e-06, 8.786137e-06, 8.809529e-06, 8.851895e-06, 8.892019e-06, 
    8.883217e-06, 8.912682e-06, 8.834664e-06, 8.867366e-06, 8.854708e-06, 
    8.887667e-06, 8.815657e-06, 8.877166e-06, 8.799942e-06, 8.806691e-06, 
    8.827604e-06, 8.869727e-06, 8.879015e-06, 8.888977e-06, 8.882809e-06, 
    8.853035e-06, 8.848143e-06, 8.827034e-06, 8.821205e-06, 8.805137e-06, 
    8.791823e-06, 8.803975e-06, 8.816719e-06, 8.852972e-06, 8.885659e-06, 
    8.921315e-06, 8.930039e-06, 8.971768e-06, 8.937796e-06, 8.993862e-06, 
    8.946198e-06, 9.028701e-06, 8.880689e-06, 8.94496e-06, 8.828554e-06, 
    8.841064e-06, 8.863732e-06, 8.915733e-06, 8.887621e-06, 8.920481e-06, 
    8.847945e-06, 8.810357e-06, 8.800615e-06, 8.782491e-06, 8.801012e-06, 
    8.799506e-06, 8.817242e-06, 8.811523e-06, 8.85415e-06, 8.831244e-06, 
    8.896328e-06, 8.920112e-06, 8.987308e-06, 9.028542e-06, 9.070541e-06, 
    9.089084e-06, 9.09473e-06, 9.097082e-06,
  4.949503e-06, 4.986646e-06, 4.979417e-06, 5.009434e-06, 4.992773e-06, 
    5.012441e-06, 4.957024e-06, 4.988125e-06, 4.968261e-06, 4.95284e-06, 
    5.067877e-06, 5.010774e-06, 5.127414e-06, 5.090822e-06, 5.182911e-06, 
    5.121716e-06, 5.19528e-06, 5.181138e-06, 5.223731e-06, 5.211517e-06, 
    5.266137e-06, 5.229372e-06, 5.294521e-06, 5.257346e-06, 5.263158e-06, 
    5.228162e-06, 5.022243e-06, 5.060756e-06, 5.019966e-06, 5.02545e-06, 
    5.022988e-06, 4.993119e-06, 4.978093e-06, 4.946665e-06, 4.952365e-06, 
    4.975449e-06, 5.027917e-06, 5.010081e-06, 5.055066e-06, 5.054048e-06, 
    5.104295e-06, 5.081618e-06, 5.166329e-06, 5.142202e-06, 5.212026e-06, 
    5.194436e-06, 5.2112e-06, 5.206114e-06, 5.211266e-06, 5.185477e-06, 
    5.196521e-06, 5.173846e-06, 5.085864e-06, 5.111668e-06, 5.034846e-06, 
    4.988859e-06, 4.958387e-06, 4.936808e-06, 4.939856e-06, 4.945671e-06, 
    4.975584e-06, 5.003764e-06, 5.025279e-06, 5.039689e-06, 5.053902e-06, 
    5.09702e-06, 5.119884e-06, 5.171215e-06, 5.161934e-06, 5.177657e-06, 
    5.192687e-06, 5.217961e-06, 5.213797e-06, 5.224943e-06, 5.177239e-06, 
    5.208928e-06, 5.156652e-06, 5.170932e-06, 5.057783e-06, 5.01489e-06, 
    4.996711e-06, 4.980806e-06, 4.942201e-06, 4.968851e-06, 4.958339e-06, 
    4.983356e-06, 4.999278e-06, 4.9914e-06, 5.040084e-06, 5.021137e-06, 
    5.12124e-06, 5.078037e-06, 5.190933e-06, 5.163839e-06, 5.197434e-06, 
    5.180281e-06, 5.209685e-06, 5.183219e-06, 5.229092e-06, 5.239101e-06, 
    5.232261e-06, 5.258549e-06, 5.181753e-06, 5.211201e-06, 4.991181e-06, 
    4.992465e-06, 4.998449e-06, 4.972163e-06, 4.970556e-06, 4.94651e-06, 
    4.967903e-06, 4.977024e-06, 5.0002e-06, 5.01393e-06, 5.026992e-06, 
    5.055756e-06, 5.08795e-06, 5.133084e-06, 5.165593e-06, 5.187426e-06, 
    5.174034e-06, 5.185856e-06, 5.172641e-06, 5.166451e-06, 5.235352e-06, 
    5.196625e-06, 5.254765e-06, 5.251542e-06, 5.225209e-06, 5.251905e-06, 
    4.993367e-06, 4.985976e-06, 4.960353e-06, 4.980402e-06, 4.943894e-06, 
    4.964319e-06, 4.976078e-06, 5.021536e-06, 5.03154e-06, 5.040827e-06, 
    5.059184e-06, 5.082778e-06, 5.124262e-06, 5.160451e-06, 5.193561e-06, 
    5.191133e-06, 5.191988e-06, 5.199395e-06, 5.181055e-06, 5.202408e-06, 
    5.205996e-06, 5.196619e-06, 5.25111e-06, 5.235522e-06, 5.251473e-06, 
    5.241321e-06, 4.988378e-06, 5.000817e-06, 4.994094e-06, 5.006739e-06, 
    4.997831e-06, 5.037491e-06, 5.049403e-06, 5.105273e-06, 5.082315e-06, 
    5.118867e-06, 5.086022e-06, 5.091837e-06, 5.120067e-06, 5.087794e-06, 
    5.158456e-06, 5.110518e-06, 5.199684e-06, 5.151684e-06, 5.202697e-06, 
    5.193418e-06, 5.208782e-06, 5.222557e-06, 5.239901e-06, 5.271961e-06, 
    5.264531e-06, 5.291377e-06, 5.01938e-06, 5.035553e-06, 5.034125e-06, 
    5.051067e-06, 5.06361e-06, 5.09083e-06, 5.134596e-06, 5.118122e-06, 
    5.148378e-06, 5.15446e-06, 5.108498e-06, 5.136704e-06, 5.046385e-06, 
    5.060942e-06, 5.052271e-06, 5.020656e-06, 5.121921e-06, 5.069864e-06, 
    5.166132e-06, 5.137823e-06, 5.220592e-06, 5.179375e-06, 5.260442e-06, 
    5.295237e-06, 5.328041e-06, 5.36648e-06, 5.044385e-06, 5.033387e-06, 
    5.053082e-06, 5.080382e-06, 5.10575e-06, 5.139549e-06, 5.143009e-06, 
    5.149352e-06, 5.165791e-06, 5.179628e-06, 5.151361e-06, 5.183098e-06, 
    5.064326e-06, 5.126446e-06, 5.029233e-06, 5.058441e-06, 5.07877e-06, 
    5.069846e-06, 5.11624e-06, 5.127196e-06, 5.171806e-06, 5.148727e-06, 
    5.286645e-06, 5.225472e-06, 5.3958e-06, 5.348017e-06, 5.029547e-06, 
    5.044345e-06, 5.095973e-06, 5.071385e-06, 5.141806e-06, 5.159193e-06, 
    5.17334e-06, 5.191449e-06, 5.193403e-06, 5.204144e-06, 5.186548e-06, 
    5.203447e-06, 5.13962e-06, 5.16811e-06, 5.090059e-06, 5.10902e-06, 
    5.100293e-06, 5.090729e-06, 5.120267e-06, 5.151806e-06, 5.152477e-06, 
    5.162605e-06, 5.191192e-06, 5.142092e-06, 5.294567e-06, 5.200228e-06, 
    5.0605e-06, 5.089086e-06, 5.093169e-06, 5.082086e-06, 5.157449e-06, 
    5.130098e-06, 5.203881e-06, 5.183903e-06, 5.21665e-06, 5.200369e-06, 
    5.197975e-06, 5.177093e-06, 5.164108e-06, 5.131352e-06, 5.104753e-06, 
    5.083692e-06, 5.088586e-06, 5.11173e-06, 5.153737e-06, 5.193583e-06, 
    5.184846e-06, 5.214159e-06, 5.136689e-06, 5.169127e-06, 5.156582e-06, 
    5.189312e-06, 5.117685e-06, 5.178672e-06, 5.102139e-06, 5.108832e-06, 
    5.129556e-06, 5.171332e-06, 5.180584e-06, 5.190477e-06, 5.184371e-06, 
    5.154804e-06, 5.149963e-06, 5.129051e-06, 5.123284e-06, 5.107374e-06, 
    5.094218e-06, 5.106239e-06, 5.118875e-06, 5.154815e-06, 5.187279e-06, 
    5.222754e-06, 5.231446e-06, 5.273034e-06, 5.239177e-06, 5.295094e-06, 
    5.247551e-06, 5.329938e-06, 5.182206e-06, 5.246146e-06, 5.130498e-06, 
    5.142913e-06, 5.165399e-06, 5.217093e-06, 5.189158e-06, 5.22183e-06, 
    5.149774e-06, 5.112532e-06, 5.102906e-06, 5.084973e-06, 5.103316e-06, 
    5.101823e-06, 5.119396e-06, 5.113746e-06, 5.156009e-06, 5.133292e-06, 
    5.197916e-06, 5.221571e-06, 5.288563e-06, 5.329778e-06, 5.371835e-06, 
    5.39044e-06, 5.396107e-06, 5.398477e-06,
  4.464165e-06, 4.503465e-06, 4.495813e-06, 4.527595e-06, 4.509952e-06, 
    4.53078e-06, 4.47212e-06, 4.505029e-06, 4.484009e-06, 4.467695e-06, 
    4.589539e-06, 4.529014e-06, 4.652746e-06, 4.613891e-06, 4.711746e-06, 
    4.646692e-06, 4.724908e-06, 4.709862e-06, 4.755199e-06, 4.742193e-06, 
    4.80038e-06, 4.761207e-06, 4.830652e-06, 4.791012e-06, 4.797205e-06, 
    4.759917e-06, 4.541165e-06, 4.581986e-06, 4.538752e-06, 4.544562e-06, 
    4.541954e-06, 4.510317e-06, 4.494411e-06, 4.461166e-06, 4.467193e-06, 
    4.491613e-06, 4.547176e-06, 4.528281e-06, 4.575957e-06, 4.574878e-06, 
    4.628193e-06, 4.604124e-06, 4.694111e-06, 4.668462e-06, 4.742735e-06, 
    4.724011e-06, 4.741855e-06, 4.736441e-06, 4.741926e-06, 4.714478e-06, 
    4.72623e-06, 4.702106e-06, 4.608628e-06, 4.636022e-06, 4.55452e-06, 
    4.505805e-06, 4.473562e-06, 4.450742e-06, 4.453965e-06, 4.460113e-06, 
    4.491756e-06, 4.521591e-06, 4.544382e-06, 4.559654e-06, 4.574723e-06, 
    4.620466e-06, 4.644747e-06, 4.699306e-06, 4.689438e-06, 4.706158e-06, 
    4.722151e-06, 4.749053e-06, 4.744621e-06, 4.756489e-06, 4.705715e-06, 
    4.739436e-06, 4.683821e-06, 4.699006e-06, 4.578833e-06, 4.533375e-06, 
    4.514119e-06, 4.497284e-06, 4.456444e-06, 4.484632e-06, 4.473511e-06, 
    4.499984e-06, 4.516839e-06, 4.508499e-06, 4.560072e-06, 4.539993e-06, 
    4.646187e-06, 4.600322e-06, 4.720284e-06, 4.691462e-06, 4.727202e-06, 
    4.708951e-06, 4.740242e-06, 4.712077e-06, 4.760908e-06, 4.77157e-06, 
    4.764283e-06, 4.792294e-06, 4.710517e-06, 4.741856e-06, 4.508266e-06, 
    4.509626e-06, 4.515962e-06, 4.488137e-06, 4.486436e-06, 4.461001e-06, 
    4.483629e-06, 4.493281e-06, 4.517817e-06, 4.532357e-06, 4.546197e-06, 
    4.576688e-06, 4.610841e-06, 4.658771e-06, 4.693329e-06, 4.716552e-06, 
    4.702306e-06, 4.714883e-06, 4.700824e-06, 4.694241e-06, 4.767574e-06, 
    4.72634e-06, 4.788261e-06, 4.784826e-06, 4.756772e-06, 4.785213e-06, 
    4.510581e-06, 4.502757e-06, 4.475642e-06, 4.496856e-06, 4.458234e-06, 
    4.479837e-06, 4.492279e-06, 4.540415e-06, 4.551017e-06, 4.56086e-06, 
    4.580324e-06, 4.605354e-06, 4.649399e-06, 4.68786e-06, 4.723081e-06, 
    4.720497e-06, 4.721407e-06, 4.729289e-06, 4.709774e-06, 4.732496e-06, 
    4.736315e-06, 4.726334e-06, 4.784366e-06, 4.767758e-06, 4.784753e-06, 
    4.773936e-06, 4.505299e-06, 4.518469e-06, 4.511351e-06, 4.524741e-06, 
    4.515307e-06, 4.557322e-06, 4.569951e-06, 4.629231e-06, 4.604862e-06, 
    4.643667e-06, 4.608797e-06, 4.614968e-06, 4.644939e-06, 4.610677e-06, 
    4.685738e-06, 4.634799e-06, 4.729596e-06, 4.678537e-06, 4.732803e-06, 
    4.722929e-06, 4.739281e-06, 4.753947e-06, 4.772423e-06, 4.806592e-06, 
    4.79867e-06, 4.8273e-06, 4.538132e-06, 4.555269e-06, 4.553757e-06, 
    4.571717e-06, 4.585018e-06, 4.613899e-06, 4.660379e-06, 4.642877e-06, 
    4.675026e-06, 4.681491e-06, 4.632657e-06, 4.662617e-06, 4.566752e-06, 
    4.582187e-06, 4.572993e-06, 4.539484e-06, 4.64691e-06, 4.591651e-06, 
    4.693901e-06, 4.663807e-06, 4.751856e-06, 4.707986e-06, 4.794312e-06, 
    4.831415e-06, 4.86643e-06, 4.907489e-06, 4.564631e-06, 4.552974e-06, 
    4.573853e-06, 4.60281e-06, 4.629738e-06, 4.665641e-06, 4.66932e-06, 
    4.676061e-06, 4.693539e-06, 4.708256e-06, 4.678195e-06, 4.711948e-06, 
    4.585773e-06, 4.651719e-06, 4.548572e-06, 4.579534e-06, 4.6011e-06, 
    4.591633e-06, 4.640878e-06, 4.652517e-06, 4.699935e-06, 4.675397e-06, 
    4.822249e-06, 4.757051e-06, 4.938837e-06, 4.887761e-06, 4.548905e-06, 
    4.56459e-06, 4.619358e-06, 4.593266e-06, 4.668041e-06, 4.686523e-06, 
    4.701568e-06, 4.720832e-06, 4.722913e-06, 4.734344e-06, 4.715618e-06, 
    4.733603e-06, 4.665717e-06, 4.696004e-06, 4.613082e-06, 4.63321e-06, 
    4.623945e-06, 4.613793e-06, 4.645156e-06, 4.678669e-06, 4.679383e-06, 
    4.69015e-06, 4.720554e-06, 4.668344e-06, 4.830696e-06, 4.730171e-06, 
    4.58172e-06, 4.612047e-06, 4.616381e-06, 4.60462e-06, 4.684669e-06, 
    4.655599e-06, 4.734065e-06, 4.712805e-06, 4.747658e-06, 4.730326e-06, 
    4.727779e-06, 4.70556e-06, 4.691749e-06, 4.656931e-06, 4.628679e-06, 
    4.606325e-06, 4.611519e-06, 4.636088e-06, 4.680721e-06, 4.723103e-06, 
    4.713806e-06, 4.745005e-06, 4.662602e-06, 4.697085e-06, 4.683746e-06, 
    4.718559e-06, 4.642413e-06, 4.707234e-06, 4.625905e-06, 4.633011e-06, 
    4.655023e-06, 4.699431e-06, 4.709274e-06, 4.719798e-06, 4.713302e-06, 
    4.681855e-06, 4.67671e-06, 4.654487e-06, 4.64836e-06, 4.631464e-06, 
    4.617496e-06, 4.630258e-06, 4.643677e-06, 4.681868e-06, 4.716396e-06, 
    4.754157e-06, 4.763415e-06, 4.807733e-06, 4.771648e-06, 4.831258e-06, 
    4.780566e-06, 4.86845e-06, 4.710996e-06, 4.779072e-06, 4.656025e-06, 
    4.669217e-06, 4.693121e-06, 4.748127e-06, 4.718395e-06, 4.753172e-06, 
    4.676509e-06, 4.636938e-06, 4.626719e-06, 4.607683e-06, 4.627154e-06, 
    4.62557e-06, 4.644231e-06, 4.63823e-06, 4.683138e-06, 4.658993e-06, 
    4.727715e-06, 4.752896e-06, 4.824297e-06, 4.868282e-06, 4.913215e-06, 
    4.933107e-06, 4.939167e-06, 4.941701e-06,
  4.333261e-06, 4.374273e-06, 4.366284e-06, 4.399469e-06, 4.381045e-06, 
    4.402797e-06, 4.341559e-06, 4.375906e-06, 4.353964e-06, 4.336944e-06, 
    4.464212e-06, 4.400952e-06, 4.53036e-06, 4.489686e-06, 4.592185e-06, 
    4.524021e-06, 4.605987e-06, 4.590208e-06, 4.637766e-06, 4.624118e-06, 
    4.685206e-06, 4.644071e-06, 4.717015e-06, 4.675365e-06, 4.681871e-06, 
    4.642718e-06, 4.413645e-06, 4.456314e-06, 4.411124e-06, 4.417195e-06, 
    4.41447e-06, 4.381427e-06, 4.364822e-06, 4.330132e-06, 4.336419e-06, 
    4.361901e-06, 4.419926e-06, 4.400186e-06, 4.450008e-06, 4.448881e-06, 
    4.504654e-06, 4.479467e-06, 4.573697e-06, 4.54682e-06, 4.624687e-06, 
    4.605046e-06, 4.623764e-06, 4.618084e-06, 4.623838e-06, 4.595049e-06, 
    4.607374e-06, 4.582078e-06, 4.484179e-06, 4.512849e-06, 4.4276e-06, 
    4.376716e-06, 4.343064e-06, 4.319261e-06, 4.322622e-06, 4.329034e-06, 
    4.362051e-06, 4.393198e-06, 4.417006e-06, 4.432966e-06, 4.448718e-06, 
    4.496568e-06, 4.521984e-06, 4.579143e-06, 4.568799e-06, 4.586326e-06, 
    4.603095e-06, 4.631317e-06, 4.626665e-06, 4.63912e-06, 4.585861e-06, 
    4.621226e-06, 4.562913e-06, 4.578828e-06, 4.453017e-06, 4.405507e-06, 
    4.385396e-06, 4.36782e-06, 4.325208e-06, 4.354614e-06, 4.343011e-06, 
    4.370638e-06, 4.388237e-06, 4.379528e-06, 4.433403e-06, 4.412421e-06, 
    4.523492e-06, 4.475491e-06, 4.601137e-06, 4.570921e-06, 4.608393e-06, 
    4.589253e-06, 4.622072e-06, 4.592531e-06, 4.643759e-06, 4.65495e-06, 
    4.647301e-06, 4.676712e-06, 4.590896e-06, 4.623766e-06, 4.379284e-06, 
    4.380704e-06, 4.387321e-06, 4.358273e-06, 4.356498e-06, 4.32996e-06, 
    4.353569e-06, 4.363641e-06, 4.389257e-06, 4.404444e-06, 4.418903e-06, 
    4.450773e-06, 4.486496e-06, 4.53667e-06, 4.572877e-06, 4.597224e-06, 
    4.582287e-06, 4.595473e-06, 4.580734e-06, 4.573833e-06, 4.650756e-06, 
    4.607489e-06, 4.672476e-06, 4.668868e-06, 4.639417e-06, 4.669275e-06, 
    4.381701e-06, 4.373533e-06, 4.345234e-06, 4.367373e-06, 4.327074e-06, 
    4.349612e-06, 4.362596e-06, 4.412862e-06, 4.42394e-06, 4.434227e-06, 
    4.454575e-06, 4.480754e-06, 4.526855e-06, 4.567145e-06, 4.60407e-06, 
    4.60136e-06, 4.602314e-06, 4.610582e-06, 4.590117e-06, 4.613946e-06, 
    4.617952e-06, 4.607483e-06, 4.668385e-06, 4.650948e-06, 4.668792e-06, 
    4.657434e-06, 4.376187e-06, 4.389939e-06, 4.382506e-06, 4.396489e-06, 
    4.386636e-06, 4.43053e-06, 4.44373e-06, 4.50574e-06, 4.480239e-06, 
    4.520853e-06, 4.484356e-06, 4.490813e-06, 4.522186e-06, 4.486324e-06, 
    4.564922e-06, 4.511569e-06, 4.610903e-06, 4.557377e-06, 4.614268e-06, 
    4.60391e-06, 4.621063e-06, 4.636453e-06, 4.655845e-06, 4.691731e-06, 
    4.683409e-06, 4.713491e-06, 4.410476e-06, 4.428383e-06, 4.426803e-06, 
    4.445576e-06, 4.459483e-06, 4.489695e-06, 4.538354e-06, 4.520026e-06, 
    4.553697e-06, 4.560471e-06, 4.509326e-06, 4.540699e-06, 4.440386e-06, 
    4.456523e-06, 4.44691e-06, 4.411889e-06, 4.52425e-06, 4.46642e-06, 
    4.573477e-06, 4.541945e-06, 4.634257e-06, 4.588242e-06, 4.678831e-06, 
    4.717817e-06, 4.754636e-06, 4.797847e-06, 4.438169e-06, 4.425985e-06, 
    4.44781e-06, 4.478093e-06, 4.506271e-06, 4.543866e-06, 4.547719e-06, 
    4.554782e-06, 4.573098e-06, 4.588525e-06, 4.557018e-06, 4.592396e-06, 
    4.460274e-06, 4.529285e-06, 4.421384e-06, 4.45375e-06, 4.476304e-06, 
    4.466401e-06, 4.517933e-06, 4.53012e-06, 4.579802e-06, 4.554086e-06, 
    4.708183e-06, 4.63971e-06, 4.830863e-06, 4.777082e-06, 4.421732e-06, 
    4.438125e-06, 4.495407e-06, 4.468109e-06, 4.546379e-06, 4.565745e-06, 
    4.581514e-06, 4.601713e-06, 4.603894e-06, 4.615884e-06, 4.596244e-06, 
    4.615106e-06, 4.543946e-06, 4.575681e-06, 4.488839e-06, 4.509905e-06, 
    4.500208e-06, 4.489583e-06, 4.522412e-06, 4.557514e-06, 4.558262e-06, 
    4.569546e-06, 4.601422e-06, 4.546698e-06, 4.717062e-06, 4.611508e-06, 
    4.456035e-06, 4.487757e-06, 4.492292e-06, 4.479986e-06, 4.563802e-06, 
    4.533348e-06, 4.615591e-06, 4.593294e-06, 4.629852e-06, 4.611669e-06, 
    4.608997e-06, 4.585698e-06, 4.571222e-06, 4.534743e-06, 4.505163e-06, 
    4.48177e-06, 4.487204e-06, 4.512919e-06, 4.559665e-06, 4.604093e-06, 
    4.594344e-06, 4.627069e-06, 4.540683e-06, 4.576815e-06, 4.562835e-06, 
    4.599329e-06, 4.51954e-06, 4.587454e-06, 4.502259e-06, 4.509698e-06, 
    4.532745e-06, 4.579273e-06, 4.589592e-06, 4.600628e-06, 4.593816e-06, 
    4.560854e-06, 4.555463e-06, 4.532183e-06, 4.525767e-06, 4.508077e-06, 
    4.493458e-06, 4.506815e-06, 4.520863e-06, 4.560866e-06, 4.59706e-06, 
    4.636673e-06, 4.64639e-06, 4.692931e-06, 4.655033e-06, 4.717654e-06, 
    4.664397e-06, 4.756763e-06, 4.591399e-06, 4.662828e-06, 4.533793e-06, 
    4.547612e-06, 4.57266e-06, 4.630345e-06, 4.599156e-06, 4.635639e-06, 
    4.555251e-06, 4.513809e-06, 4.503111e-06, 4.483191e-06, 4.503567e-06, 
    4.501908e-06, 4.521443e-06, 4.515161e-06, 4.562197e-06, 4.536902e-06, 
    4.608931e-06, 4.63535e-06, 4.710336e-06, 4.756586e-06, 4.803876e-06, 
    4.824826e-06, 4.83121e-06, 4.833881e-06,
  4.365279e-06, 4.405926e-06, 4.398006e-06, 4.430915e-06, 4.412641e-06, 
    4.434216e-06, 4.3735e-06, 4.407545e-06, 4.385794e-06, 4.368927e-06, 
    4.495183e-06, 4.432386e-06, 4.560928e-06, 4.520489e-06, 4.622458e-06, 
    4.554624e-06, 4.636205e-06, 4.620489e-06, 4.667872e-06, 4.654269e-06, 
    4.715187e-06, 4.674157e-06, 4.746938e-06, 4.705367e-06, 4.711858e-06, 
    4.672808e-06, 4.444979e-06, 4.487339e-06, 4.442477e-06, 4.448502e-06, 
    4.445797e-06, 4.41302e-06, 4.396557e-06, 4.362178e-06, 4.368407e-06, 
    4.393661e-06, 4.451212e-06, 4.431626e-06, 4.481074e-06, 4.479954e-06, 
    4.535367e-06, 4.510334e-06, 4.604049e-06, 4.5773e-06, 4.654836e-06, 
    4.635267e-06, 4.653916e-06, 4.648256e-06, 4.65399e-06, 4.625309e-06, 
    4.637585e-06, 4.612392e-06, 4.515017e-06, 4.543514e-06, 4.458828e-06, 
    4.40835e-06, 4.374991e-06, 4.35141e-06, 4.354739e-06, 4.361091e-06, 
    4.393809e-06, 4.424694e-06, 4.448314e-06, 4.464154e-06, 4.479793e-06, 
    4.52733e-06, 4.552597e-06, 4.609471e-06, 4.599173e-06, 4.616623e-06, 
    4.633323e-06, 4.661443e-06, 4.656808e-06, 4.669222e-06, 4.616159e-06, 
    4.651387e-06, 4.593314e-06, 4.609157e-06, 4.484064e-06, 4.436904e-06, 
    4.416957e-06, 4.399529e-06, 4.3573e-06, 4.386438e-06, 4.374939e-06, 
    4.402322e-06, 4.419773e-06, 4.411137e-06, 4.464588e-06, 4.443764e-06, 
    4.554097e-06, 4.506384e-06, 4.631373e-06, 4.601286e-06, 4.638601e-06, 
    4.619537e-06, 4.65223e-06, 4.622801e-06, 4.673845e-06, 4.685005e-06, 
    4.677378e-06, 4.70671e-06, 4.621173e-06, 4.653918e-06, 4.410895e-06, 
    4.412303e-06, 4.418865e-06, 4.390065e-06, 4.388306e-06, 4.362008e-06, 
    4.385402e-06, 4.395386e-06, 4.420785e-06, 4.43585e-06, 4.450197e-06, 
    4.481833e-06, 4.517319e-06, 4.567204e-06, 4.603232e-06, 4.627475e-06, 
    4.6126e-06, 4.625731e-06, 4.611054e-06, 4.604184e-06, 4.680823e-06, 
    4.637701e-06, 4.702485e-06, 4.698886e-06, 4.669518e-06, 4.699291e-06, 
    4.413292e-06, 4.405192e-06, 4.377142e-06, 4.399085e-06, 4.359149e-06, 
    4.38148e-06, 4.39435e-06, 4.444202e-06, 4.455194e-06, 4.465406e-06, 
    4.485608e-06, 4.511613e-06, 4.557441e-06, 4.597528e-06, 4.634295e-06, 
    4.631595e-06, 4.632545e-06, 4.640782e-06, 4.620397e-06, 4.644133e-06, 
    4.648125e-06, 4.637694e-06, 4.698404e-06, 4.681013e-06, 4.698809e-06, 
    4.687481e-06, 4.407824e-06, 4.421461e-06, 4.414089e-06, 4.427958e-06, 
    4.418186e-06, 4.461736e-06, 4.474841e-06, 4.536447e-06, 4.511101e-06, 
    4.551473e-06, 4.515192e-06, 4.521609e-06, 4.552799e-06, 4.517147e-06, 
    4.595315e-06, 4.542242e-06, 4.641102e-06, 4.587807e-06, 4.644454e-06, 
    4.634135e-06, 4.651225e-06, 4.666563e-06, 4.685897e-06, 4.721697e-06, 
    4.713392e-06, 4.743419e-06, 4.441834e-06, 4.459606e-06, 4.458037e-06, 
    4.476672e-06, 4.490483e-06, 4.520497e-06, 4.568878e-06, 4.550649e-06, 
    4.584143e-06, 4.590885e-06, 4.540011e-06, 4.571211e-06, 4.47152e-06, 
    4.487544e-06, 4.477997e-06, 4.443236e-06, 4.55485e-06, 4.497374e-06, 
    4.60383e-06, 4.57245e-06, 4.664375e-06, 4.618531e-06, 4.708825e-06, 
    4.74774e-06, 4.784519e-06, 4.827724e-06, 4.469319e-06, 4.457224e-06, 
    4.47889e-06, 4.50897e-06, 4.536974e-06, 4.574361e-06, 4.578195e-06, 
    4.585223e-06, 4.603452e-06, 4.618812e-06, 4.587449e-06, 4.622667e-06, 
    4.491271e-06, 4.559857e-06, 4.452659e-06, 4.48479e-06, 4.507192e-06, 
    4.497354e-06, 4.548568e-06, 4.560687e-06, 4.610127e-06, 4.58453e-06, 
    4.73812e-06, 4.66981e-06, 4.860762e-06, 4.806956e-06, 4.453004e-06, 
    4.469276e-06, 4.526175e-06, 4.499051e-06, 4.576862e-06, 4.596133e-06, 
    4.611831e-06, 4.631946e-06, 4.634119e-06, 4.646064e-06, 4.6265e-06, 
    4.645289e-06, 4.574441e-06, 4.606024e-06, 4.519647e-06, 4.540586e-06, 
    4.530946e-06, 4.520386e-06, 4.553021e-06, 4.587942e-06, 4.588685e-06, 
    4.599917e-06, 4.63166e-06, 4.577179e-06, 4.746988e-06, 4.641707e-06, 
    4.487058e-06, 4.518573e-06, 4.523079e-06, 4.51085e-06, 4.594199e-06, 
    4.563899e-06, 4.645772e-06, 4.623561e-06, 4.659983e-06, 4.641865e-06, 
    4.639202e-06, 4.615997e-06, 4.601585e-06, 4.565286e-06, 4.535872e-06, 
    4.512622e-06, 4.518022e-06, 4.543582e-06, 4.590082e-06, 4.634318e-06, 
    4.624608e-06, 4.65721e-06, 4.571194e-06, 4.607153e-06, 4.593237e-06, 
    4.629571e-06, 4.550167e-06, 4.617749e-06, 4.532985e-06, 4.54038e-06, 
    4.563298e-06, 4.609601e-06, 4.619874e-06, 4.630866e-06, 4.624081e-06, 
    4.591265e-06, 4.5859e-06, 4.562739e-06, 4.556359e-06, 4.538769e-06, 
    4.524237e-06, 4.537514e-06, 4.551482e-06, 4.591277e-06, 4.627312e-06, 
    4.666782e-06, 4.676469e-06, 4.722896e-06, 4.685089e-06, 4.747579e-06, 
    4.69443e-06, 4.786647e-06, 4.621676e-06, 4.692863e-06, 4.564341e-06, 
    4.578088e-06, 4.603017e-06, 4.660476e-06, 4.6294e-06, 4.665753e-06, 
    4.58569e-06, 4.544468e-06, 4.533832e-06, 4.514034e-06, 4.534285e-06, 
    4.532636e-06, 4.552058e-06, 4.545811e-06, 4.592602e-06, 4.567434e-06, 
    4.639137e-06, 4.665464e-06, 4.740268e-06, 4.786468e-06, 4.833754e-06, 
    4.854718e-06, 4.861109e-06, 4.863782e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWDP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWLIQ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_DEPTH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SINKS =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 SNOW_SOURCES =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 SOIL1C =
  5.777963, 5.777942, 5.777946, 5.77793, 5.777939, 5.777928, 5.777958, 
    5.777942, 5.777952, 5.777961, 5.777898, 5.777929, 5.777866, 5.777886, 
    5.777836, 5.777869, 5.77783, 5.777837, 5.777815, 5.777821, 5.777792, 
    5.777812, 5.777777, 5.777797, 5.777794, 5.777812, 5.777923, 5.777902, 
    5.777924, 5.777921, 5.777923, 5.777939, 5.777947, 5.777964, 5.777961, 
    5.777948, 5.77792, 5.77793, 5.777905, 5.777906, 5.777879, 5.777891, 
    5.777845, 5.777858, 5.777821, 5.777831, 5.777822, 5.777824, 5.777822, 
    5.777835, 5.777829, 5.777842, 5.777889, 5.777875, 5.777916, 5.777941, 
    5.777958, 5.777969, 5.777968, 5.777965, 5.777948, 5.777933, 5.777921, 
    5.777914, 5.777906, 5.777883, 5.77787, 5.777843, 5.777848, 5.777839, 
    5.777832, 5.777818, 5.77782, 5.777814, 5.77784, 5.777822, 5.777851, 
    5.777843, 5.777904, 5.777927, 5.777937, 5.777946, 5.777966, 5.777952, 
    5.777958, 5.777944, 5.777936, 5.77794, 5.777914, 5.777924, 5.77787, 
    5.777893, 5.777832, 5.777847, 5.777829, 5.777838, 5.777822, 5.777836, 
    5.777812, 5.777807, 5.77781, 5.777796, 5.777837, 5.777822, 5.77794, 
    5.777939, 5.777936, 5.77795, 5.777951, 5.777964, 5.777953, 5.777947, 
    5.777935, 5.777927, 5.77792, 5.777905, 5.777887, 5.777864, 5.777846, 
    5.777834, 5.777841, 5.777835, 5.777842, 5.777845, 5.777809, 5.777829, 
    5.777798, 5.7778, 5.777814, 5.7778, 5.777939, 5.777943, 5.777956, 
    5.777946, 5.777966, 5.777955, 5.777948, 5.777924, 5.777918, 5.777913, 
    5.777903, 5.77789, 5.777868, 5.777849, 5.777831, 5.777832, 5.777832, 
    5.777828, 5.777838, 5.777826, 5.777824, 5.777829, 5.7778, 5.777809, 
    5.7778, 5.777805, 5.777941, 5.777935, 5.777938, 5.777931, 5.777936, 
    5.777915, 5.777908, 5.777878, 5.777891, 5.777871, 5.777889, 5.777885, 
    5.77787, 5.777888, 5.77785, 5.777875, 5.777828, 5.777853, 5.777826, 
    5.777831, 5.777822, 5.777815, 5.777806, 5.777789, 5.777793, 5.777779, 
    5.777925, 5.777916, 5.777916, 5.777907, 5.777901, 5.777886, 5.777863, 
    5.777871, 5.777855, 5.777852, 5.777876, 5.777861, 5.77791, 5.777902, 
    5.777907, 5.777924, 5.777869, 5.777897, 5.777845, 5.777861, 5.777816, 
    5.777838, 5.777795, 5.777777, 5.777759, 5.777739, 5.777911, 5.777917, 
    5.777906, 5.777892, 5.777878, 5.77786, 5.777858, 5.777854, 5.777846, 
    5.777838, 5.777853, 5.777836, 5.7779, 5.777867, 5.777919, 5.777904, 
    5.777893, 5.777897, 5.777872, 5.777866, 5.777843, 5.777855, 5.777781, 
    5.777814, 5.777723, 5.777749, 5.777919, 5.777911, 5.777883, 5.777896, 
    5.777859, 5.777849, 5.777842, 5.777832, 5.777831, 5.777825, 5.777834, 
    5.777825, 5.77786, 5.777844, 5.777886, 5.777876, 5.777881, 5.777886, 
    5.77787, 5.777853, 5.777853, 5.777847, 5.777832, 5.777858, 5.777777, 
    5.777827, 5.777902, 5.777887, 5.777885, 5.777891, 5.77785, 5.777865, 
    5.777825, 5.777836, 5.777819, 5.777827, 5.777829, 5.77784, 5.777847, 
    5.777864, 5.777878, 5.77789, 5.777887, 5.777875, 5.777852, 5.777831, 
    5.777835, 5.77782, 5.777861, 5.777844, 5.777851, 5.777833, 5.777872, 
    5.777839, 5.77788, 5.777876, 5.777865, 5.777843, 5.777838, 5.777833, 
    5.777836, 5.777852, 5.777854, 5.777865, 5.777869, 5.777877, 5.777884, 
    5.777878, 5.777871, 5.777852, 5.777834, 5.777815, 5.777811, 5.777789, 
    5.777806, 5.777777, 5.777802, 5.777758, 5.777837, 5.777803, 5.777864, 
    5.777858, 5.777846, 5.777818, 5.777833, 5.777816, 5.777854, 5.777874, 
    5.77788, 5.777889, 5.777879, 5.77788, 5.777871, 5.777874, 5.777851, 
    5.777863, 5.777829, 5.777816, 5.77778, 5.777759, 5.777736, 5.777726, 
    5.777723, 5.777722 ;

 SOIL1C_TO_SOIL2C =
  3.18083e-08, 3.194808e-08, 3.192091e-08, 3.203365e-08, 3.197111e-08, 
    3.204494e-08, 3.183664e-08, 3.195364e-08, 3.187895e-08, 3.182088e-08, 
    3.225245e-08, 3.203868e-08, 3.247448e-08, 3.233815e-08, 3.26806e-08, 
    3.245327e-08, 3.272643e-08, 3.267403e-08, 3.283173e-08, 3.278655e-08, 
    3.298826e-08, 3.285258e-08, 3.309281e-08, 3.295585e-08, 3.297728e-08, 
    3.28481e-08, 3.20817e-08, 3.222584e-08, 3.207316e-08, 3.209372e-08, 
    3.208449e-08, 3.197241e-08, 3.191592e-08, 3.179761e-08, 3.181909e-08, 
    3.190598e-08, 3.210296e-08, 3.203609e-08, 3.22046e-08, 3.22008e-08, 
    3.238839e-08, 3.230381e-08, 3.261911e-08, 3.25295e-08, 3.278844e-08, 
    3.272332e-08, 3.278538e-08, 3.276656e-08, 3.278562e-08, 3.269012e-08, 
    3.273104e-08, 3.264699e-08, 3.231965e-08, 3.241586e-08, 3.212892e-08, 
    3.195638e-08, 3.184177e-08, 3.176044e-08, 3.177194e-08, 3.179386e-08, 
    3.190649e-08, 3.201238e-08, 3.209308e-08, 3.214706e-08, 3.220025e-08, 
    3.236125e-08, 3.244645e-08, 3.263723e-08, 3.26028e-08, 3.266112e-08, 
    3.271684e-08, 3.281039e-08, 3.279499e-08, 3.28362e-08, 3.265958e-08, 
    3.277697e-08, 3.258318e-08, 3.263618e-08, 3.221473e-08, 3.205413e-08, 
    3.198588e-08, 3.192613e-08, 3.178078e-08, 3.188116e-08, 3.184159e-08, 
    3.193573e-08, 3.199554e-08, 3.196596e-08, 3.214854e-08, 3.207756e-08, 
    3.24515e-08, 3.229043e-08, 3.271034e-08, 3.260986e-08, 3.273442e-08, 
    3.267086e-08, 3.277977e-08, 3.268175e-08, 3.285154e-08, 3.288851e-08, 
    3.286325e-08, 3.296029e-08, 3.267632e-08, 3.278538e-08, 3.196513e-08, 
    3.196995e-08, 3.199243e-08, 3.189362e-08, 3.188758e-08, 3.179703e-08, 
    3.18776e-08, 3.191191e-08, 3.199901e-08, 3.205053e-08, 3.20995e-08, 
    3.220718e-08, 3.232743e-08, 3.249558e-08, 3.261637e-08, 3.269735e-08, 
    3.264769e-08, 3.269153e-08, 3.264253e-08, 3.261956e-08, 3.287466e-08, 
    3.273142e-08, 3.294634e-08, 3.293444e-08, 3.283718e-08, 3.293578e-08, 
    3.197334e-08, 3.194558e-08, 3.184918e-08, 3.192462e-08, 3.178716e-08, 
    3.18641e-08, 3.190835e-08, 3.207904e-08, 3.211654e-08, 3.215132e-08, 
    3.222e-08, 3.230814e-08, 3.246276e-08, 3.259728e-08, 3.272008e-08, 
    3.271108e-08, 3.271425e-08, 3.274168e-08, 3.267373e-08, 3.275284e-08, 
    3.276612e-08, 3.27314e-08, 3.293285e-08, 3.28753e-08, 3.293419e-08, 
    3.289672e-08, 3.19546e-08, 3.200132e-08, 3.197608e-08, 3.202355e-08, 
    3.19901e-08, 3.213882e-08, 3.218341e-08, 3.239203e-08, 3.230641e-08, 
    3.244267e-08, 3.232025e-08, 3.234194e-08, 3.244712e-08, 3.232686e-08, 
    3.258987e-08, 3.241157e-08, 3.274275e-08, 3.256471e-08, 3.275391e-08, 
    3.271955e-08, 3.277643e-08, 3.282738e-08, 3.289147e-08, 3.300973e-08, 
    3.298235e-08, 3.308125e-08, 3.207097e-08, 3.213157e-08, 3.212623e-08, 
    3.218964e-08, 3.223654e-08, 3.233819e-08, 3.250121e-08, 3.243991e-08, 
    3.255245e-08, 3.257504e-08, 3.240406e-08, 3.250904e-08, 3.217212e-08, 
    3.222656e-08, 3.219414e-08, 3.207575e-08, 3.245404e-08, 3.22599e-08, 
    3.261837e-08, 3.251321e-08, 3.282012e-08, 3.266749e-08, 3.296728e-08, 
    3.309543e-08, 3.321603e-08, 3.335698e-08, 3.216464e-08, 3.212346e-08, 
    3.219719e-08, 3.229919e-08, 3.239382e-08, 3.251963e-08, 3.253249e-08, 
    3.255607e-08, 3.261711e-08, 3.266844e-08, 3.256352e-08, 3.268131e-08, 
    3.223919e-08, 3.247089e-08, 3.21079e-08, 3.221721e-08, 3.229317e-08, 
    3.225985e-08, 3.24329e-08, 3.247369e-08, 3.263942e-08, 3.255375e-08, 
    3.306381e-08, 3.283814e-08, 3.346429e-08, 3.328932e-08, 3.210908e-08, 
    3.216449e-08, 3.235736e-08, 3.22656e-08, 3.252802e-08, 3.259262e-08, 
    3.264512e-08, 3.271225e-08, 3.271949e-08, 3.275926e-08, 3.269409e-08, 
    3.275669e-08, 3.251989e-08, 3.262571e-08, 3.233531e-08, 3.2406e-08, 
    3.237348e-08, 3.233781e-08, 3.244789e-08, 3.256517e-08, 3.256767e-08, 
    3.260528e-08, 3.271126e-08, 3.252908e-08, 3.309294e-08, 3.274473e-08, 
    3.222492e-08, 3.233167e-08, 3.234691e-08, 3.230556e-08, 3.258614e-08, 
    3.248448e-08, 3.275829e-08, 3.268429e-08, 3.280554e-08, 3.274529e-08, 
    3.273643e-08, 3.265904e-08, 3.261086e-08, 3.248914e-08, 3.23901e-08, 
    3.231156e-08, 3.232982e-08, 3.24161e-08, 3.257234e-08, 3.272015e-08, 
    3.268777e-08, 3.279633e-08, 3.2509e-08, 3.262948e-08, 3.258291e-08, 
    3.270434e-08, 3.243828e-08, 3.266485e-08, 3.238036e-08, 3.240531e-08, 
    3.248246e-08, 3.263766e-08, 3.267198e-08, 3.270865e-08, 3.268602e-08, 
    3.257631e-08, 3.255833e-08, 3.248059e-08, 3.245912e-08, 3.239987e-08, 
    3.235083e-08, 3.239564e-08, 3.244271e-08, 3.257635e-08, 3.26968e-08, 
    3.282811e-08, 3.286024e-08, 3.301367e-08, 3.288878e-08, 3.309488e-08, 
    3.291967e-08, 3.322296e-08, 3.267798e-08, 3.29145e-08, 3.248597e-08, 
    3.253214e-08, 3.261565e-08, 3.280716e-08, 3.270376e-08, 3.282468e-08, 
    3.255763e-08, 3.241907e-08, 3.238322e-08, 3.231633e-08, 3.238475e-08, 
    3.237918e-08, 3.244465e-08, 3.242361e-08, 3.258079e-08, 3.249636e-08, 
    3.27362e-08, 3.282373e-08, 3.307088e-08, 3.32224e-08, 3.337661e-08, 
    3.34447e-08, 3.346542e-08, 3.347408e-08 ;

 SOIL1C_TO_SOIL3C =
  3.772561e-10, 3.789146e-10, 3.785922e-10, 3.799299e-10, 3.791878e-10, 
    3.800637e-10, 3.775923e-10, 3.789805e-10, 3.780943e-10, 3.774054e-10, 
    3.825259e-10, 3.799895e-10, 3.851602e-10, 3.835427e-10, 3.876058e-10, 
    3.849085e-10, 3.881497e-10, 3.87528e-10, 3.893991e-10, 3.88863e-10, 
    3.912564e-10, 3.896465e-10, 3.924969e-10, 3.908719e-10, 3.911261e-10, 
    3.895934e-10, 3.804999e-10, 3.822101e-10, 3.803986e-10, 3.806425e-10, 
    3.80533e-10, 3.792031e-10, 3.78533e-10, 3.771293e-10, 3.773841e-10, 
    3.784151e-10, 3.807521e-10, 3.799588e-10, 3.819581e-10, 3.81913e-10, 
    3.841388e-10, 3.831352e-10, 3.868762e-10, 3.85813e-10, 3.888854e-10, 
    3.881127e-10, 3.888491e-10, 3.886258e-10, 3.88852e-10, 3.877188e-10, 
    3.882043e-10, 3.872072e-10, 3.833232e-10, 3.844647e-10, 3.810602e-10, 
    3.79013e-10, 3.776532e-10, 3.766883e-10, 3.768247e-10, 3.770848e-10, 
    3.784211e-10, 3.796775e-10, 3.806349e-10, 3.812754e-10, 3.819065e-10, 
    3.838167e-10, 3.848276e-10, 3.870912e-10, 3.866827e-10, 3.873748e-10, 
    3.880359e-10, 3.891458e-10, 3.889631e-10, 3.894522e-10, 3.873565e-10, 
    3.887493e-10, 3.8645e-10, 3.870789e-10, 3.820782e-10, 3.801728e-10, 
    3.79363e-10, 3.786541e-10, 3.769296e-10, 3.781205e-10, 3.77651e-10, 
    3.787679e-10, 3.794776e-10, 3.791266e-10, 3.812929e-10, 3.804508e-10, 
    3.848876e-10, 3.829765e-10, 3.879587e-10, 3.867665e-10, 3.882445e-10, 
    3.874903e-10, 3.887826e-10, 3.876195e-10, 3.896342e-10, 3.900728e-10, 
    3.897731e-10, 3.909246e-10, 3.875551e-10, 3.888491e-10, 3.791168e-10, 
    3.791741e-10, 3.794408e-10, 3.782684e-10, 3.781967e-10, 3.771223e-10, 
    3.780783e-10, 3.784854e-10, 3.795188e-10, 3.8013e-10, 3.807111e-10, 
    3.819887e-10, 3.834155e-10, 3.854106e-10, 3.868438e-10, 3.878046e-10, 
    3.872154e-10, 3.877356e-10, 3.871541e-10, 3.868816e-10, 3.899085e-10, 
    3.882089e-10, 3.90759e-10, 3.906178e-10, 3.894638e-10, 3.906337e-10, 
    3.792142e-10, 3.788848e-10, 3.777411e-10, 3.786362e-10, 3.770053e-10, 
    3.779182e-10, 3.784431e-10, 3.804684e-10, 3.809133e-10, 3.813259e-10, 
    3.821408e-10, 3.831866e-10, 3.850211e-10, 3.866173e-10, 3.880743e-10, 
    3.879675e-10, 3.880051e-10, 3.883306e-10, 3.875244e-10, 3.88463e-10, 
    3.886206e-10, 3.882087e-10, 3.905989e-10, 3.89916e-10, 3.906148e-10, 
    3.901702e-10, 3.789919e-10, 3.795462e-10, 3.792467e-10, 3.7981e-10, 
    3.794131e-10, 3.811776e-10, 3.817066e-10, 3.841819e-10, 3.83166e-10, 
    3.847828e-10, 3.833302e-10, 3.835876e-10, 3.848356e-10, 3.834087e-10, 
    3.865293e-10, 3.844137e-10, 3.883433e-10, 3.862308e-10, 3.884757e-10, 
    3.88068e-10, 3.88743e-10, 3.893475e-10, 3.90108e-10, 3.915112e-10, 
    3.911863e-10, 3.923598e-10, 3.803726e-10, 3.810916e-10, 3.810282e-10, 
    3.817806e-10, 3.823371e-10, 3.835431e-10, 3.854774e-10, 3.8475e-10, 
    3.860853e-10, 3.863534e-10, 3.843247e-10, 3.855703e-10, 3.815727e-10, 
    3.822186e-10, 3.81834e-10, 3.804293e-10, 3.849177e-10, 3.826143e-10, 
    3.868675e-10, 3.856198e-10, 3.892613e-10, 3.874503e-10, 3.910074e-10, 
    3.925281e-10, 3.939591e-10, 3.956316e-10, 3.814839e-10, 3.809954e-10, 
    3.818701e-10, 3.830803e-10, 3.842031e-10, 3.856959e-10, 3.858486e-10, 
    3.861282e-10, 3.868525e-10, 3.874616e-10, 3.862167e-10, 3.876142e-10, 
    3.823685e-10, 3.851176e-10, 3.808107e-10, 3.821077e-10, 3.83009e-10, 
    3.826136e-10, 3.846669e-10, 3.851508e-10, 3.871173e-10, 3.861007e-10, 
    3.921528e-10, 3.894752e-10, 3.969049e-10, 3.948287e-10, 3.808247e-10, 
    3.814822e-10, 3.837706e-10, 3.826818e-10, 3.857955e-10, 3.865619e-10, 
    3.871849e-10, 3.879814e-10, 3.880674e-10, 3.885392e-10, 3.87766e-10, 
    3.885087e-10, 3.856991e-10, 3.869546e-10, 3.83509e-10, 3.843477e-10, 
    3.839619e-10, 3.835387e-10, 3.848448e-10, 3.862363e-10, 3.86266e-10, 
    3.867122e-10, 3.879696e-10, 3.858081e-10, 3.924985e-10, 3.883668e-10, 
    3.821992e-10, 3.834657e-10, 3.836466e-10, 3.83156e-10, 3.864851e-10, 
    3.852788e-10, 3.885277e-10, 3.876497e-10, 3.890883e-10, 3.883734e-10, 
    3.882683e-10, 3.873501e-10, 3.867784e-10, 3.853342e-10, 3.84159e-10, 
    3.832271e-10, 3.834438e-10, 3.844675e-10, 3.863214e-10, 3.880752e-10, 
    3.87691e-10, 3.88979e-10, 3.855697e-10, 3.869993e-10, 3.864468e-10, 
    3.878875e-10, 3.847307e-10, 3.87419e-10, 3.840435e-10, 3.843394e-10, 
    3.852549e-10, 3.870964e-10, 3.875037e-10, 3.879387e-10, 3.876702e-10, 
    3.863684e-10, 3.861552e-10, 3.852327e-10, 3.84978e-10, 3.84275e-10, 
    3.83693e-10, 3.842248e-10, 3.847832e-10, 3.86369e-10, 3.87798e-10, 
    3.893561e-10, 3.897374e-10, 3.915579e-10, 3.90076e-10, 3.925215e-10, 
    3.904425e-10, 3.940413e-10, 3.875748e-10, 3.903812e-10, 3.852965e-10, 
    3.858443e-10, 3.868351e-10, 3.891076e-10, 3.878807e-10, 3.893155e-10, 
    3.861468e-10, 3.845028e-10, 3.840774e-10, 3.832838e-10, 3.840955e-10, 
    3.840295e-10, 3.848063e-10, 3.845567e-10, 3.864216e-10, 3.854199e-10, 
    3.882656e-10, 3.893041e-10, 3.922368e-10, 3.940346e-10, 3.958645e-10, 
    3.966724e-10, 3.969183e-10, 3.970211e-10 ;

 SOIL1C_vr =
  19.9794, 19.97934, 19.97935, 19.97931, 19.97933, 19.97931, 19.97939, 
    19.97934, 19.97937, 19.97939, 19.97923, 19.97931, 19.97914, 19.97919, 
    19.97906, 19.97915, 19.97904, 19.97906, 19.979, 19.97902, 19.97894, 
    19.979, 19.9789, 19.97896, 19.97895, 19.979, 19.97929, 19.97924, 19.9793, 
    19.97929, 19.97929, 19.97933, 19.97935, 19.9794, 19.97939, 19.97936, 
    19.97928, 19.97931, 19.97924, 19.97925, 19.97917, 19.97921, 19.97909, 
    19.97912, 19.97902, 19.97905, 19.97902, 19.97903, 19.97902, 19.97906, 
    19.97904, 19.97907, 19.9792, 19.97916, 19.97927, 19.97934, 19.97938, 
    19.97942, 19.97941, 19.9794, 19.97936, 19.97932, 19.97929, 19.97927, 
    19.97925, 19.97919, 19.97915, 19.97908, 19.97909, 19.97907, 19.97905, 
    19.97901, 19.97902, 19.979, 19.97907, 19.97902, 19.9791, 19.97908, 
    19.97924, 19.9793, 19.97933, 19.97935, 19.97941, 19.97937, 19.97938, 
    19.97935, 19.97932, 19.97934, 19.97927, 19.97929, 19.97915, 19.97921, 
    19.97905, 19.97909, 19.97904, 19.97906, 19.97902, 19.97906, 19.979, 
    19.97898, 19.97899, 19.97895, 19.97906, 19.97902, 19.97934, 19.97934, 
    19.97933, 19.97936, 19.97937, 19.9794, 19.97937, 19.97936, 19.97932, 
    19.9793, 19.97928, 19.97924, 19.9792, 19.97913, 19.97909, 19.97906, 
    19.97907, 19.97906, 19.97908, 19.97909, 19.97899, 19.97904, 19.97896, 
    19.97896, 19.979, 19.97896, 19.97933, 19.97934, 19.97938, 19.97935, 
    19.97941, 19.97938, 19.97936, 19.97929, 19.97928, 19.97927, 19.97924, 
    19.9792, 19.97915, 19.97909, 19.97905, 19.97905, 19.97905, 19.97904, 
    19.97906, 19.97903, 19.97903, 19.97904, 19.97897, 19.97899, 19.97897, 
    19.97898, 19.97934, 19.97932, 19.97933, 19.97931, 19.97933, 19.97927, 
    19.97925, 19.97917, 19.97921, 19.97915, 19.9792, 19.97919, 19.97915, 
    19.9792, 19.9791, 19.97916, 19.97904, 19.97911, 19.97903, 19.97905, 
    19.97902, 19.97901, 19.97898, 19.97894, 19.97895, 19.97891, 19.9793, 
    19.97927, 19.97927, 19.97925, 19.97923, 19.97919, 19.97913, 19.97915, 
    19.97911, 19.9791, 19.97917, 19.97913, 19.97926, 19.97924, 19.97925, 
    19.97929, 19.97915, 19.97922, 19.97909, 19.97913, 19.97901, 19.97907, 
    19.97895, 19.9789, 19.97886, 19.9788, 19.97926, 19.97928, 19.97925, 
    19.97921, 19.97917, 19.97912, 19.97912, 19.97911, 19.97909, 19.97907, 
    19.97911, 19.97906, 19.97923, 19.97914, 19.97928, 19.97924, 19.97921, 
    19.97922, 19.97916, 19.97914, 19.97908, 19.97911, 19.97892, 19.979, 
    19.97876, 19.97883, 19.97928, 19.97926, 19.97919, 19.97922, 19.97912, 
    19.9791, 19.97907, 19.97905, 19.97905, 19.97903, 19.97906, 19.97903, 
    19.97912, 19.97908, 19.97919, 19.97917, 19.97918, 19.97919, 19.97915, 
    19.97911, 19.9791, 19.97909, 19.97905, 19.97912, 19.9789, 19.97904, 
    19.97924, 19.9792, 19.97919, 19.97921, 19.9791, 19.97914, 19.97903, 
    19.97906, 19.97901, 19.97904, 19.97904, 19.97907, 19.97909, 19.97914, 
    19.97917, 19.9792, 19.9792, 19.97916, 19.9791, 19.97905, 19.97906, 
    19.97902, 19.97913, 19.97908, 19.9791, 19.97905, 19.97915, 19.97907, 
    19.97918, 19.97917, 19.97914, 19.97908, 19.97906, 19.97905, 19.97906, 
    19.9791, 19.97911, 19.97914, 19.97915, 19.97917, 19.97919, 19.97917, 
    19.97915, 19.9791, 19.97906, 19.97901, 19.97899, 19.97894, 19.97898, 
    19.9789, 19.97897, 19.97886, 19.97906, 19.97897, 19.97914, 19.97912, 
    19.97909, 19.97901, 19.97905, 19.97901, 19.97911, 19.97916, 19.97918, 
    19.9792, 19.97918, 19.97918, 19.97915, 19.97916, 19.9791, 19.97913, 
    19.97904, 19.97901, 19.97891, 19.97886, 19.9788, 19.97877, 19.97876, 
    19.97876,
  19.981, 19.98093, 19.98094, 19.98088, 19.98092, 19.98088, 19.98099, 
    19.98093, 19.98096, 19.98099, 19.98077, 19.98088, 19.98066, 19.98073, 
    19.98056, 19.98067, 19.98053, 19.98056, 19.98048, 19.9805, 19.9804, 
    19.98047, 19.98035, 19.98042, 19.98041, 19.98047, 19.98086, 19.98079, 
    19.98087, 19.98085, 19.98086, 19.98092, 19.98095, 19.981, 19.98099, 
    19.98095, 19.98085, 19.98088, 19.9808, 19.9808, 19.98071, 19.98075, 
    19.98059, 19.98063, 19.9805, 19.98054, 19.9805, 19.98051, 19.9805, 
    19.98055, 19.98053, 19.98057, 19.98074, 19.98069, 19.98084, 19.98092, 
    19.98098, 19.98102, 19.98102, 19.98101, 19.98095, 19.9809, 19.98085, 
    19.98083, 19.9808, 19.98072, 19.98068, 19.98058, 19.9806, 19.98057, 
    19.98054, 19.98049, 19.9805, 19.98048, 19.98057, 19.98051, 19.98061, 
    19.98058, 19.98079, 19.98088, 19.98091, 19.98094, 19.98101, 19.98096, 
    19.98098, 19.98093, 19.9809, 19.98092, 19.98083, 19.98086, 19.98067, 
    19.98075, 19.98054, 19.98059, 19.98053, 19.98056, 19.98051, 19.98056, 
    19.98047, 19.98045, 19.98046, 19.98042, 19.98056, 19.9805, 19.98092, 
    19.98092, 19.98091, 19.98096, 19.98096, 19.981, 19.98096, 19.98095, 
    19.9809, 19.98088, 19.98085, 19.9808, 19.98074, 19.98065, 19.98059, 
    19.98055, 19.98057, 19.98055, 19.98058, 19.98059, 19.98046, 19.98053, 
    19.98042, 19.98043, 19.98048, 19.98043, 19.98092, 19.98093, 19.98098, 
    19.98094, 19.98101, 19.98097, 19.98095, 19.98086, 19.98084, 19.98083, 
    19.98079, 19.98075, 19.98067, 19.9806, 19.98054, 19.98054, 19.98054, 
    19.98053, 19.98056, 19.98052, 19.98051, 19.98053, 19.98043, 19.98046, 
    19.98043, 19.98045, 19.98092, 19.9809, 19.98092, 19.98089, 19.98091, 
    19.98083, 19.98081, 19.9807, 19.98075, 19.98068, 19.98074, 19.98073, 
    19.98067, 19.98074, 19.9806, 19.98069, 19.98053, 19.98062, 19.98052, 
    19.98054, 19.98051, 19.98048, 19.98045, 19.98039, 19.98041, 19.98036, 
    19.98087, 19.98083, 19.98084, 19.98081, 19.98078, 19.98073, 19.98065, 
    19.98068, 19.98062, 19.98061, 19.9807, 19.98064, 19.98081, 19.98079, 
    19.9808, 19.98086, 19.98067, 19.98077, 19.98059, 19.98064, 19.98049, 
    19.98056, 19.98041, 19.98035, 19.98029, 19.98022, 19.98082, 19.98084, 
    19.9808, 19.98075, 19.9807, 19.98064, 19.98063, 19.98062, 19.98059, 
    19.98056, 19.98062, 19.98056, 19.98078, 19.98066, 19.98085, 19.98079, 
    19.98075, 19.98077, 19.98068, 19.98066, 19.98058, 19.98062, 19.98036, 
    19.98048, 19.98016, 19.98025, 19.98085, 19.98082, 19.98072, 19.98077, 
    19.98063, 19.9806, 19.98058, 19.98054, 19.98054, 19.98052, 19.98055, 
    19.98052, 19.98064, 19.98059, 19.98073, 19.9807, 19.98071, 19.98073, 
    19.98067, 19.98062, 19.98061, 19.98059, 19.98054, 19.98063, 19.98035, 
    19.98053, 19.98079, 19.98073, 19.98073, 19.98075, 19.98061, 19.98066, 
    19.98052, 19.98056, 19.98049, 19.98052, 19.98053, 19.98057, 19.98059, 
    19.98065, 19.98071, 19.98074, 19.98074, 19.98069, 19.98061, 19.98054, 
    19.98055, 19.9805, 19.98064, 19.98058, 19.98061, 19.98055, 19.98068, 
    19.98057, 19.98071, 19.9807, 19.98066, 19.98058, 19.98056, 19.98054, 
    19.98055, 19.98061, 19.98062, 19.98066, 19.98067, 19.9807, 19.98072, 
    19.9807, 19.98068, 19.98061, 19.98055, 19.98048, 19.98047, 19.98039, 
    19.98045, 19.98035, 19.98044, 19.98028, 19.98056, 19.98044, 19.98066, 
    19.98063, 19.98059, 19.98049, 19.98055, 19.98048, 19.98062, 19.98069, 
    19.98071, 19.98074, 19.98071, 19.98071, 19.98068, 19.98069, 19.98061, 
    19.98065, 19.98053, 19.98049, 19.98036, 19.98028, 19.98021, 19.98017, 
    19.98016, 19.98016,
  19.98272, 19.98265, 19.98266, 19.9826, 19.98263, 19.98259, 19.98271, 
    19.98264, 19.98268, 19.98272, 19.98248, 19.9826, 19.98236, 19.98244, 
    19.98225, 19.98237, 19.98223, 19.98225, 19.98217, 19.98219, 19.98208, 
    19.98216, 19.98203, 19.9821, 19.98209, 19.98216, 19.98257, 19.9825, 
    19.98258, 19.98257, 19.98257, 19.98263, 19.98266, 19.98273, 19.98272, 
    19.98267, 19.98256, 19.9826, 19.98251, 19.98251, 19.98241, 19.98245, 
    19.98228, 19.98233, 19.98219, 19.98223, 19.98219, 19.9822, 19.98219, 
    19.98224, 19.98222, 19.98227, 19.98244, 19.98239, 19.98255, 19.98264, 
    19.9827, 19.98275, 19.98274, 19.98273, 19.98267, 19.98261, 19.98257, 
    19.98254, 19.98251, 19.98242, 19.98238, 19.98227, 19.98229, 19.98226, 
    19.98223, 19.98218, 19.98219, 19.98217, 19.98226, 19.9822, 19.9823, 
    19.98228, 19.9825, 19.98259, 19.98263, 19.98266, 19.98274, 19.98268, 
    19.9827, 19.98265, 19.98262, 19.98264, 19.98254, 19.98258, 19.98237, 
    19.98246, 19.98223, 19.98229, 19.98222, 19.98226, 19.9822, 19.98225, 
    19.98216, 19.98214, 19.98215, 19.9821, 19.98225, 19.98219, 19.98264, 
    19.98264, 19.98262, 19.98268, 19.98268, 19.98273, 19.98269, 19.98267, 
    19.98262, 19.98259, 19.98256, 19.98251, 19.98244, 19.98235, 19.98228, 
    19.98224, 19.98227, 19.98224, 19.98227, 19.98228, 19.98215, 19.98222, 
    19.98211, 19.98211, 19.98217, 19.98211, 19.98263, 19.98265, 19.9827, 
    19.98266, 19.98273, 19.98269, 19.98267, 19.98258, 19.98256, 19.98254, 
    19.9825, 19.98245, 19.98237, 19.9823, 19.98223, 19.98223, 19.98223, 
    19.98222, 19.98225, 19.98221, 19.9822, 19.98222, 19.98211, 19.98215, 
    19.98211, 19.98213, 19.98264, 19.98262, 19.98263, 19.9826, 19.98262, 
    19.98254, 19.98252, 19.98241, 19.98245, 19.98238, 19.98244, 19.98243, 
    19.98238, 19.98244, 19.9823, 19.9824, 19.98222, 19.98231, 19.98221, 
    19.98223, 19.9822, 19.98217, 19.98214, 19.98207, 19.98209, 19.98203, 
    19.98258, 19.98255, 19.98255, 19.98252, 19.98249, 19.98244, 19.98235, 
    19.98238, 19.98232, 19.98231, 19.9824, 19.98234, 19.98252, 19.9825, 
    19.98251, 19.98258, 19.98237, 19.98248, 19.98228, 19.98234, 19.98218, 
    19.98226, 19.9821, 19.98203, 19.98196, 19.98189, 19.98253, 19.98255, 
    19.98251, 19.98246, 19.9824, 19.98234, 19.98233, 19.98232, 19.98228, 
    19.98226, 19.98231, 19.98225, 19.98249, 19.98236, 19.98256, 19.9825, 
    19.98246, 19.98248, 19.98238, 19.98236, 19.98227, 19.98232, 19.98204, 
    19.98216, 19.98183, 19.98192, 19.98256, 19.98253, 19.98243, 19.98248, 
    19.98233, 19.9823, 19.98227, 19.98223, 19.98223, 19.98221, 19.98224, 
    19.98221, 19.98234, 19.98228, 19.98244, 19.9824, 19.98242, 19.98244, 
    19.98238, 19.98231, 19.98231, 19.98229, 19.98223, 19.98233, 19.98203, 
    19.98222, 19.9825, 19.98244, 19.98243, 19.98245, 19.9823, 19.98236, 
    19.98221, 19.98225, 19.98218, 19.98222, 19.98222, 19.98226, 19.98229, 
    19.98235, 19.98241, 19.98245, 19.98244, 19.98239, 19.98231, 19.98223, 
    19.98225, 19.98219, 19.98234, 19.98228, 19.9823, 19.98224, 19.98238, 
    19.98226, 19.98241, 19.9824, 19.98236, 19.98227, 19.98225, 19.98223, 
    19.98225, 19.98231, 19.98232, 19.98236, 19.98237, 19.9824, 19.98243, 
    19.9824, 19.98238, 19.98231, 19.98224, 19.98217, 19.98215, 19.98207, 
    19.98214, 19.98203, 19.98212, 19.98196, 19.98225, 19.98212, 19.98236, 
    19.98233, 19.98228, 19.98218, 19.98224, 19.98217, 19.98232, 19.98239, 
    19.98241, 19.98245, 19.98241, 19.98241, 19.98238, 19.98239, 19.9823, 
    19.98235, 19.98222, 19.98217, 19.98204, 19.98196, 19.98187, 19.98184, 
    19.98183, 19.98182,
  19.9841, 19.98402, 19.98404, 19.98398, 19.98401, 19.98397, 19.98408, 
    19.98402, 19.98406, 19.98409, 19.98386, 19.98397, 19.98374, 19.98381, 
    19.98363, 19.98375, 19.98361, 19.98363, 19.98355, 19.98357, 19.98347, 
    19.98354, 19.98341, 19.98348, 19.98347, 19.98354, 19.98395, 19.98388, 
    19.98396, 19.98395, 19.98395, 19.98401, 19.98404, 19.9841, 19.98409, 
    19.98405, 19.98394, 19.98398, 19.98389, 19.98389, 19.98379, 19.98383, 
    19.98366, 19.98371, 19.98357, 19.98361, 19.98357, 19.98359, 19.98357, 
    19.98363, 19.9836, 19.98365, 19.98382, 19.98377, 19.98393, 19.98402, 
    19.98408, 19.98413, 19.98412, 19.98411, 19.98405, 19.98399, 19.98395, 
    19.98392, 19.98389, 19.9838, 19.98376, 19.98365, 19.98367, 19.98364, 
    19.98361, 19.98356, 19.98357, 19.98355, 19.98364, 19.98358, 19.98368, 
    19.98365, 19.98388, 19.98397, 19.984, 19.98404, 19.98411, 19.98406, 
    19.98408, 19.98403, 19.984, 19.98401, 19.98392, 19.98396, 19.98375, 
    19.98384, 19.98362, 19.98367, 19.9836, 19.98364, 19.98358, 19.98363, 
    19.98354, 19.98352, 19.98353, 19.98348, 19.98363, 19.98357, 19.98401, 
    19.98401, 19.984, 19.98405, 19.98406, 19.98411, 19.98406, 19.98404, 
    19.984, 19.98397, 19.98394, 19.98388, 19.98382, 19.98373, 19.98367, 
    19.98362, 19.98365, 19.98363, 19.98365, 19.98366, 19.98353, 19.9836, 
    19.98349, 19.9835, 19.98355, 19.98349, 19.98401, 19.98403, 19.98408, 
    19.98404, 19.98411, 19.98407, 19.98405, 19.98395, 19.98393, 19.98392, 
    19.98388, 19.98383, 19.98375, 19.98368, 19.98361, 19.98361, 19.98361, 
    19.9836, 19.98363, 19.98359, 19.98359, 19.9836, 19.9835, 19.98353, 
    19.9835, 19.98351, 19.98402, 19.984, 19.98401, 19.98398, 19.984, 
    19.98392, 19.9839, 19.98379, 19.98383, 19.98376, 19.98382, 19.98381, 
    19.98376, 19.98382, 19.98368, 19.98378, 19.9836, 19.98369, 19.98359, 
    19.98361, 19.98358, 19.98355, 19.98352, 19.98345, 19.98347, 19.98342, 
    19.98396, 19.98392, 19.98393, 19.98389, 19.98387, 19.98381, 19.98373, 
    19.98376, 19.9837, 19.98369, 19.98378, 19.98372, 19.9839, 19.98388, 
    19.98389, 19.98396, 19.98375, 19.98386, 19.98366, 19.98372, 19.98356, 
    19.98364, 19.98348, 19.98341, 19.98334, 19.98327, 19.98391, 19.98393, 
    19.98389, 19.98384, 19.98379, 19.98372, 19.98371, 19.9837, 19.98367, 
    19.98364, 19.98369, 19.98363, 19.98387, 19.98374, 19.98394, 19.98388, 
    19.98384, 19.98386, 19.98376, 19.98374, 19.98365, 19.9837, 19.98343, 
    19.98355, 19.98321, 19.9833, 19.98394, 19.98391, 19.9838, 19.98385, 
    19.98371, 19.98368, 19.98365, 19.98361, 19.98361, 19.98359, 19.98362, 
    19.98359, 19.98372, 19.98366, 19.98382, 19.98378, 19.9838, 19.98381, 
    19.98376, 19.98369, 19.98369, 19.98367, 19.98361, 19.98371, 19.98341, 
    19.9836, 19.98388, 19.98382, 19.98381, 19.98383, 19.98368, 19.98374, 
    19.98359, 19.98363, 19.98356, 19.9836, 19.9836, 19.98364, 19.98367, 
    19.98373, 19.98379, 19.98383, 19.98382, 19.98377, 19.98369, 19.98361, 
    19.98363, 19.98357, 19.98372, 19.98366, 19.98368, 19.98362, 19.98376, 
    19.98364, 19.98379, 19.98378, 19.98374, 19.98365, 19.98363, 19.98362, 
    19.98363, 19.98369, 19.9837, 19.98374, 19.98375, 19.98378, 19.98381, 
    19.98378, 19.98376, 19.98369, 19.98362, 19.98355, 19.98353, 19.98345, 
    19.98352, 19.98341, 19.9835, 19.98334, 19.98363, 19.98351, 19.98374, 
    19.98371, 19.98367, 19.98356, 19.98362, 19.98355, 19.9837, 19.98377, 
    19.98379, 19.98383, 19.98379, 19.98379, 19.98376, 19.98377, 19.98368, 
    19.98373, 19.9836, 19.98355, 19.98342, 19.98334, 19.98326, 19.98322, 
    19.98321, 19.98321,
  19.9857, 19.98564, 19.98565, 19.9856, 19.98563, 19.98559, 19.98569, 
    19.98564, 19.98567, 19.9857, 19.98549, 19.9856, 19.98539, 19.98545, 
    19.98529, 19.9854, 19.98527, 19.98529, 19.98522, 19.98524, 19.98514, 
    19.98521, 19.98509, 19.98516, 19.98515, 19.98521, 19.98557, 19.98551, 
    19.98558, 19.98557, 19.98557, 19.98563, 19.98565, 19.98571, 19.9857, 
    19.98566, 19.98557, 19.9856, 19.98552, 19.98552, 19.98543, 19.98547, 
    19.98532, 19.98536, 19.98524, 19.98527, 19.98524, 19.98525, 19.98524, 
    19.98528, 19.98527, 19.98531, 19.98546, 19.98542, 19.98555, 19.98563, 
    19.98569, 19.98573, 19.98572, 19.98571, 19.98566, 19.98561, 19.98557, 
    19.98554, 19.98552, 19.98544, 19.9854, 19.98531, 19.98533, 19.9853, 
    19.98527, 19.98523, 19.98524, 19.98521, 19.9853, 19.98524, 19.98534, 
    19.98531, 19.98551, 19.98559, 19.98562, 19.98565, 19.98572, 19.98567, 
    19.98569, 19.98564, 19.98561, 19.98563, 19.98554, 19.98558, 19.9854, 
    19.98548, 19.98528, 19.98532, 19.98526, 19.98529, 19.98524, 19.98529, 
    19.98521, 19.98519, 19.9852, 19.98516, 19.98529, 19.98524, 19.98563, 
    19.98563, 19.98562, 19.98566, 19.98567, 19.98571, 19.98567, 19.98565, 
    19.98561, 19.98559, 19.98557, 19.98552, 19.98546, 19.98538, 19.98532, 
    19.98528, 19.98531, 19.98528, 19.98531, 19.98532, 19.9852, 19.98527, 
    19.98516, 19.98517, 19.98521, 19.98517, 19.98563, 19.98564, 19.98569, 
    19.98565, 19.98571, 19.98568, 19.98566, 19.98558, 19.98556, 19.98554, 
    19.98551, 19.98547, 19.98539, 19.98533, 19.98527, 19.98528, 19.98527, 
    19.98526, 19.98529, 19.98525, 19.98525, 19.98527, 19.98517, 19.9852, 
    19.98517, 19.98519, 19.98564, 19.98561, 19.98562, 19.9856, 19.98562, 
    19.98555, 19.98553, 19.98543, 19.98547, 19.9854, 19.98546, 19.98545, 
    19.9854, 19.98546, 19.98533, 19.98542, 19.98526, 19.98534, 19.98525, 
    19.98527, 19.98524, 19.98522, 19.98519, 19.98513, 19.98515, 19.9851, 
    19.98558, 19.98555, 19.98555, 19.98552, 19.9855, 19.98545, 19.98537, 
    19.9854, 19.98535, 19.98534, 19.98542, 19.98537, 19.98553, 19.98551, 
    19.98552, 19.98558, 19.9854, 19.98549, 19.98532, 19.98537, 19.98522, 
    19.9853, 19.98515, 19.98509, 19.98503, 19.98497, 19.98553, 19.98556, 
    19.98552, 19.98547, 19.98543, 19.98537, 19.98536, 19.98535, 19.98532, 
    19.98529, 19.98535, 19.98529, 19.9855, 19.98539, 19.98556, 19.98551, 
    19.98547, 19.98549, 19.98541, 19.98539, 19.98531, 19.98535, 19.98511, 
    19.98521, 19.98491, 19.985, 19.98556, 19.98553, 19.98544, 19.98549, 
    19.98536, 19.98533, 19.98531, 19.98527, 19.98527, 19.98525, 19.98528, 
    19.98525, 19.98537, 19.98532, 19.98545, 19.98542, 19.98544, 19.98545, 
    19.9854, 19.98534, 19.98534, 19.98532, 19.98528, 19.98536, 19.98509, 
    19.98526, 19.98551, 19.98546, 19.98545, 19.98547, 19.98533, 19.98538, 
    19.98525, 19.98529, 19.98523, 19.98526, 19.98526, 19.9853, 19.98532, 
    19.98538, 19.98543, 19.98547, 19.98546, 19.98541, 19.98534, 19.98527, 
    19.98529, 19.98523, 19.98537, 19.98531, 19.98534, 19.98528, 19.9854, 
    19.9853, 19.98543, 19.98542, 19.98538, 19.98531, 19.98529, 19.98528, 
    19.98529, 19.98534, 19.98535, 19.98538, 19.9854, 19.98542, 19.98545, 
    19.98543, 19.9854, 19.98534, 19.98528, 19.98522, 19.9852, 19.98513, 
    19.98519, 19.98509, 19.98517, 19.98503, 19.98529, 19.98518, 19.98538, 
    19.98536, 19.98532, 19.98523, 19.98528, 19.98522, 19.98535, 19.98541, 
    19.98543, 19.98546, 19.98543, 19.98543, 19.9854, 19.98541, 19.98534, 
    19.98538, 19.98526, 19.98522, 19.9851, 19.98503, 19.98496, 19.98492, 
    19.98491, 19.98491,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N =
  0.7222453, 0.7222428, 0.7222433, 0.7222412, 0.7222424, 0.722241, 0.7222448, 
    0.7222427, 0.722244, 0.7222451, 0.7222373, 0.7222412, 0.7222333, 
    0.7222357, 0.7222295, 0.7222337, 0.7222288, 0.7222297, 0.7222269, 
    0.7222276, 0.722224, 0.7222264, 0.7222221, 0.7222246, 0.7222242, 
    0.7222266, 0.7222404, 0.7222378, 0.7222405, 0.7222401, 0.7222403, 
    0.7222424, 0.7222434, 0.7222455, 0.7222451, 0.7222435, 0.72224, 
    0.7222412, 0.7222382, 0.7222382, 0.7222348, 0.7222364, 0.7222307, 
    0.7222323, 0.7222276, 0.7222288, 0.7222277, 0.722228, 0.7222277, 
    0.7222294, 0.7222286, 0.7222302, 0.7222361, 0.7222344, 0.7222396, 
    0.7222427, 0.7222447, 0.7222462, 0.722246, 0.7222456, 0.7222435, 
    0.7222416, 0.7222401, 0.7222392, 0.7222382, 0.7222353, 0.7222338, 
    0.7222304, 0.722231, 0.7222299, 0.7222289, 0.7222272, 0.7222275, 
    0.7222267, 0.72223, 0.7222278, 0.7222313, 0.7222304, 0.722238, 0.7222409, 
    0.7222421, 0.7222432, 0.7222458, 0.722244, 0.7222447, 0.722243, 
    0.7222419, 0.7222425, 0.7222392, 0.7222404, 0.7222337, 0.7222366, 
    0.722229, 0.7222309, 0.7222286, 0.7222297, 0.7222278, 0.7222295, 
    0.7222265, 0.7222258, 0.7222263, 0.7222245, 0.7222297, 0.7222277, 
    0.7222425, 0.7222424, 0.722242, 0.7222438, 0.7222439, 0.7222455, 
    0.7222441, 0.7222434, 0.7222419, 0.7222409, 0.72224, 0.7222381, 
    0.7222359, 0.7222329, 0.7222307, 0.7222292, 0.7222301, 0.7222294, 
    0.7222303, 0.7222307, 0.7222261, 0.7222286, 0.7222248, 0.722225, 
    0.7222267, 0.722225, 0.7222424, 0.7222428, 0.7222446, 0.7222432, 
    0.7222457, 0.7222443, 0.7222435, 0.7222404, 0.7222397, 0.7222391, 
    0.7222379, 0.7222363, 0.7222335, 0.7222311, 0.7222289, 0.722229, 
    0.7222289, 0.7222285, 0.7222297, 0.7222283, 0.7222281, 0.7222286, 
    0.722225, 0.7222261, 0.722225, 0.7222257, 0.7222427, 0.7222418, 
    0.7222423, 0.7222414, 0.7222421, 0.7222394, 0.7222385, 0.7222348, 
    0.7222363, 0.7222339, 0.7222361, 0.7222357, 0.7222338, 0.722236, 
    0.7222312, 0.7222344, 0.7222285, 0.7222317, 0.7222282, 0.7222289, 
    0.7222278, 0.7222269, 0.7222258, 0.7222236, 0.7222241, 0.7222223, 
    0.7222406, 0.7222395, 0.7222396, 0.7222384, 0.7222376, 0.7222357, 
    0.7222328, 0.7222339, 0.7222319, 0.7222314, 0.7222345, 0.7222326, 
    0.7222387, 0.7222378, 0.7222384, 0.7222405, 0.7222337, 0.7222372, 
    0.7222307, 0.7222326, 0.722227, 0.7222298, 0.7222244, 0.7222221, 
    0.7222199, 0.7222174, 0.7222389, 0.7222396, 0.7222383, 0.7222365, 
    0.7222347, 0.7222325, 0.7222322, 0.7222318, 0.7222307, 0.7222298, 
    0.7222317, 0.7222295, 0.7222375, 0.7222334, 0.7222399, 0.7222379, 
    0.7222366, 0.7222372, 0.722234, 0.7222333, 0.7222303, 0.7222319, 
    0.7222226, 0.7222267, 0.7222154, 0.7222186, 0.7222399, 0.7222389, 
    0.7222354, 0.7222371, 0.7222323, 0.7222311, 0.7222302, 0.722229, 
    0.7222289, 0.7222282, 0.7222293, 0.7222282, 0.7222325, 0.7222306, 
    0.7222358, 0.7222345, 0.7222351, 0.7222357, 0.7222338, 0.7222316, 
    0.7222316, 0.7222309, 0.722229, 0.7222323, 0.7222221, 0.7222284, 
    0.7222378, 0.7222359, 0.7222356, 0.7222363, 0.7222313, 0.7222331, 
    0.7222282, 0.7222295, 0.7222273, 0.7222284, 0.7222286, 0.72223, 
    0.7222309, 0.722233, 0.7222348, 0.7222362, 0.7222359, 0.7222344, 
    0.7222315, 0.7222289, 0.7222294, 0.7222275, 0.7222326, 0.7222305, 
    0.7222313, 0.7222291, 0.722234, 0.7222298, 0.722235, 0.7222345, 
    0.7222331, 0.7222303, 0.7222297, 0.7222291, 0.7222295, 0.7222314, 
    0.7222318, 0.7222332, 0.7222336, 0.7222346, 0.7222355, 0.7222347, 
    0.7222339, 0.7222314, 0.7222293, 0.7222269, 0.7222263, 0.7222236, 
    0.7222258, 0.7222221, 0.7222252, 0.7222198, 0.7222296, 0.7222254, 
    0.7222331, 0.7222322, 0.7222307, 0.7222273, 0.7222291, 0.722227, 
    0.7222318, 0.7222343, 0.722235, 0.7222362, 0.7222349, 0.722235, 
    0.7222338, 0.7222342, 0.7222314, 0.7222329, 0.7222286, 0.722227, 
    0.7222225, 0.7222198, 0.722217, 0.7222158, 0.7222154, 0.7222152 ;

 SOIL1N_TNDNCY_VERT_TRANS =
  -5.139921e-21, -1.541976e-20, 5.139921e-21, 3.597945e-20, -2.569961e-20, 
    -2.006177e-36, -5.139921e-21, -2.006177e-36, 1.027984e-20, 5.139921e-21, 
    -1.541976e-20, -3.083953e-20, -2.569961e-20, 5.139921e-21, 1.027984e-20, 
    2.006177e-36, 5.139921e-21, 2.006177e-36, -1.027984e-20, -2.569961e-20, 
    -2.569961e-20, 5.139921e-21, 3.083953e-20, -5.139921e-21, 1.541976e-20, 
    -5.139921e-21, 5.139921e-21, 6.681898e-20, 1.027984e-20, 2.055969e-20, 
    -1.541976e-20, 2.006177e-36, 1.541976e-20, -1.027984e-20, -2.055969e-20, 
    1.027984e-20, -1.027984e-20, -1.541976e-20, 3.597945e-20, 5.139921e-21, 
    5.139921e-21, -1.027984e-20, 5.139921e-21, 1.027984e-20, -1.541976e-20, 
    -2.055969e-20, 1.541976e-20, -1.027984e-20, 1.027984e-20, 1.027984e-20, 
    -2.055969e-20, 5.139921e-21, -5.139921e-21, -3.597945e-20, -5.139921e-21, 
    -2.055969e-20, 0, -2.006177e-36, 3.597945e-20, 2.569961e-20, 
    5.139921e-21, -1.541976e-20, 1.027984e-20, 5.139921e-21, 1.027984e-20, 
    5.139921e-21, -1.541976e-20, 1.541976e-20, -1.027984e-20, 5.139921e-20, 
    2.569961e-20, 2.569961e-20, -1.027984e-20, 1.027984e-20, -5.139921e-21, 
    -1.541976e-20, 3.083953e-20, -4.111937e-20, 1.541976e-20, 5.139921e-21, 
    5.139921e-21, 2.006177e-36, 5.139921e-21, -5.139921e-21, 1.541976e-20, 
    -1.027984e-20, -1.027984e-20, 3.083953e-20, -5.139921e-21, -1.541976e-20, 
    2.569961e-20, 1.027984e-20, -2.006177e-36, 1.541976e-20, -1.027984e-20, 
    -1.541976e-20, -1.541976e-20, -1.541976e-20, 1.541976e-20, 4.111937e-20, 
    5.139921e-21, 0, -2.055969e-20, 1.541976e-20, 2.055969e-20, 
    -5.139921e-20, 2.006177e-36, 1.027984e-20, 2.055969e-20, 2.569961e-20, 
    2.055969e-20, -5.139921e-20, 2.006177e-36, 2.569961e-20, 0, 
    -1.541976e-20, -5.139921e-21, 1.541976e-20, 1.541976e-20, 0, 
    2.055969e-20, 2.569961e-20, 1.541976e-20, -2.055969e-20, 5.139921e-21, 
    1.541976e-20, 1.541976e-20, 5.139921e-21, 5.139921e-21, 1.541976e-20, 
    -2.055969e-20, -5.139921e-21, 1.027984e-20, -3.083953e-20, 1.541976e-20, 
    3.597945e-20, -1.541976e-20, 2.055969e-20, 1.541976e-20, 2.055969e-20, 
    -3.083953e-20, -1.027984e-20, -4.625929e-20, 5.139921e-21, 1.027984e-20, 
    -1.541976e-20, 0, -5.139921e-21, 0, 0, -2.569961e-20, -2.569961e-20, 
    1.027984e-20, 2.006177e-36, 5.139921e-21, 5.139921e-21, -5.139921e-21, 
    2.569961e-20, 1.027984e-20, 3.083953e-20, 1.541976e-20, -3.597945e-20, 0, 
    -2.055969e-20, -1.541976e-20, -1.027984e-20, 0, 0, -5.139921e-21, 
    2.569961e-20, 1.027984e-20, -5.139921e-21, -2.055969e-20, 5.139921e-21, 
    0, 1.027984e-20, 1.027984e-20, -1.541976e-20, -1.541976e-20, 
    2.055969e-20, 3.597945e-20, 1.541976e-20, -2.569961e-20, 3.597945e-20, 
    -2.055969e-20, 1.027984e-20, 0, 3.597945e-20, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, -5.139921e-21, 1.541976e-20, 1.541976e-20, 
    2.569961e-20, -1.027984e-20, -1.027984e-20, 1.027984e-20, 5.139921e-21, 
    -1.541976e-20, -1.027984e-20, -2.055969e-20, 2.569961e-20, -1.541976e-20, 
    1.027984e-20, 2.006177e-36, 2.569961e-20, 1.027984e-20, 2.055969e-20, 
    -2.006177e-36, -1.027984e-20, -6.167906e-20, 0, -1.027984e-20, 
    4.625929e-20, 3.083953e-20, 4.625929e-20, 5.139921e-21, -1.027984e-20, 0, 
    1.027984e-20, -5.139921e-21, 1.541976e-20, 1.541976e-20, -5.139921e-21, 
    -1.027984e-20, 1.027984e-20, -2.055969e-20, 2.006177e-36, 5.139921e-21, 
    5.139921e-21, 1.541976e-20, -1.027984e-20, -1.027984e-20, 1.027984e-20, 
    5.139921e-21, -1.541976e-20, 1.027984e-20, -2.055969e-20, -1.541976e-20, 
    -2.569961e-20, -5.139921e-21, -1.541976e-20, -1.541976e-20, 
    -1.541976e-20, 1.541976e-20, 1.541976e-20, -5.139921e-21, 0, 
    -5.139921e-21, 0, 5.139921e-21, -1.541976e-20, 2.006177e-36, 
    -1.541976e-20, 5.139921e-21, 2.006177e-36, 5.139921e-21, -3.597945e-20, 
    -5.139921e-21, 3.083953e-20, -5.139921e-21, -1.541976e-20, -5.139921e-21, 
    2.569961e-20, 1.541976e-20, 2.569961e-20, 2.055969e-20, 1.027984e-20, 
    -2.055969e-20, 1.027984e-20, 2.569961e-20, -5.139921e-21, 1.541976e-20, 
    1.541976e-20, -2.569961e-20, 2.569961e-20, -5.139921e-21, 5.139921e-21, 
    1.541976e-20, 5.139921e-21, 3.083953e-20, -1.541976e-20, -5.139921e-21, 
    1.027984e-20, 5.139921e-21, -1.541976e-20, -1.027984e-20, 0, 
    1.027984e-20, 3.083953e-20, 2.569961e-20, -5.139921e-21, -2.055969e-20, 
    1.541976e-20, -1.541976e-20, 1.027984e-20, 1.027984e-20, -1.541976e-20, 
    -3.083953e-20, -2.055969e-20, 1.541976e-20, -2.006177e-36, 0, 
    1.027984e-20, -5.139921e-21, 2.569961e-20, 1.027984e-20, -2.055969e-20, 
    0, 0, 1.541976e-20, 2.569961e-20, 0, 1.541976e-20, 2.055969e-20, 
    -3.083953e-20, 5.139921e-21, 5.139921e-21, 0, -1.541976e-20, 
    -2.569961e-20, 1.541976e-20, 0, -5.139921e-21, 1.027984e-20, 
    1.027984e-20, -2.569961e-20, -1.027984e-20, -5.139921e-21, 1.541976e-20, 
    5.139921e-21, -1.541976e-20, 2.006177e-36, -2.055969e-20, 2.055969e-20, 
    5.139921e-21, 5.139921e-21,
  -1.541976e-20, 5.139921e-21, -1.027984e-20, 1.027984e-20, 2.055969e-20, 
    -5.139921e-21, 5.139921e-21, 1.027984e-20, -1.027984e-20, 0, 
    -1.027984e-20, 5.139921e-21, 5.139921e-21, 3.083953e-20, 2.055969e-20, 
    2.006177e-36, -5.139921e-21, -5.139921e-21, 2.055969e-20, 2.006177e-36, 
    0, -4.625929e-20, -2.006177e-36, 2.055969e-20, 5.139921e-21, 
    2.055969e-20, -2.569961e-20, 1.027984e-20, -5.139921e-21, -2.006177e-36, 
    1.541976e-20, -2.569961e-20, 1.027984e-20, -1.027984e-20, 1.027984e-20, 
    0, -1.027984e-20, -5.139921e-21, -1.027984e-20, -3.083953e-20, 
    -3.083953e-20, 1.541976e-20, -5.139921e-21, 1.027984e-20, -1.541976e-20, 
    3.083953e-20, 0, -1.027984e-20, -5.139921e-21, 0, -2.055969e-20, 
    -1.541976e-20, -5.139921e-21, 5.139921e-21, -2.055969e-20, 1.027984e-20, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, 2.055969e-20, -1.541976e-20, 
    2.055969e-20, -1.027984e-20, 1.541976e-20, 1.027984e-20, 5.139921e-21, 
    -2.006177e-36, 0, 1.027984e-20, 1.027984e-20, 5.139921e-21, 5.139921e-21, 
    0, 1.027984e-20, -1.027984e-20, 5.139921e-21, 0, 1.541976e-20, 
    1.541976e-20, 0, 5.139921e-21, 2.006177e-36, -2.569961e-20, 
    -1.541976e-20, -1.541976e-20, 2.006177e-36, -5.139921e-21, -5.139921e-21, 
    1.027984e-20, 0, 5.139921e-21, -2.055969e-20, 1.027984e-20, 
    -1.027984e-20, 3.083953e-20, -2.006177e-36, -5.139921e-21, -5.139921e-21, 
    -2.055969e-20, -1.541976e-20, -2.006177e-36, 1.027984e-20, 1.541976e-20, 
    1.541976e-20, 5.139921e-21, 5.139921e-21, 1.027984e-20, 5.139921e-21, 
    1.541976e-20, 1.027984e-20, 1.541976e-20, -3.083953e-20, -5.139921e-21, 
    5.139921e-21, 1.541976e-20, -2.055969e-20, 2.055969e-20, 0, 
    -1.541976e-20, 0, 1.541976e-20, 1.027984e-20, 3.083953e-20, 
    -1.027984e-20, -2.055969e-20, -1.027984e-20, -5.139921e-21, 2.006177e-36, 
    1.027984e-20, 1.027984e-20, 0, 1.027984e-20, 0, 1.027984e-20, 
    -5.139921e-21, 5.139921e-21, 1.541976e-20, -1.541976e-20, -4.625929e-20, 
    -2.055969e-20, 2.569961e-20, -1.027984e-20, -1.541976e-20, -1.027984e-20, 
    -1.027984e-20, 1.027984e-20, -1.027984e-20, -2.006177e-36, 5.139921e-21, 
    1.027984e-20, 1.541976e-20, 5.139921e-21, -5.139921e-21, 0, 
    -1.541976e-20, -1.027984e-20, -1.541976e-20, 1.541976e-20, -1.027984e-20, 
    1.027984e-20, 2.055969e-20, 1.541976e-20, 0, -2.055969e-20, 0, 
    1.027984e-20, 1.541976e-20, 0, 2.055969e-20, -1.027984e-20, 1.541976e-20, 
    5.139921e-21, -1.027984e-20, -5.139921e-21, 2.569961e-20, 5.139921e-21, 
    -1.027984e-20, 0, 0, 0, 1.027984e-20, -1.027984e-20, 5.139921e-21, 
    5.139921e-21, -2.006177e-36, -1.541976e-20, 0, -5.139921e-21, 
    -5.139921e-21, 2.569961e-20, 5.139921e-21, 5.139921e-21, -1.027984e-20, 
    -5.139921e-21, 5.139921e-21, -1.541976e-20, 3.083953e-20, -2.055969e-20, 
    1.027984e-20, -1.027984e-20, 5.139921e-21, 2.569961e-20, 5.139921e-21, 
    -1.027984e-20, 1.541976e-20, -2.055969e-20, 1.541976e-20, -2.569961e-20, 
    5.139921e-21, 5.139921e-21, 0, 1.027984e-20, 2.006177e-36, 1.541976e-20, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20, -2.006177e-36, 2.006177e-36, 
    -1.541976e-20, -5.139921e-21, -1.541976e-20, 1.541976e-20, -1.541976e-20, 
    1.027984e-20, 1.541976e-20, 5.139921e-21, 2.569961e-20, -1.027984e-20, 0, 
    0, 1.027984e-20, 2.569961e-20, -2.055969e-20, 0, -5.139921e-21, 
    1.541976e-20, 1.027984e-20, -5.139921e-21, -1.027984e-20, 0, 
    -1.027984e-20, -5.139921e-21, -2.055969e-20, -2.569961e-20, 
    -2.055969e-20, 3.083953e-20, 2.569961e-20, 1.027984e-20, 1.541976e-20, 
    1.027984e-20, 1.027984e-20, 2.055969e-20, -5.139921e-21, -1.541976e-20, 
    -1.027984e-20, 0, 1.027984e-20, -3.083953e-20, -1.027984e-20, 
    -5.139921e-20, -5.139921e-21, 1.027984e-20, -3.597945e-20, -1.027984e-20, 
    -1.541976e-20, -2.055969e-20, -1.541976e-20, 5.139921e-21, -1.027984e-20, 
    1.541976e-20, 1.027984e-20, 5.139921e-21, 0, 0, -1.541976e-20, 
    1.027984e-20, 2.055969e-20, -1.027984e-20, 1.027984e-20, -5.139921e-21, 
    2.569961e-20, -5.139921e-21, -1.027984e-20, 1.541976e-20, 1.027984e-20, 
    0, 0, -1.027984e-20, -1.027984e-20, -2.055969e-20, 5.139921e-21, 
    -1.541976e-20, 3.083953e-20, -1.541976e-20, 2.569961e-20, 1.027984e-20, 
    2.055969e-20, -3.597945e-20, -2.055969e-20, -1.541976e-20, -2.055969e-20, 
    -5.139921e-21, -5.139921e-21, -5.139921e-21, 2.055969e-20, -2.055969e-20, 
    2.569961e-20, 5.139921e-21, -1.027984e-20, -1.541976e-20, -1.541976e-20, 
    1.541976e-20, -1.027984e-20, -2.569961e-20, 5.139921e-21, -2.569961e-20, 
    -1.027984e-20, 1.541976e-20, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    -1.027984e-20, 1.027984e-20, 5.139921e-21, 4.111937e-20, -5.139921e-21, 
    -1.541976e-20, 2.006177e-36, 1.027984e-20, 5.139921e-21, 0, 
    -1.027984e-20, -1.541976e-20, -5.139921e-21, -2.006177e-36, 0, 
    5.139921e-21,
  1.541976e-20, -1.541976e-20, 1.541976e-20, 5.139921e-21, 1.541976e-20, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20, -4.111937e-20, 1.027984e-20, 
    -2.055969e-20, 1.027984e-20, 1.027984e-20, -5.139921e-21, -1.541976e-20, 
    3.083953e-20, -3.597945e-20, 3.597945e-20, -1.541976e-20, 2.569961e-20, 
    1.541976e-20, 2.055969e-20, -1.541976e-20, 0, 1.027984e-20, 
    -1.027984e-20, 3.597945e-20, 0, -1.027984e-20, -1.541976e-20, 
    -1.027984e-20, -1.027984e-20, -2.055969e-20, 2.006177e-36, 5.139921e-21, 
    1.027984e-20, 0, -2.055969e-20, 0, 5.139921e-21, 5.139921e-21, 
    -2.569961e-20, 2.006177e-36, 5.139921e-21, 1.027984e-20, -5.139921e-21, 
    1.027984e-20, 5.139921e-21, -2.569961e-20, -1.541976e-20, 1.541976e-20, 
    -5.139921e-21, -1.027984e-20, -1.541976e-20, 1.027984e-20, 2.006177e-36, 
    -5.139921e-21, 2.006177e-36, 0, -5.139921e-21, 1.027984e-20, 
    -2.055969e-20, 3.083953e-20, 1.027984e-20, 2.055969e-20, -2.569961e-20, 
    -4.111937e-20, -5.139921e-21, 1.027984e-20, -2.006177e-36, 3.083953e-20, 
    -1.541976e-20, -1.541976e-20, 1.541976e-20, -1.027984e-20, 1.541976e-20, 
    2.055969e-20, -2.569961e-20, 2.055969e-20, -1.541976e-20, 2.569961e-20, 
    1.027984e-20, 1.541976e-20, 5.139921e-21, -5.139921e-21, 0, 1.541976e-20, 
    1.027984e-20, 2.006177e-36, -1.541976e-20, -5.139921e-21, 1.027984e-20, 
    5.139921e-21, 2.569961e-20, -5.139921e-21, -1.027984e-20, -1.541976e-20, 
    -1.027984e-20, 1.541976e-20, 2.569961e-20, 1.027984e-20, 3.597945e-20, 
    -5.139921e-21, -2.055969e-20, -1.027984e-20, -5.139921e-21, 5.139921e-21, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, -5.139921e-21, 1.027984e-20, 
    1.541976e-20, 0, 5.139921e-21, -2.055969e-20, 1.027984e-20, 3.083953e-20, 
    -5.139921e-21, 1.541976e-20, 1.541976e-20, -1.027984e-20, 1.027984e-20, 
    1.027984e-20, -1.541976e-20, 1.027984e-20, -1.541976e-20, 2.055969e-20, 
    -1.541976e-20, 3.083953e-20, -1.027984e-20, 1.027984e-20, 5.139921e-21, 
    -2.055969e-20, 1.027984e-20, 2.569961e-20, 0, 5.139921e-21, 5.139921e-21, 
    -5.139921e-21, -1.027984e-20, -5.139921e-21, 1.027984e-20, -5.139921e-20, 
    1.027984e-20, 1.027984e-20, -2.055969e-20, -1.027984e-20, -2.055969e-20, 
    5.139921e-21, -2.569961e-20, 2.569961e-20, 1.027984e-20, -1.027984e-20, 
    -5.139921e-21, -1.541976e-20, -2.006177e-36, 1.027984e-20, -3.083953e-20, 
    -5.139921e-21, 1.027984e-20, 0, 2.055969e-20, 0, 0, 0, -1.027984e-20, 
    5.139921e-21, 3.083953e-20, -2.569961e-20, -2.569961e-20, 2.055969e-20, 
    2.006177e-36, 2.006177e-36, 2.569961e-20, -4.111937e-20, -2.006177e-36, 
    1.027984e-20, -1.027984e-20, -2.055969e-20, 1.027984e-20, -5.139921e-21, 
    1.027984e-20, -1.027984e-20, 5.139921e-21, 5.139921e-21, -3.597945e-20, 
    1.541976e-20, -1.541976e-20, 1.027984e-20, 0, -1.027984e-20, 
    -5.139921e-21, 3.597945e-20, 1.027984e-20, 1.027984e-20, -1.027984e-20, 
    2.055969e-20, 3.597945e-20, 5.139921e-21, -1.027984e-20, 1.541976e-20, 0, 
    0, 3.083953e-20, 2.569961e-20, -2.055969e-20, -1.027984e-20, 0, 0, 
    2.569961e-20, -2.569961e-20, -1.541976e-20, 0, 3.083953e-20, 
    -2.006177e-36, -3.597945e-20, 5.139921e-21, 5.139921e-21, 4.111937e-20, 
    2.569961e-20, 0, -2.055969e-20, 2.569961e-20, 5.139921e-21, 
    -1.541976e-20, 1.027984e-20, 0, 1.541976e-20, -5.139921e-21, 
    -5.139921e-21, -1.541976e-20, -1.027984e-20, 1.541976e-20, -1.027984e-20, 
    1.027984e-20, -2.569961e-20, 1.027984e-20, -2.055969e-20, -5.653913e-20, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20, -2.055969e-20, 1.027984e-20, 
    5.139921e-21, 1.027984e-20, -1.027984e-20, -5.139921e-21, 1.027984e-20, 
    0, -5.139921e-21, 0, 1.027984e-20, 1.027984e-20, 3.597945e-20, 
    -2.055969e-20, 3.083953e-20, 1.027984e-20, -1.027984e-20, 1.027984e-20, 
    -1.027984e-20, 5.139921e-21, 3.597945e-20, -1.541976e-20, -5.139921e-21, 
    5.139921e-21, -2.569961e-20, -5.139921e-21, 0, 2.055969e-20, 
    2.006177e-36, -2.055969e-20, 0, -3.083953e-20, 5.139921e-21, 
    1.541976e-20, 2.569961e-20, 1.027984e-20, -1.541976e-20, 3.083953e-20, 
    -1.027984e-20, -3.083953e-20, -2.006177e-36, 2.006177e-36, 2.055969e-20, 
    -1.541976e-20, 2.569961e-20, 1.541976e-20, -1.541976e-20, 1.027984e-20, 
    -5.139921e-21, -1.541976e-20, 5.139921e-21, -3.083953e-20, -1.027984e-20, 
    -1.027984e-20, 1.027984e-20, 5.139921e-21, 0, -2.006177e-36, 
    -5.139921e-21, 0, -2.569961e-20, -1.027984e-20, -1.541976e-20, 
    -1.027984e-20, -1.027984e-20, -1.027984e-20, 5.139921e-21, 1.027984e-20, 
    1.541976e-20, 1.027984e-20, 1.027984e-20, -2.569961e-20, -5.139921e-21, 
    -1.541976e-20, 2.055969e-20, 1.027984e-20, 1.027984e-20, -2.055969e-20, 
    -1.027984e-20, -1.541976e-20, 1.027984e-20, 5.139921e-21, -2.055969e-20, 
    -1.541976e-20, 0, -1.027984e-20, 5.139921e-21, -1.541976e-20, 
    -1.027984e-20, 0, -2.055969e-20, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, -5.139921e-21,
  -1.027984e-20, 1.027984e-20, 5.139921e-21, -1.541976e-20, -1.541976e-20, 
    5.139921e-21, 1.541976e-20, -1.541976e-20, 3.597945e-20, -5.139921e-21, 
    -2.569961e-20, 0, -5.139921e-21, -1.027984e-20, 1.541976e-20, 
    -1.541976e-20, -3.083953e-20, 5.139921e-21, 5.139921e-21, -2.055969e-20, 
    -1.541976e-20, -2.569961e-20, -3.083953e-20, -2.055969e-20, 4.111937e-20, 
    -5.139921e-21, 0, 3.597945e-20, -5.139921e-21, -2.006177e-36, 
    2.055969e-20, 1.541976e-20, 5.139921e-21, -1.541976e-20, -2.569961e-20, 
    -1.541976e-20, -5.139921e-21, -1.541976e-20, 2.055969e-20, 1.541976e-20, 
    1.541976e-20, 1.027984e-20, -5.139921e-21, -3.083953e-20, -5.139921e-21, 
    5.139921e-21, -2.569961e-20, -1.541976e-20, -5.139921e-21, 1.027984e-20, 
    2.006177e-36, -5.139921e-21, -1.027984e-20, -4.111937e-20, -2.055969e-20, 
    1.027984e-20, -1.027984e-20, 2.055969e-20, 0, 5.139921e-21, 
    -1.541976e-20, 3.083953e-20, -1.027984e-20, 3.083953e-20, 5.139921e-21, 
    -1.541976e-20, 4.111937e-20, -5.139921e-21, 0, 3.083953e-20, 
    -1.027984e-20, -1.541976e-20, -5.139921e-21, 2.569961e-20, -1.541976e-20, 
    2.055969e-20, -1.027984e-20, -3.083953e-20, 5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 1.541976e-20, 4.111937e-20, 5.139921e-21, -1.027984e-20, 
    2.569961e-20, -1.027984e-20, -6.167906e-20, 2.006177e-36, -1.027984e-20, 
    1.541976e-20, 1.541976e-20, -5.139921e-21, -1.541976e-20, -1.027984e-20, 
    2.569961e-20, 1.027984e-20, -1.027984e-20, 3.597945e-20, 1.027984e-20, 
    1.541976e-20, -4.111937e-20, -1.541976e-20, 1.027984e-20, 5.139921e-21, 
    1.541976e-20, -4.111937e-20, 3.083953e-20, -4.111937e-20, 1.541976e-20, 
    1.027984e-20, 1.027984e-20, 3.083953e-20, -2.569961e-20, 2.055969e-20, 
    1.027984e-20, 1.027984e-20, 1.027984e-20, -1.541976e-20, 2.055969e-20, 
    1.027984e-20, 2.569961e-20, 1.027984e-20, -5.139921e-21, -2.055969e-20, 
    3.083953e-20, -5.139921e-21, -4.111937e-20, -3.083953e-20, -1.027984e-20, 
    1.541976e-20, 2.055969e-20, 2.569961e-20, 1.541976e-20, 2.569961e-20, 
    -1.027984e-20, -1.541976e-20, 0, 2.569961e-20, -5.139921e-21, 
    5.139921e-21, 1.541976e-20, 0, 1.027984e-20, 5.139921e-21, 2.055969e-20, 
    0, 0, 1.027984e-20, -1.027984e-20, 3.083953e-20, 2.055969e-20, 
    3.083953e-20, -2.569961e-20, 1.541976e-20, 2.569961e-20, -1.027984e-20, 
    -1.027984e-20, -5.139921e-21, 1.027984e-20, 5.139921e-21, 5.139921e-21, 
    5.139921e-21, 1.027984e-20, -1.541976e-20, -1.027984e-20, -1.027984e-20, 
    -3.083953e-20, -5.139921e-21, 1.541976e-20, -1.541976e-20, -1.027984e-20, 
    1.541976e-20, 2.055969e-20, 1.541976e-20, 2.006177e-36, -2.569961e-20, 
    -1.027984e-20, 4.625929e-20, 2.569961e-20, 1.027984e-20, 1.027984e-20, 
    -2.055969e-20, 0, -4.625929e-20, -2.055969e-20, 2.055969e-20, 
    2.569961e-20, 2.055969e-20, 2.055969e-20, -2.055969e-20, -1.027984e-20, 
    -5.139921e-20, -5.139921e-21, 1.027984e-20, -5.139921e-21, 2.569961e-20, 
    1.541976e-20, 1.541976e-20, 2.569961e-20, -1.541976e-20, -5.139921e-21, 
    4.111937e-20, 5.139921e-21, 3.083953e-20, -2.055969e-20, -1.027984e-20, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, 1.027984e-20, -1.541976e-20, 
    2.006177e-36, 2.055969e-20, -2.055969e-20, 1.541976e-20, -2.055969e-20, 
    -1.027984e-20, 3.083953e-20, -1.541976e-20, 1.027984e-20, -2.055969e-20, 
    -1.027984e-20, -2.055969e-20, -5.139921e-21, -5.139921e-21, 
    -3.083953e-20, 5.139921e-21, -1.027984e-20, 2.055969e-20, 2.569961e-20, 
    2.006177e-36, -2.055969e-20, 1.027984e-20, 0, -5.139921e-21, 
    2.006177e-36, -1.027984e-20, 1.027984e-20, -2.569961e-20, 2.055969e-20, 
    -2.569961e-20, -2.055969e-20, 1.027984e-20, 3.083953e-20, -1.027984e-20, 
    -5.139921e-21, 2.055969e-20, 5.139921e-21, 1.027984e-20, -2.569961e-20, 
    1.541976e-20, 1.027984e-20, 5.139921e-21, -2.055969e-20, 4.625929e-20, 
    1.541976e-20, 2.055969e-20, -5.139921e-21, -1.027984e-20, -5.653913e-20, 
    -1.541976e-20, -5.139921e-21, -5.139921e-21, 0, 1.027984e-20, 0, 
    1.027984e-20, -2.055969e-20, -5.139921e-21, 0, 3.597945e-20, 
    1.027984e-20, 1.027984e-20, -5.139921e-21, -1.541976e-20, -5.139921e-21, 
    -1.027984e-20, -2.569961e-20, 1.027984e-20, 1.027984e-20, 5.139921e-21, 
    -2.569961e-20, 2.569961e-20, 5.139921e-21, 2.055969e-20, 5.139921e-21, 
    -1.541976e-20, -5.139921e-21, 3.083953e-20, -3.083953e-20, 5.653913e-20, 
    5.139921e-21, 1.541976e-20, -3.597945e-20, -2.569961e-20, 0, 
    5.139921e-21, 5.139921e-21, -3.597945e-20, 2.055969e-20, -2.055969e-20, 
    5.139921e-21, 2.055969e-20, 5.139921e-21, -1.027984e-20, -2.055969e-20, 
    1.541976e-20, 4.111937e-20, 5.139921e-21, -2.569961e-20, 2.055969e-20, 
    2.569961e-20, -2.569961e-20, 3.083953e-20, 2.569961e-20, 0, 
    -1.541976e-20, -5.139921e-21, -1.027984e-20, 2.569961e-20, -1.541976e-20, 
    -5.139921e-21, 1.541976e-20, 1.541976e-20, -1.027984e-20, 5.139921e-21, 
    1.027984e-20, 2.569961e-20, -1.027984e-20, -5.139921e-21, -5.139921e-20, 
    5.139921e-21, -1.541976e-20, -5.139921e-21, 1.027984e-20, -2.055969e-20, 
    3.083953e-20,
  1.027984e-20, -1.027984e-20, 3.083953e-20, 5.139921e-21, 1.027984e-20, 
    5.139921e-21, -2.055969e-20, -1.027984e-20, 2.569961e-20, 2.569961e-20, 
    0, 2.569961e-20, 5.139921e-21, 2.006177e-36, 1.027984e-20, -1.027984e-20, 
    1.027984e-20, 1.027984e-20, -2.055969e-20, -1.027984e-20, -1.541976e-20, 
    3.597945e-20, -3.083953e-20, -1.541976e-20, 2.055969e-20, 5.139921e-21, 
    -5.139921e-21, -1.027984e-20, -2.055969e-20, -1.541976e-20, 1.027984e-20, 
    -2.569961e-20, -2.569961e-20, 1.541976e-20, -5.139921e-21, 1.027984e-20, 
    -1.027984e-20, -1.027984e-20, -1.027984e-20, 2.569961e-20, 1.027984e-20, 
    -2.055969e-20, 5.139921e-21, 2.569961e-20, 1.027984e-20, 1.541976e-20, 
    1.027984e-20, -2.055969e-20, -1.541976e-20, 5.139921e-21, 1.541976e-20, 
    1.027984e-20, -2.569961e-20, -5.139921e-21, 2.055969e-20, 2.569961e-20, 
    -2.569961e-20, 0, 2.569961e-20, 1.027984e-20, 0, -5.139921e-21, 
    2.006177e-36, -3.083953e-20, -2.055969e-20, -3.083953e-20, -1.541976e-20, 
    1.541976e-20, -2.006177e-36, -5.139921e-21, 1.027984e-20, 3.083953e-20, 
    0, -2.006177e-36, 1.027984e-20, -2.569961e-20, 1.027984e-20, 
    -1.541976e-20, -2.569961e-20, -1.541976e-20, 1.027984e-20, -5.139921e-21, 
    2.006177e-36, 3.083953e-20, 2.055969e-20, 5.139921e-21, -3.597945e-20, 
    -5.139921e-21, -1.027984e-20, -1.027984e-20, 5.139921e-21, -5.139921e-21, 
    1.027984e-20, -4.111937e-20, -1.541976e-20, -1.027984e-20, -1.027984e-20, 
    -5.139921e-21, 2.569961e-20, 5.139921e-21, -4.111937e-20, 0, 0, 
    -1.541976e-20, 0, -2.055969e-20, 5.139921e-21, -5.139921e-21, 
    -2.055969e-20, 0, -4.111937e-20, 5.139921e-21, -1.541976e-20, 
    5.139921e-21, -5.139921e-21, 2.569961e-20, -3.083953e-20, 2.055969e-20, 
    1.027984e-20, 2.569961e-20, 5.139921e-21, -2.006177e-36, -2.055969e-20, 
    5.139921e-21, -5.139921e-21, -1.541976e-20, -1.541976e-20, 5.139921e-21, 
    -2.055969e-20, 5.139921e-21, 5.139921e-21, 2.055969e-20, -1.027984e-20, 
    -2.569961e-20, -2.055969e-20, -1.027984e-20, 3.083953e-20, -1.541976e-20, 
    0, -3.083953e-20, 1.027984e-20, 1.541976e-20, 5.139921e-21, 
    -1.541976e-20, 1.541976e-20, 3.083953e-20, -2.055969e-20, 0, 
    2.055969e-20, 1.027984e-20, 1.027984e-20, -5.139921e-21, 5.139921e-21, 
    5.139921e-21, 1.027984e-20, -1.541976e-20, -2.055969e-20, 1.541976e-20, 
    -5.139921e-21, 2.055969e-20, -2.569961e-20, 0, -3.597945e-20, 
    1.541976e-20, 5.139921e-21, 3.597945e-20, -1.541976e-20, -5.139921e-21, 
    -1.027984e-20, 3.083953e-20, -5.139921e-21, -1.541976e-20, -3.597945e-20, 
    -2.569961e-20, 1.541976e-20, 5.139921e-21, 0, -5.139921e-21, 
    5.139921e-21, 1.541976e-20, 0, -2.569961e-20, -5.139921e-21, 
    -2.055969e-20, 1.541976e-20, 5.139921e-21, -5.139921e-21, 5.139921e-21, 
    1.541976e-20, 1.027984e-20, -1.541976e-20, 0, -1.027984e-20, 
    -2.055969e-20, 2.569961e-20, -1.541976e-20, -5.139921e-21, -1.541976e-20, 
    -2.055969e-20, -2.055969e-20, -2.055969e-20, 5.139921e-21, 0, 0, 
    -2.055969e-20, -1.027984e-20, 2.006177e-36, 1.027984e-20, 2.006177e-36, 
    -2.055969e-20, 2.055969e-20, 1.541976e-20, 3.083953e-20, -1.027984e-20, 
    2.006177e-36, 2.569961e-20, 1.027984e-20, 1.027984e-20, 5.139921e-21, 
    -5.139921e-21, 1.027984e-20, 1.541976e-20, -1.541976e-20, -1.541976e-20, 
    -2.055969e-20, -5.139921e-21, -1.027984e-20, -1.027984e-20, 0, 
    -1.541976e-20, 2.055969e-20, 0, 1.027984e-20, 2.055969e-20, 
    -1.027984e-20, 3.597945e-20, 1.027984e-20, 0, -1.027984e-20, 
    -1.027984e-20, -1.541976e-20, -1.541976e-20, 1.541976e-20, 1.027984e-20, 
    1.027984e-20, -1.027984e-20, -1.541976e-20, -5.139921e-21, 2.569961e-20, 
    -2.006177e-36, -5.139921e-21, 5.139921e-21, -1.541976e-20, -1.027984e-20, 
    2.569961e-20, 5.139921e-21, -3.083953e-20, 5.139921e-21, 1.541976e-20, 
    1.541976e-20, 1.541976e-20, -5.139921e-21, 1.027984e-20, -3.083953e-20, 
    5.139921e-21, -1.541976e-20, -1.027984e-20, 2.055969e-20, 2.055969e-20, 
    4.111937e-20, -1.541976e-20, 2.006177e-36, 1.027984e-20, -1.027984e-20, 
    5.139921e-21, -2.055969e-20, -1.027984e-20, -3.083953e-20, 1.027984e-20, 
    0, 1.541976e-20, 5.139921e-21, -5.139921e-21, -1.541976e-20, 
    2.006177e-36, 0, 3.083953e-20, -5.139921e-21, 5.139921e-21, 1.027984e-20, 
    -2.006177e-36, 1.541976e-20, 1.027984e-20, 2.569961e-20, -5.139921e-21, 
    7.709882e-20, -1.541976e-20, -1.541976e-20, 0, 1.541976e-20, 
    1.541976e-20, -3.083953e-20, -3.083953e-20, -1.541976e-20, -1.541976e-20, 
    3.083953e-20, -2.055969e-20, -1.541976e-20, -1.541976e-20, -1.541976e-20, 
    5.139921e-21, -3.083953e-20, -1.027984e-20, 0, 5.139921e-21, 0, 
    2.006177e-36, -3.083953e-20, 1.027984e-20, 5.139921e-21, 0, 3.597945e-20, 
    2.055969e-20, -1.541976e-20, -1.027984e-20, 5.139921e-21, 0, 
    5.139921e-21, 1.027984e-20, 0, -5.139921e-21, -1.027984e-20, 
    -3.597945e-20, -2.006177e-36, 1.541976e-20, 5.139921e-21, -2.006177e-36, 
    -5.139921e-21,
  8.598663e-29, 8.598634e-29, 8.59864e-29, 8.598617e-29, 8.59863e-29, 
    8.598615e-29, 8.598657e-29, 8.598634e-29, 8.598649e-29, 8.598661e-29, 
    8.598572e-29, 8.598616e-29, 8.598527e-29, 8.598555e-29, 8.598485e-29, 
    8.598531e-29, 8.598475e-29, 8.598486e-29, 8.598453e-29, 8.598463e-29, 
    8.598421e-29, 8.598449e-29, 8.5984e-29, 8.598428e-29, 8.598424e-29, 
    8.59845e-29, 8.598607e-29, 8.598578e-29, 8.598609e-29, 8.598605e-29, 
    8.598607e-29, 8.59863e-29, 8.598641e-29, 8.598666e-29, 8.598661e-29, 
    8.598643e-29, 8.598603e-29, 8.598616e-29, 8.598582e-29, 8.598583e-29, 
    8.598545e-29, 8.598562e-29, 8.598497e-29, 8.598516e-29, 8.598462e-29, 
    8.598476e-29, 8.598463e-29, 8.598467e-29, 8.598463e-29, 8.598483e-29, 
    8.598474e-29, 8.598491e-29, 8.598559e-29, 8.598539e-29, 8.598598e-29, 
    8.598633e-29, 8.598657e-29, 8.598673e-29, 8.598671e-29, 8.598666e-29, 
    8.598643e-29, 8.598622e-29, 8.598605e-29, 8.598594e-29, 8.598583e-29, 
    8.59855e-29, 8.598533e-29, 8.598494e-29, 8.598501e-29, 8.598489e-29, 
    8.598477e-29, 8.598458e-29, 8.598461e-29, 8.598453e-29, 8.598489e-29, 
    8.598465e-29, 8.598504e-29, 8.598494e-29, 8.59858e-29, 8.598613e-29, 
    8.598627e-29, 8.598639e-29, 8.598669e-29, 8.598648e-29, 8.598657e-29, 
    8.598637e-29, 8.598625e-29, 8.598631e-29, 8.598593e-29, 8.598608e-29, 
    8.598532e-29, 8.598565e-29, 8.598479e-29, 8.598499e-29, 8.598474e-29, 
    8.598486e-29, 8.598464e-29, 8.598485e-29, 8.59845e-29, 8.598442e-29, 
    8.598447e-29, 8.598427e-29, 8.598485e-29, 8.598463e-29, 8.598631e-29, 
    8.59863e-29, 8.598625e-29, 8.598646e-29, 8.598647e-29, 8.598666e-29, 
    8.598649e-29, 8.598642e-29, 8.598624e-29, 8.598614e-29, 8.598604e-29, 
    8.598581e-29, 8.598557e-29, 8.598522e-29, 8.598498e-29, 8.598481e-29, 
    8.598491e-29, 8.598482e-29, 8.598492e-29, 8.598497e-29, 8.598445e-29, 
    8.598474e-29, 8.59843e-29, 8.598432e-29, 8.598453e-29, 8.598432e-29, 
    8.59863e-29, 8.598635e-29, 8.598655e-29, 8.598639e-29, 8.598668e-29, 
    8.598652e-29, 8.598643e-29, 8.598608e-29, 8.5986e-29, 8.598593e-29, 
    8.598579e-29, 8.598561e-29, 8.598529e-29, 8.598501e-29, 8.598477e-29, 
    8.598479e-29, 8.598478e-29, 8.598472e-29, 8.598486e-29, 8.59847e-29, 
    8.598467e-29, 8.598474e-29, 8.598433e-29, 8.598445e-29, 8.598432e-29, 
    8.59844e-29, 8.598633e-29, 8.598624e-29, 8.598629e-29, 8.598619e-29, 
    8.598626e-29, 8.598596e-29, 8.598586e-29, 8.598544e-29, 8.598561e-29, 
    8.598533e-29, 8.598559e-29, 8.598554e-29, 8.598533e-29, 8.598557e-29, 
    8.598503e-29, 8.59854e-29, 8.598472e-29, 8.598508e-29, 8.59847e-29, 
    8.598477e-29, 8.598465e-29, 8.598454e-29, 8.598441e-29, 8.598417e-29, 
    8.598423e-29, 8.598402e-29, 8.59861e-29, 8.598597e-29, 8.598598e-29, 
    8.598585e-29, 8.598575e-29, 8.598555e-29, 8.598521e-29, 8.598534e-29, 
    8.598511e-29, 8.598506e-29, 8.598541e-29, 8.598519e-29, 8.598589e-29, 
    8.598578e-29, 8.598584e-29, 8.598609e-29, 8.598531e-29, 8.598571e-29, 
    8.598497e-29, 8.598519e-29, 8.598456e-29, 8.598487e-29, 8.598426e-29, 
    8.598399e-29, 8.598374e-29, 8.598346e-29, 8.59859e-29, 8.598599e-29, 
    8.598584e-29, 8.598563e-29, 8.598544e-29, 8.598518e-29, 8.598515e-29, 
    8.59851e-29, 8.598498e-29, 8.598487e-29, 8.598509e-29, 8.598485e-29, 
    8.598575e-29, 8.598527e-29, 8.598602e-29, 8.59858e-29, 8.598564e-29, 
    8.598571e-29, 8.598535e-29, 8.598527e-29, 8.598493e-29, 8.59851e-29, 
    8.598406e-29, 8.598452e-29, 8.598323e-29, 8.598359e-29, 8.598602e-29, 
    8.59859e-29, 8.598551e-29, 8.598569e-29, 8.598516e-29, 8.598503e-29, 
    8.598492e-29, 8.598478e-29, 8.598477e-29, 8.598468e-29, 8.598482e-29, 
    8.598469e-29, 8.598518e-29, 8.598496e-29, 8.598556e-29, 8.598541e-29, 
    8.598548e-29, 8.598555e-29, 8.598532e-29, 8.598508e-29, 8.598507e-29, 
    8.5985e-29, 8.598479e-29, 8.598516e-29, 8.5984e-29, 8.598471e-29, 
    8.598578e-29, 8.598556e-29, 8.598553e-29, 8.598562e-29, 8.598504e-29, 
    8.598525e-29, 8.598468e-29, 8.598484e-29, 8.598459e-29, 8.598471e-29, 
    8.598473e-29, 8.598489e-29, 8.598499e-29, 8.598524e-29, 8.598544e-29, 
    8.59856e-29, 8.598557e-29, 8.598539e-29, 8.598507e-29, 8.598476e-29, 
    8.598483e-29, 8.59846e-29, 8.598519e-29, 8.598495e-29, 8.598504e-29, 
    8.59848e-29, 8.598535e-29, 8.598488e-29, 8.598546e-29, 8.598541e-29, 
    8.598525e-29, 8.598494e-29, 8.598486e-29, 8.598479e-29, 8.598483e-29, 
    8.598506e-29, 8.59851e-29, 8.598525e-29, 8.59853e-29, 8.598542e-29, 
    8.598552e-29, 8.598543e-29, 8.598533e-29, 8.598506e-29, 8.598481e-29, 
    8.598454e-29, 8.598448e-29, 8.598416e-29, 8.598442e-29, 8.5984e-29, 
    8.598435e-29, 8.598373e-29, 8.598485e-29, 8.598436e-29, 8.598524e-29, 
    8.598515e-29, 8.598498e-29, 8.598459e-29, 8.59848e-29, 8.598455e-29, 
    8.59851e-29, 8.598538e-29, 8.598545e-29, 8.598559e-29, 8.598545e-29, 
    8.598547e-29, 8.598533e-29, 8.598538e-29, 8.598505e-29, 8.598522e-29, 
    8.598473e-29, 8.598455e-29, 8.598405e-29, 8.598373e-29, 8.598341e-29, 
    8.598327e-29, 8.598323e-29, 8.598321e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N_TO_SOIL2N =
  1.165102e-08, 1.170224e-08, 1.169228e-08, 1.173359e-08, 1.171068e-08, 
    1.173773e-08, 1.16614e-08, 1.170427e-08, 1.16769e-08, 1.165563e-08, 
    1.181377e-08, 1.173544e-08, 1.189512e-08, 1.184517e-08, 1.197065e-08, 
    1.188735e-08, 1.198745e-08, 1.196825e-08, 1.202603e-08, 1.200948e-08, 
    1.208339e-08, 1.203367e-08, 1.212171e-08, 1.207152e-08, 1.207937e-08, 
    1.203203e-08, 1.17512e-08, 1.180401e-08, 1.174807e-08, 1.17556e-08, 
    1.175222e-08, 1.171115e-08, 1.169045e-08, 1.16471e-08, 1.165497e-08, 
    1.168681e-08, 1.175899e-08, 1.173449e-08, 1.179623e-08, 1.179484e-08, 
    1.186358e-08, 1.183259e-08, 1.194812e-08, 1.191528e-08, 1.201017e-08, 
    1.198631e-08, 1.200905e-08, 1.200215e-08, 1.200914e-08, 1.197414e-08, 
    1.198914e-08, 1.195834e-08, 1.183839e-08, 1.187364e-08, 1.17685e-08, 
    1.170528e-08, 1.166328e-08, 1.163348e-08, 1.163769e-08, 1.164573e-08, 
    1.1687e-08, 1.17258e-08, 1.175537e-08, 1.177515e-08, 1.179464e-08, 
    1.185363e-08, 1.188485e-08, 1.195476e-08, 1.194214e-08, 1.196352e-08, 
    1.198393e-08, 1.201821e-08, 1.201257e-08, 1.202767e-08, 1.196295e-08, 
    1.200597e-08, 1.193496e-08, 1.195438e-08, 1.179994e-08, 1.17411e-08, 
    1.171609e-08, 1.169419e-08, 1.164093e-08, 1.167771e-08, 1.166322e-08, 
    1.169771e-08, 1.171963e-08, 1.170879e-08, 1.177569e-08, 1.174968e-08, 
    1.18867e-08, 1.182768e-08, 1.198155e-08, 1.194473e-08, 1.199038e-08, 
    1.196709e-08, 1.200699e-08, 1.197108e-08, 1.203329e-08, 1.204684e-08, 
    1.203758e-08, 1.207315e-08, 1.196909e-08, 1.200905e-08, 1.170848e-08, 
    1.171025e-08, 1.171849e-08, 1.168228e-08, 1.168007e-08, 1.164689e-08, 
    1.167641e-08, 1.168898e-08, 1.17209e-08, 1.173978e-08, 1.175772e-08, 
    1.179718e-08, 1.184124e-08, 1.190286e-08, 1.194712e-08, 1.197679e-08, 
    1.19586e-08, 1.197466e-08, 1.19567e-08, 1.194829e-08, 1.204177e-08, 
    1.198928e-08, 1.206803e-08, 1.206367e-08, 1.202803e-08, 1.206416e-08, 
    1.171149e-08, 1.170132e-08, 1.1666e-08, 1.169364e-08, 1.164327e-08, 
    1.167147e-08, 1.168768e-08, 1.175022e-08, 1.176396e-08, 1.177671e-08, 
    1.180187e-08, 1.183417e-08, 1.189083e-08, 1.194012e-08, 1.198512e-08, 
    1.198182e-08, 1.198298e-08, 1.199304e-08, 1.196814e-08, 1.199713e-08, 
    1.200199e-08, 1.198927e-08, 1.206309e-08, 1.2042e-08, 1.206358e-08, 
    1.204985e-08, 1.170462e-08, 1.172174e-08, 1.171249e-08, 1.172989e-08, 
    1.171763e-08, 1.177213e-08, 1.178847e-08, 1.186491e-08, 1.183354e-08, 
    1.188347e-08, 1.183861e-08, 1.184656e-08, 1.18851e-08, 1.184103e-08, 
    1.193741e-08, 1.187207e-08, 1.199343e-08, 1.192819e-08, 1.199752e-08, 
    1.198493e-08, 1.200577e-08, 1.202444e-08, 1.204793e-08, 1.209126e-08, 
    1.208123e-08, 1.211747e-08, 1.174727e-08, 1.176947e-08, 1.176751e-08, 
    1.179075e-08, 1.180794e-08, 1.184518e-08, 1.190492e-08, 1.188246e-08, 
    1.192369e-08, 1.193197e-08, 1.186932e-08, 1.190779e-08, 1.178433e-08, 
    1.180428e-08, 1.17924e-08, 1.174902e-08, 1.188763e-08, 1.18165e-08, 
    1.194785e-08, 1.190932e-08, 1.202178e-08, 1.196585e-08, 1.20757e-08, 
    1.212267e-08, 1.216686e-08, 1.221852e-08, 1.178159e-08, 1.17665e-08, 
    1.179351e-08, 1.183089e-08, 1.186557e-08, 1.191167e-08, 1.191638e-08, 
    1.192502e-08, 1.194739e-08, 1.19662e-08, 1.192775e-08, 1.197091e-08, 
    1.180891e-08, 1.189381e-08, 1.17608e-08, 1.180085e-08, 1.182869e-08, 
    1.181647e-08, 1.187989e-08, 1.189483e-08, 1.195557e-08, 1.192417e-08, 
    1.211108e-08, 1.202839e-08, 1.225784e-08, 1.219372e-08, 1.176123e-08, 
    1.178153e-08, 1.185221e-08, 1.181858e-08, 1.191474e-08, 1.193841e-08, 
    1.195765e-08, 1.198225e-08, 1.198491e-08, 1.199948e-08, 1.19756e-08, 
    1.199854e-08, 1.191176e-08, 1.195054e-08, 1.184413e-08, 1.187003e-08, 
    1.185811e-08, 1.184504e-08, 1.188538e-08, 1.192836e-08, 1.192927e-08, 
    1.194305e-08, 1.198189e-08, 1.191513e-08, 1.212176e-08, 1.199415e-08, 
    1.180368e-08, 1.184279e-08, 1.184838e-08, 1.183323e-08, 1.193604e-08, 
    1.189879e-08, 1.199912e-08, 1.197201e-08, 1.201644e-08, 1.199436e-08, 
    1.199111e-08, 1.196275e-08, 1.19451e-08, 1.19005e-08, 1.18642e-08, 
    1.183542e-08, 1.184212e-08, 1.187373e-08, 1.193099e-08, 1.198515e-08, 
    1.197328e-08, 1.201306e-08, 1.190777e-08, 1.195192e-08, 1.193486e-08, 
    1.197935e-08, 1.188186e-08, 1.196488e-08, 1.186064e-08, 1.186978e-08, 
    1.189805e-08, 1.195492e-08, 1.19675e-08, 1.198093e-08, 1.197264e-08, 
    1.193244e-08, 1.192585e-08, 1.189736e-08, 1.18895e-08, 1.186779e-08, 
    1.184981e-08, 1.186623e-08, 1.188348e-08, 1.193245e-08, 1.197659e-08, 
    1.202471e-08, 1.203648e-08, 1.209271e-08, 1.204694e-08, 1.212247e-08, 
    1.205826e-08, 1.21694e-08, 1.196969e-08, 1.205637e-08, 1.189933e-08, 
    1.191625e-08, 1.194685e-08, 1.201703e-08, 1.197914e-08, 1.202345e-08, 
    1.192559e-08, 1.187482e-08, 1.186168e-08, 1.183717e-08, 1.186224e-08, 
    1.18602e-08, 1.188419e-08, 1.187648e-08, 1.193408e-08, 1.190314e-08, 
    1.199103e-08, 1.20231e-08, 1.211367e-08, 1.21692e-08, 1.222571e-08, 
    1.225066e-08, 1.225825e-08, 1.226143e-08 ;

 SOIL1N_TO_SOIL3N =
  1.382354e-10, 1.388434e-10, 1.387252e-10, 1.392155e-10, 1.389435e-10, 
    1.392646e-10, 1.383587e-10, 1.388675e-10, 1.385427e-10, 1.382901e-10, 
    1.401671e-10, 1.392374e-10, 1.411328e-10, 1.405399e-10, 1.420293e-10, 
    1.410406e-10, 1.422287e-10, 1.420008e-10, 1.426867e-10, 1.424902e-10, 
    1.433676e-10, 1.427774e-10, 1.438223e-10, 1.432266e-10, 1.433198e-10, 
    1.427579e-10, 1.394245e-10, 1.400514e-10, 1.393873e-10, 1.394767e-10, 
    1.394366e-10, 1.389491e-10, 1.387035e-10, 1.381889e-10, 1.382824e-10, 
    1.386603e-10, 1.395169e-10, 1.392261e-10, 1.39959e-10, 1.399425e-10, 
    1.407584e-10, 1.403905e-10, 1.417619e-10, 1.413721e-10, 1.424984e-10, 
    1.422151e-10, 1.424851e-10, 1.424032e-10, 1.424862e-10, 1.420707e-10, 
    1.422487e-10, 1.418832e-10, 1.404594e-10, 1.408779e-10, 1.396298e-10, 
    1.388794e-10, 1.38381e-10, 1.380273e-10, 1.380773e-10, 1.381726e-10, 
    1.386625e-10, 1.39123e-10, 1.39474e-10, 1.397088e-10, 1.399401e-10, 
    1.406403e-10, 1.410109e-10, 1.418407e-10, 1.416909e-10, 1.419446e-10, 
    1.42187e-10, 1.425939e-10, 1.425269e-10, 1.427062e-10, 1.419379e-10, 
    1.424485e-10, 1.416056e-10, 1.418362e-10, 1.40003e-10, 1.393046e-10, 
    1.390077e-10, 1.387479e-10, 1.381157e-10, 1.385523e-10, 1.383802e-10, 
    1.387896e-10, 1.390498e-10, 1.389211e-10, 1.397152e-10, 1.394065e-10, 
    1.410329e-10, 1.403323e-10, 1.421587e-10, 1.417217e-10, 1.422635e-10, 
    1.41987e-10, 1.424607e-10, 1.420344e-10, 1.427729e-10, 1.429337e-10, 
    1.428238e-10, 1.432459e-10, 1.420107e-10, 1.424851e-10, 1.389175e-10, 
    1.389385e-10, 1.390362e-10, 1.386065e-10, 1.385802e-10, 1.381864e-10, 
    1.385368e-10, 1.38686e-10, 1.390648e-10, 1.392889e-10, 1.395019e-10, 
    1.399702e-10, 1.404932e-10, 1.412246e-10, 1.4175e-10, 1.421022e-10, 
    1.418862e-10, 1.420769e-10, 1.418637e-10, 1.417638e-10, 1.428734e-10, 
    1.422504e-10, 1.431852e-10, 1.431335e-10, 1.427104e-10, 1.431393e-10, 
    1.389532e-10, 1.388324e-10, 1.384132e-10, 1.387413e-10, 1.381435e-10, 
    1.384781e-10, 1.386705e-10, 1.394129e-10, 1.39576e-10, 1.397273e-10, 
    1.40026e-10, 1.404093e-10, 1.410818e-10, 1.416669e-10, 1.422011e-10, 
    1.421619e-10, 1.421757e-10, 1.42295e-10, 1.419995e-10, 1.423436e-10, 
    1.424013e-10, 1.422503e-10, 1.431266e-10, 1.428762e-10, 1.431324e-10, 
    1.429694e-10, 1.388717e-10, 1.390749e-10, 1.389651e-10, 1.391716e-10, 
    1.390261e-10, 1.396729e-10, 1.398668e-10, 1.407742e-10, 1.404018e-10, 
    1.409945e-10, 1.40462e-10, 1.405563e-10, 1.410138e-10, 1.404908e-10, 
    1.416347e-10, 1.408592e-10, 1.422997e-10, 1.415253e-10, 1.423482e-10, 
    1.421988e-10, 1.424462e-10, 1.426678e-10, 1.429466e-10, 1.43461e-10, 
    1.433419e-10, 1.43772e-10, 1.393778e-10, 1.396414e-10, 1.396182e-10, 
    1.398939e-10, 1.400979e-10, 1.4054e-10, 1.412491e-10, 1.409824e-10, 
    1.414719e-10, 1.415702e-10, 1.408265e-10, 1.412831e-10, 1.398177e-10, 
    1.400545e-10, 1.399135e-10, 1.393986e-10, 1.410439e-10, 1.401995e-10, 
    1.417587e-10, 1.413013e-10, 1.426362e-10, 1.419723e-10, 1.432763e-10, 
    1.438338e-10, 1.443584e-10, 1.449715e-10, 1.397852e-10, 1.396061e-10, 
    1.399268e-10, 1.403704e-10, 1.40782e-10, 1.413292e-10, 1.413852e-10, 
    1.414877e-10, 1.417532e-10, 1.419764e-10, 1.415201e-10, 1.420324e-10, 
    1.401095e-10, 1.411172e-10, 1.395384e-10, 1.400138e-10, 1.403442e-10, 
    1.401993e-10, 1.40952e-10, 1.411294e-10, 1.418502e-10, 1.414776e-10, 
    1.436962e-10, 1.427146e-10, 1.454383e-10, 1.446772e-10, 1.395435e-10, 
    1.397846e-10, 1.406234e-10, 1.402243e-10, 1.413657e-10, 1.416466e-10, 
    1.41875e-10, 1.42167e-10, 1.421985e-10, 1.423715e-10, 1.42088e-10, 
    1.423603e-10, 1.413303e-10, 1.417906e-10, 1.405275e-10, 1.40835e-10, 
    1.406935e-10, 1.405384e-10, 1.410172e-10, 1.415273e-10, 1.415382e-10, 
    1.417017e-10, 1.421627e-10, 1.413703e-10, 1.438229e-10, 1.423083e-10, 
    1.400474e-10, 1.405117e-10, 1.40578e-10, 1.403981e-10, 1.416185e-10, 
    1.411763e-10, 1.423673e-10, 1.420454e-10, 1.425728e-10, 1.423107e-10, 
    1.422722e-10, 1.419356e-10, 1.41726e-10, 1.411966e-10, 1.407658e-10, 
    1.404242e-10, 1.405036e-10, 1.408789e-10, 1.415585e-10, 1.422014e-10, 
    1.420605e-10, 1.425327e-10, 1.412829e-10, 1.41807e-10, 1.416045e-10, 
    1.421326e-10, 1.409754e-10, 1.419609e-10, 1.407235e-10, 1.408319e-10, 
    1.411675e-10, 1.418426e-10, 1.419919e-10, 1.421513e-10, 1.420529e-10, 
    1.415757e-10, 1.414975e-10, 1.411594e-10, 1.41066e-10, 1.408083e-10, 
    1.40595e-10, 1.407899e-10, 1.409946e-10, 1.415759e-10, 1.420998e-10, 
    1.426709e-10, 1.428107e-10, 1.434781e-10, 1.429348e-10, 1.438313e-10, 
    1.430692e-10, 1.443885e-10, 1.420179e-10, 1.430467e-10, 1.411828e-10, 
    1.413836e-10, 1.417468e-10, 1.425798e-10, 1.421301e-10, 1.426561e-10, 
    1.414945e-10, 1.408918e-10, 1.407359e-10, 1.40445e-10, 1.407425e-10, 
    1.407183e-10, 1.410031e-10, 1.409116e-10, 1.415952e-10, 1.41228e-10, 
    1.422712e-10, 1.426519e-10, 1.43727e-10, 1.44386e-10, 1.450569e-10, 
    1.453531e-10, 1.454432e-10, 1.454809e-10 ;

 SOIL1N_vr =
  2.497425, 2.497418, 2.497419, 2.497414, 2.497417, 2.497413, 2.497423, 
    2.497418, 2.497421, 2.497424, 2.497403, 2.497414, 2.497393, 2.497399, 
    2.497383, 2.497394, 2.49738, 2.497383, 2.497375, 2.497378, 2.497368, 
    2.497375, 2.497363, 2.49737, 2.497369, 2.497375, 2.497411, 2.497405, 
    2.497412, 2.497411, 2.497411, 2.497417, 2.497419, 2.497425, 2.497424, 
    2.49742, 2.497411, 2.497414, 2.497406, 2.497406, 2.497397, 2.497401, 
    2.497386, 2.49739, 2.497378, 2.497381, 2.497378, 2.497379, 2.497378, 
    2.497382, 2.49738, 2.497384, 2.4974, 2.497396, 2.497409, 2.497417, 
    2.497423, 2.497427, 2.497427, 2.497425, 2.49742, 2.497415, 2.497411, 
    2.497408, 2.497406, 2.497398, 2.497394, 2.497385, 2.497386, 2.497384, 
    2.497381, 2.497376, 2.497377, 2.497375, 2.497384, 2.497378, 2.497387, 
    2.497385, 2.497405, 2.497413, 2.497416, 2.497419, 2.497426, 2.497421, 
    2.497423, 2.497418, 2.497416, 2.497417, 2.497408, 2.497412, 2.497394, 
    2.497401, 2.497381, 2.497386, 2.49738, 2.497383, 2.497378, 2.497383, 
    2.497375, 2.497373, 2.497374, 2.497369, 2.497383, 2.497378, 2.497417, 
    2.497417, 2.497416, 2.497421, 2.497421, 2.497425, 2.497421, 2.49742, 
    2.497416, 2.497413, 2.497411, 2.497406, 2.4974, 2.497392, 2.497386, 
    2.497382, 2.497384, 2.497382, 2.497385, 2.497386, 2.497373, 2.49738, 
    2.49737, 2.49737, 2.497375, 2.49737, 2.497417, 2.497418, 2.497423, 
    2.497419, 2.497426, 2.497422, 2.49742, 2.497411, 2.49741, 2.497408, 
    2.497405, 2.497401, 2.497393, 2.497387, 2.497381, 2.497381, 2.497381, 
    2.49738, 2.497383, 2.497379, 2.497379, 2.49738, 2.497371, 2.497373, 
    2.497371, 2.497372, 2.497418, 2.497415, 2.497416, 2.497414, 2.497416, 
    2.497409, 2.497406, 2.497396, 2.497401, 2.497394, 2.4974, 2.497399, 
    2.497394, 2.4974, 2.497387, 2.497396, 2.49738, 2.497388, 2.497379, 
    2.497381, 2.497378, 2.497376, 2.497373, 2.497367, 2.497368, 2.497364, 
    2.497412, 2.497409, 2.497409, 2.497406, 2.497404, 2.497399, 2.497391, 
    2.497394, 2.497389, 2.497388, 2.497396, 2.497391, 2.497407, 2.497405, 
    2.497406, 2.497412, 2.497394, 2.497403, 2.497386, 2.497391, 2.497376, 
    2.497383, 2.497369, 2.497363, 2.497357, 2.49735, 2.497407, 2.49741, 
    2.497406, 2.497401, 2.497396, 2.497391, 2.49739, 2.497389, 2.497386, 
    2.497383, 2.497388, 2.497383, 2.497404, 2.497393, 2.49741, 2.497405, 
    2.497401, 2.497403, 2.497395, 2.497393, 2.497385, 2.497389, 2.497365, 
    2.497375, 2.497345, 2.497354, 2.49741, 2.497407, 2.497398, 2.497403, 
    2.49739, 2.497387, 2.497384, 2.497381, 2.497381, 2.497379, 2.497382, 
    2.497379, 2.497391, 2.497385, 2.497399, 2.497396, 2.497397, 2.497399, 
    2.497394, 2.497388, 2.497388, 2.497386, 2.497381, 2.49739, 2.497363, 
    2.49738, 2.497405, 2.4974, 2.497399, 2.497401, 2.497387, 2.497392, 
    2.497379, 2.497383, 2.497377, 2.49738, 2.49738, 2.497384, 2.497386, 
    2.497392, 2.497397, 2.497401, 2.4974, 2.497396, 2.497388, 2.497381, 
    2.497382, 2.497377, 2.497391, 2.497385, 2.497387, 2.497382, 2.497394, 
    2.497383, 2.497397, 2.497396, 2.497392, 2.497385, 2.497383, 2.497381, 
    2.497382, 2.497388, 2.497389, 2.497392, 2.497393, 2.497396, 2.497399, 
    2.497396, 2.497394, 2.497388, 2.497382, 2.497376, 2.497374, 2.497367, 
    2.497373, 2.497363, 2.497371, 2.497357, 2.497383, 2.497371, 2.497392, 
    2.49739, 2.497386, 2.497377, 2.497382, 2.497376, 2.497389, 2.497395, 
    2.497397, 2.4974, 2.497397, 2.497397, 2.497394, 2.497395, 2.497387, 
    2.497391, 2.49738, 2.497376, 2.497364, 2.497357, 2.49735, 2.497346, 
    2.497345, 2.497345,
  2.497625, 2.497616, 2.497618, 2.497611, 2.497615, 2.49761, 2.497623, 
    2.497616, 2.49762, 2.497624, 2.497597, 2.49761, 2.497583, 2.497591, 
    2.49757, 2.497584, 2.497567, 2.49757, 2.49756, 2.497563, 2.49755, 
    2.497559, 2.497544, 2.497552, 2.497551, 2.497559, 2.497607, 2.497598, 
    2.497608, 2.497607, 2.497607, 2.497615, 2.497618, 2.497626, 2.497624, 
    2.497619, 2.497606, 2.497611, 2.4976, 2.4976, 2.497588, 2.497593, 
    2.497574, 2.497579, 2.497563, 2.497567, 2.497563, 2.497564, 2.497563, 
    2.497569, 2.497566, 2.497572, 2.497592, 2.497586, 2.497605, 2.497616, 
    2.497623, 2.497628, 2.497627, 2.497626, 2.497619, 2.497612, 2.497607, 
    2.497603, 2.4976, 2.49759, 2.497585, 2.497572, 2.497575, 2.497571, 
    2.497567, 2.497561, 2.497562, 2.49756, 2.497571, 2.497564, 2.497576, 
    2.497572, 2.497599, 2.497609, 2.497614, 2.497617, 2.497627, 2.49762, 
    2.497623, 2.497617, 2.497613, 2.497615, 2.497603, 2.497608, 2.497584, 
    2.497594, 2.497568, 2.497574, 2.497566, 2.49757, 2.497563, 2.49757, 
    2.497559, 2.497557, 2.497558, 2.497552, 2.49757, 2.497563, 2.497615, 
    2.497615, 2.497613, 2.49762, 2.49762, 2.497626, 2.497621, 2.497618, 
    2.497613, 2.49761, 2.497607, 2.4976, 2.497592, 2.497581, 2.497574, 
    2.497569, 2.497572, 2.497569, 2.497572, 2.497574, 2.497557, 2.497566, 
    2.497553, 2.497554, 2.49756, 2.497554, 2.497614, 2.497616, 2.497622, 
    2.497617, 2.497626, 2.497621, 2.497619, 2.497608, 2.497605, 2.497603, 
    2.497599, 2.497593, 2.497583, 2.497575, 2.497567, 2.497568, 2.497568, 
    2.497566, 2.49757, 2.497565, 2.497564, 2.497566, 2.497554, 2.497557, 
    2.497554, 2.497556, 2.497616, 2.497613, 2.497614, 2.497611, 2.497613, 
    2.497604, 2.497601, 2.497588, 2.497593, 2.497585, 2.497592, 2.497591, 
    2.497584, 2.497592, 2.497576, 2.497587, 2.497566, 2.497577, 2.497565, 
    2.497567, 2.497564, 2.497561, 2.497556, 2.497549, 2.497551, 2.497545, 
    2.497608, 2.497604, 2.497605, 2.497601, 2.497598, 2.497591, 2.497581, 
    2.497585, 2.497578, 2.497576, 2.497587, 2.497581, 2.497602, 2.497598, 
    2.497601, 2.497608, 2.497584, 2.497596, 2.497574, 2.49758, 2.497561, 
    2.497571, 2.497552, 2.497544, 2.497536, 2.497527, 2.497602, 2.497605, 
    2.4976, 2.497594, 2.497588, 2.49758, 2.497579, 2.497578, 2.497574, 
    2.497571, 2.497577, 2.49757, 2.497598, 2.497583, 2.497606, 2.497599, 
    2.497594, 2.497596, 2.497585, 2.497583, 2.497572, 2.497578, 2.497545, 
    2.49756, 2.49752, 2.497531, 2.497606, 2.497602, 2.49759, 2.497596, 
    2.497579, 2.497575, 2.497572, 2.497568, 2.497567, 2.497565, 2.497569, 
    2.497565, 2.49758, 2.497573, 2.497591, 2.497587, 2.497589, 2.497591, 
    2.497584, 2.497577, 2.497577, 2.497574, 2.497568, 2.497579, 2.497544, 
    2.497566, 2.497598, 2.497592, 2.497591, 2.497593, 2.497576, 2.497582, 
    2.497565, 2.49757, 2.497562, 2.497566, 2.497566, 2.497571, 2.497574, 
    2.497582, 2.497588, 2.497593, 2.497592, 2.497586, 2.497576, 2.497567, 
    2.497569, 2.497562, 2.497581, 2.497573, 2.497576, 2.497568, 2.497585, 
    2.497571, 2.497589, 2.497587, 2.497582, 2.497572, 2.49757, 2.497568, 
    2.497569, 2.497576, 2.497577, 2.497582, 2.497584, 2.497587, 2.497591, 
    2.497588, 2.497585, 2.497576, 2.497569, 2.497561, 2.497558, 2.497549, 
    2.497556, 2.497544, 2.497555, 2.497535, 2.49757, 2.497555, 2.497582, 
    2.497579, 2.497574, 2.497562, 2.497568, 2.497561, 2.497577, 2.497586, 
    2.497588, 2.497593, 2.497588, 2.497589, 2.497585, 2.497586, 2.497576, 
    2.497581, 2.497566, 2.497561, 2.497545, 2.497535, 2.497526, 2.497522, 
    2.49752, 2.49752,
  2.49784, 2.497831, 2.497833, 2.497825, 2.497829, 2.497824, 2.497838, 
    2.49783, 2.497835, 2.497839, 2.49781, 2.497825, 2.497795, 2.497804, 
    2.497781, 2.497797, 2.497778, 2.497782, 2.497771, 2.497774, 2.497761, 
    2.49777, 2.497753, 2.497763, 2.497761, 2.49777, 2.497822, 2.497812, 
    2.497822, 2.497821, 2.497822, 2.497829, 2.497833, 2.497841, 2.497839, 
    2.497834, 2.49782, 2.497825, 2.497813, 2.497814, 2.497801, 2.497807, 
    2.497785, 2.497792, 2.497774, 2.497778, 2.497774, 2.497776, 2.497774, 
    2.497781, 2.497778, 2.497784, 2.497806, 2.497799, 2.497818, 2.49783, 
    2.497838, 2.497844, 2.497843, 2.497841, 2.497834, 2.497826, 2.497821, 
    2.497817, 2.497814, 2.497803, 2.497797, 2.497784, 2.497787, 2.497782, 
    2.497779, 2.497772, 2.497774, 2.497771, 2.497783, 2.497775, 2.497788, 
    2.497784, 2.497813, 2.497824, 2.497828, 2.497832, 2.497842, 2.497835, 
    2.497838, 2.497832, 2.497828, 2.49783, 2.497817, 2.497822, 2.497797, 
    2.497808, 2.497779, 2.497786, 2.497778, 2.497782, 2.497775, 2.497781, 
    2.49777, 2.497767, 2.497769, 2.497762, 2.497782, 2.497774, 2.49783, 
    2.497829, 2.497828, 2.497834, 2.497835, 2.497841, 2.497836, 2.497833, 
    2.497827, 2.497824, 2.497821, 2.497813, 2.497805, 2.497794, 2.497786, 
    2.49778, 2.497783, 2.497781, 2.497784, 2.497785, 2.497768, 2.497778, 
    2.497763, 2.497764, 2.497771, 2.497764, 2.497829, 2.497831, 2.497838, 
    2.497832, 2.497842, 2.497837, 2.497833, 2.497822, 2.497819, 2.497817, 
    2.497813, 2.497807, 2.497796, 2.497787, 2.497779, 2.497779, 2.497779, 
    2.497777, 2.497782, 2.497777, 2.497776, 2.497778, 2.497764, 2.497768, 
    2.497764, 2.497767, 2.49783, 2.497827, 2.497829, 2.497826, 2.497828, 
    2.497818, 2.497815, 2.497801, 2.497807, 2.497797, 2.497806, 2.497804, 
    2.497797, 2.497805, 2.497787, 2.497799, 2.497777, 2.497789, 2.497776, 
    2.497779, 2.497775, 2.497771, 2.497767, 2.497759, 2.497761, 2.497754, 
    2.497823, 2.497818, 2.497819, 2.497814, 2.497811, 2.497804, 2.497793, 
    2.497797, 2.49779, 2.497788, 2.4978, 2.497793, 2.497816, 2.497812, 
    2.497814, 2.497822, 2.497797, 2.49781, 2.497786, 2.497792, 2.497772, 
    2.497782, 2.497762, 2.497753, 2.497745, 2.497736, 2.497816, 2.497819, 
    2.497814, 2.497807, 2.497801, 2.497792, 2.497791, 2.49779, 2.497786, 
    2.497782, 2.497789, 2.497781, 2.497811, 2.497795, 2.49782, 2.497813, 
    2.497808, 2.49781, 2.497798, 2.497795, 2.497784, 2.49779, 2.497756, 
    2.497771, 2.497729, 2.49774, 2.49782, 2.497816, 2.497803, 2.497809, 
    2.497792, 2.497787, 2.497784, 2.497779, 2.497779, 2.497776, 2.49778, 
    2.497776, 2.497792, 2.497785, 2.497805, 2.4978, 2.497802, 2.497804, 
    2.497797, 2.497789, 2.497789, 2.497786, 2.497779, 2.497792, 2.497753, 
    2.497777, 2.497812, 2.497805, 2.497804, 2.497807, 2.497788, 2.497795, 
    2.497776, 2.497781, 2.497773, 2.497777, 2.497777, 2.497783, 2.497786, 
    2.497794, 2.497801, 2.497806, 2.497805, 2.497799, 2.497789, 2.497779, 
    2.497781, 2.497773, 2.497793, 2.497785, 2.497788, 2.49778, 2.497798, 
    2.497782, 2.497802, 2.4978, 2.497795, 2.497784, 2.497782, 2.497779, 
    2.497781, 2.497788, 2.49779, 2.497795, 2.497796, 2.4978, 2.497803, 
    2.497801, 2.497797, 2.497788, 2.49778, 2.497771, 2.497769, 2.497759, 
    2.497767, 2.497753, 2.497765, 2.497745, 2.497782, 2.497766, 2.497794, 
    2.497791, 2.497786, 2.497773, 2.49778, 2.497772, 2.49779, 2.497799, 
    2.497801, 2.497806, 2.497801, 2.497802, 2.497797, 2.497799, 2.497788, 
    2.497794, 2.497777, 2.497772, 2.497755, 2.497745, 2.497734, 2.49773, 
    2.497728, 2.497728,
  2.498012, 2.498003, 2.498005, 2.497997, 2.498001, 2.497997, 2.49801, 
    2.498003, 2.498008, 2.498012, 2.497983, 2.497997, 2.497968, 2.497977, 
    2.497954, 2.497969, 2.497951, 2.497954, 2.497944, 2.497947, 2.497933, 
    2.497942, 2.497926, 2.497936, 2.497934, 2.497943, 2.497994, 2.497984, 
    2.497995, 2.497993, 2.497994, 2.498001, 2.498005, 2.498013, 2.498012, 
    2.498006, 2.497993, 2.497997, 2.497986, 2.497986, 2.497973, 2.497979, 
    2.497958, 2.497964, 2.497947, 2.497951, 2.497947, 2.497948, 2.497947, 
    2.497953, 2.497951, 2.497956, 2.497978, 2.497972, 2.497991, 2.498003, 
    2.49801, 2.498016, 2.498015, 2.498013, 2.498006, 2.497999, 2.497993, 
    2.49799, 2.497986, 2.497975, 2.49797, 2.497957, 2.497959, 2.497955, 
    2.497952, 2.497945, 2.497946, 2.497943, 2.497955, 2.497947, 2.49796, 
    2.497957, 2.497985, 2.497996, 2.498, 2.498004, 2.498014, 2.498008, 
    2.49801, 2.498004, 2.498, 2.498002, 2.49799, 2.497994, 2.497969, 2.49798, 
    2.497952, 2.497959, 2.49795, 2.497955, 2.497947, 2.497954, 2.497942, 
    2.49794, 2.497942, 2.497935, 2.497954, 2.497947, 2.498002, 2.498002, 
    2.498, 2.498007, 2.498007, 2.498013, 2.498008, 2.498005, 2.498, 2.497996, 
    2.497993, 2.497986, 2.497977, 2.497966, 2.497958, 2.497953, 2.497956, 
    2.497953, 2.497957, 2.497958, 2.497941, 2.497951, 2.497936, 2.497937, 
    2.497943, 2.497937, 2.498001, 2.498003, 2.49801, 2.498005, 2.498014, 
    2.498009, 2.498006, 2.497994, 2.497992, 2.497989, 2.497985, 2.497979, 
    2.497968, 2.497959, 2.497951, 2.497952, 2.497952, 2.49795, 2.497954, 
    2.497949, 2.497948, 2.497951, 2.497937, 2.497941, 2.497937, 2.497939, 
    2.498003, 2.497999, 2.498001, 2.497998, 2.498, 2.49799, 2.497987, 
    2.497973, 2.497979, 2.49797, 2.497978, 2.497977, 2.49797, 2.497977, 
    2.49796, 2.497972, 2.49795, 2.497962, 2.497949, 2.497951, 2.497947, 
    2.497944, 2.49794, 2.497932, 2.497934, 2.497927, 2.497995, 2.497991, 
    2.497991, 2.497987, 2.497984, 2.497977, 2.497966, 2.49797, 2.497962, 
    2.497961, 2.497972, 2.497965, 2.497988, 2.497984, 2.497987, 2.497994, 
    2.497969, 2.497982, 2.497958, 2.497965, 2.497945, 2.497955, 2.497935, 
    2.497926, 2.497918, 2.497909, 2.497988, 2.497991, 2.497986, 2.497979, 
    2.497973, 2.497965, 2.497964, 2.497962, 2.497958, 2.497955, 2.497962, 
    2.497954, 2.497983, 2.497968, 2.497992, 2.497985, 2.49798, 2.497982, 
    2.497971, 2.497968, 2.497957, 2.497962, 2.497928, 2.497943, 2.497901, 
    2.497913, 2.497992, 2.497988, 2.497976, 2.497982, 2.497964, 2.49796, 
    2.497956, 2.497952, 2.497951, 2.497949, 2.497953, 2.497949, 2.497965, 
    2.497957, 2.497977, 2.497972, 2.497974, 2.497977, 2.497969, 2.497962, 
    2.497962, 2.497959, 2.497952, 2.497964, 2.497926, 2.49795, 2.497984, 
    2.497977, 2.497976, 2.497979, 2.49796, 2.497967, 2.497949, 2.497954, 
    2.497946, 2.49795, 2.49795, 2.497955, 2.497959, 2.497967, 2.497973, 
    2.497979, 2.497977, 2.497972, 2.497961, 2.497951, 2.497953, 2.497946, 
    2.497965, 2.497957, 2.49796, 2.497952, 2.49797, 2.497955, 2.497974, 
    2.497972, 2.497967, 2.497957, 2.497954, 2.497952, 2.497953, 2.497961, 
    2.497962, 2.497967, 2.497969, 2.497973, 2.497976, 2.497973, 2.49797, 
    2.497961, 2.497953, 2.497944, 2.497942, 2.497931, 2.49794, 2.497926, 
    2.497938, 2.497918, 2.497954, 2.497938, 2.497967, 2.497964, 2.497958, 
    2.497945, 2.497952, 2.497944, 2.497962, 2.497971, 2.497974, 2.497978, 
    2.497974, 2.497974, 2.49797, 2.497971, 2.497961, 2.497966, 2.49795, 
    2.497944, 2.497928, 2.497918, 2.497907, 2.497903, 2.497901, 2.497901,
  2.498213, 2.498205, 2.498206, 2.4982, 2.498204, 2.498199, 2.498211, 
    2.498204, 2.498209, 2.498212, 2.498187, 2.498199, 2.498173, 2.498182, 
    2.498161, 2.498175, 2.498158, 2.498162, 2.498152, 2.498155, 2.498143, 
    2.498151, 2.498137, 2.498145, 2.498143, 2.498151, 2.498197, 2.498188, 
    2.498197, 2.498196, 2.498197, 2.498203, 2.498207, 2.498214, 2.498212, 
    2.498207, 2.498196, 2.498199, 2.498189, 2.49819, 2.498178, 2.498184, 
    2.498165, 2.49817, 2.498155, 2.498159, 2.498155, 2.498156, 2.498155, 
    2.498161, 2.498158, 2.498163, 2.498183, 2.498177, 2.498194, 2.498204, 
    2.498211, 2.498216, 2.498215, 2.498214, 2.498207, 2.498201, 2.498196, 
    2.498193, 2.49819, 2.49818, 2.498175, 2.498164, 2.498166, 2.498162, 
    2.498159, 2.498153, 2.498154, 2.498152, 2.498163, 2.498155, 2.498167, 
    2.498164, 2.498189, 2.498199, 2.498203, 2.498206, 2.498215, 2.498209, 
    2.498211, 2.498205, 2.498202, 2.498204, 2.498193, 2.498197, 2.498175, 
    2.498184, 2.498159, 2.498165, 2.498158, 2.498162, 2.498155, 2.498161, 
    2.498151, 2.498149, 2.49815, 2.498144, 2.498161, 2.498155, 2.498204, 
    2.498204, 2.498202, 2.498208, 2.498208, 2.498214, 2.498209, 2.498207, 
    2.498202, 2.498199, 2.498196, 2.498189, 2.498182, 2.498172, 2.498165, 
    2.49816, 2.498163, 2.498161, 2.498163, 2.498165, 2.49815, 2.498158, 
    2.498145, 2.498146, 2.498152, 2.498146, 2.498203, 2.498205, 2.498211, 
    2.498206, 2.498214, 2.49821, 2.498207, 2.498197, 2.498195, 2.498193, 
    2.498188, 2.498183, 2.498174, 2.498166, 2.498159, 2.498159, 2.498159, 
    2.498158, 2.498162, 2.498157, 2.498156, 2.498158, 2.498146, 2.49815, 
    2.498146, 2.498148, 2.498204, 2.498202, 2.498203, 2.4982, 2.498202, 
    2.498194, 2.498191, 2.498178, 2.498183, 2.498175, 2.498183, 2.498181, 
    2.498175, 2.498182, 2.498167, 2.498177, 2.498158, 2.498168, 2.498157, 
    2.498159, 2.498155, 2.498152, 2.498149, 2.498142, 2.498143, 2.498137, 
    2.498198, 2.498194, 2.498194, 2.49819, 2.498188, 2.498182, 2.498172, 
    2.498176, 2.498169, 2.498168, 2.498178, 2.498171, 2.498191, 2.498188, 
    2.49819, 2.498197, 2.498175, 2.498186, 2.498165, 2.498171, 2.498153, 
    2.498162, 2.498144, 2.498136, 2.498129, 2.498121, 2.498192, 2.498194, 
    2.49819, 2.498184, 2.498178, 2.498171, 2.49817, 2.498168, 2.498165, 
    2.498162, 2.498168, 2.498161, 2.498188, 2.498174, 2.498195, 2.498189, 
    2.498184, 2.498186, 2.498176, 2.498173, 2.498164, 2.498169, 2.498138, 
    2.498152, 2.498114, 2.498125, 2.498195, 2.498192, 2.49818, 2.498186, 
    2.49817, 2.498166, 2.498163, 2.498159, 2.498159, 2.498157, 2.49816, 
    2.498157, 2.498171, 2.498164, 2.498182, 2.498178, 2.498179, 2.498182, 
    2.498175, 2.498168, 2.498168, 2.498166, 2.498159, 2.49817, 2.498137, 
    2.498157, 2.498188, 2.498182, 2.498181, 2.498183, 2.498167, 2.498173, 
    2.498157, 2.498161, 2.498154, 2.498157, 2.498158, 2.498163, 2.498165, 
    2.498173, 2.498178, 2.498183, 2.498182, 2.498177, 2.498168, 2.498159, 
    2.498161, 2.498154, 2.498171, 2.498164, 2.498167, 2.49816, 2.498176, 
    2.498162, 2.498179, 2.498178, 2.498173, 2.498164, 2.498162, 2.498159, 
    2.498161, 2.498167, 2.498168, 2.498173, 2.498174, 2.498178, 2.498181, 
    2.498178, 2.498175, 2.498167, 2.49816, 2.498152, 2.49815, 2.498141, 
    2.498149, 2.498137, 2.498147, 2.498129, 2.498161, 2.498147, 2.498173, 
    2.49817, 2.498165, 2.498154, 2.49816, 2.498152, 2.498168, 2.498177, 
    2.498179, 2.498183, 2.498179, 2.498179, 2.498175, 2.498177, 2.498167, 
    2.498172, 2.498158, 2.498153, 2.498138, 2.498129, 2.49812, 2.498116, 
    2.498114, 2.498114,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1_HR_S2 =
  6.139984e-08, 6.166982e-08, 6.161733e-08, 6.183509e-08, 6.171429e-08, 
    6.185687e-08, 6.145457e-08, 6.168054e-08, 6.153628e-08, 6.142414e-08, 
    6.225768e-08, 6.18448e-08, 6.268651e-08, 6.24232e-08, 6.308463e-08, 
    6.264554e-08, 6.317316e-08, 6.307195e-08, 6.337655e-08, 6.328928e-08, 
    6.36789e-08, 6.341682e-08, 6.388085e-08, 6.361631e-08, 6.365769e-08, 
    6.340817e-08, 6.192788e-08, 6.220628e-08, 6.191139e-08, 6.195108e-08, 
    6.193327e-08, 6.171678e-08, 6.160769e-08, 6.13792e-08, 6.142068e-08, 
    6.15885e-08, 6.196894e-08, 6.183979e-08, 6.216526e-08, 6.21579e-08, 
    6.252024e-08, 6.235687e-08, 6.296585e-08, 6.279277e-08, 6.329292e-08, 
    6.316714e-08, 6.328702e-08, 6.325067e-08, 6.328749e-08, 6.310302e-08, 
    6.318206e-08, 6.301973e-08, 6.238747e-08, 6.257329e-08, 6.201908e-08, 
    6.168585e-08, 6.146448e-08, 6.130741e-08, 6.132962e-08, 6.137195e-08, 
    6.158948e-08, 6.1794e-08, 6.194986e-08, 6.205412e-08, 6.215684e-08, 
    6.246781e-08, 6.263237e-08, 6.300085e-08, 6.293435e-08, 6.304701e-08, 
    6.315463e-08, 6.333532e-08, 6.330558e-08, 6.338519e-08, 6.304403e-08, 
    6.327077e-08, 6.289647e-08, 6.299884e-08, 6.21848e-08, 6.187463e-08, 
    6.174282e-08, 6.162742e-08, 6.134669e-08, 6.154056e-08, 6.146414e-08, 
    6.164594e-08, 6.176148e-08, 6.170433e-08, 6.205697e-08, 6.191988e-08, 
    6.264213e-08, 6.233103e-08, 6.314207e-08, 6.2948e-08, 6.318859e-08, 
    6.306583e-08, 6.327619e-08, 6.308686e-08, 6.341482e-08, 6.348623e-08, 
    6.343743e-08, 6.362488e-08, 6.307636e-08, 6.328702e-08, 6.170274e-08, 
    6.171205e-08, 6.175546e-08, 6.156463e-08, 6.155295e-08, 6.137806e-08, 
    6.153368e-08, 6.159995e-08, 6.176817e-08, 6.186767e-08, 6.196226e-08, 
    6.217023e-08, 6.240249e-08, 6.272727e-08, 6.296058e-08, 6.311698e-08, 
    6.302108e-08, 6.310574e-08, 6.301109e-08, 6.296673e-08, 6.345947e-08, 
    6.31828e-08, 6.359792e-08, 6.357495e-08, 6.338708e-08, 6.357754e-08, 
    6.171859e-08, 6.166497e-08, 6.147879e-08, 6.162449e-08, 6.135902e-08, 
    6.150762e-08, 6.159307e-08, 6.192275e-08, 6.199517e-08, 6.206234e-08, 
    6.219499e-08, 6.236523e-08, 6.266387e-08, 6.29237e-08, 6.316089e-08, 
    6.314351e-08, 6.314963e-08, 6.320262e-08, 6.307136e-08, 6.322416e-08, 
    6.324981e-08, 6.318276e-08, 6.357187e-08, 6.34607e-08, 6.357446e-08, 
    6.350208e-08, 6.16824e-08, 6.177263e-08, 6.172387e-08, 6.181556e-08, 
    6.175097e-08, 6.20382e-08, 6.212431e-08, 6.252726e-08, 6.236188e-08, 
    6.262507e-08, 6.238862e-08, 6.243052e-08, 6.263367e-08, 6.240139e-08, 
    6.290938e-08, 6.256499e-08, 6.320468e-08, 6.286079e-08, 6.322623e-08, 
    6.315987e-08, 6.326974e-08, 6.336815e-08, 6.349195e-08, 6.372039e-08, 
    6.366749e-08, 6.385851e-08, 6.190715e-08, 6.202419e-08, 6.201388e-08, 
    6.213636e-08, 6.222695e-08, 6.242326e-08, 6.273814e-08, 6.261973e-08, 
    6.28371e-08, 6.288074e-08, 6.25505e-08, 6.275327e-08, 6.210252e-08, 
    6.220766e-08, 6.214506e-08, 6.191639e-08, 6.264703e-08, 6.227206e-08, 
    6.296444e-08, 6.276132e-08, 6.335412e-08, 6.305931e-08, 6.363837e-08, 
    6.388592e-08, 6.411888e-08, 6.439114e-08, 6.208806e-08, 6.200854e-08, 
    6.215092e-08, 6.234794e-08, 6.253071e-08, 6.277371e-08, 6.279857e-08, 
    6.284409e-08, 6.2962e-08, 6.306114e-08, 6.285849e-08, 6.3086e-08, 
    6.223206e-08, 6.267957e-08, 6.197848e-08, 6.21896e-08, 6.233632e-08, 
    6.227195e-08, 6.26062e-08, 6.268498e-08, 6.30051e-08, 6.283961e-08, 
    6.382483e-08, 6.338895e-08, 6.459844e-08, 6.426044e-08, 6.198075e-08, 
    6.208779e-08, 6.24603e-08, 6.228306e-08, 6.278993e-08, 6.291469e-08, 
    6.301611e-08, 6.314576e-08, 6.315975e-08, 6.323658e-08, 6.31107e-08, 
    6.32316e-08, 6.277423e-08, 6.297861e-08, 6.241772e-08, 6.255424e-08, 
    6.249143e-08, 6.242254e-08, 6.263516e-08, 6.286168e-08, 6.286651e-08, 
    6.293915e-08, 6.314385e-08, 6.279198e-08, 6.38811e-08, 6.32085e-08, 
    6.22045e-08, 6.241068e-08, 6.244011e-08, 6.236025e-08, 6.290218e-08, 
    6.270582e-08, 6.32347e-08, 6.309176e-08, 6.332596e-08, 6.320958e-08, 
    6.319247e-08, 6.304299e-08, 6.294994e-08, 6.271483e-08, 6.252353e-08, 
    6.237183e-08, 6.24071e-08, 6.257374e-08, 6.287554e-08, 6.316102e-08, 
    6.309849e-08, 6.330816e-08, 6.275317e-08, 6.29859e-08, 6.289595e-08, 
    6.313048e-08, 6.261659e-08, 6.305422e-08, 6.250472e-08, 6.25529e-08, 
    6.270192e-08, 6.300169e-08, 6.306799e-08, 6.313881e-08, 6.309511e-08, 
    6.28832e-08, 6.284847e-08, 6.26983e-08, 6.265685e-08, 6.254241e-08, 
    6.244768e-08, 6.253423e-08, 6.262513e-08, 6.288328e-08, 6.311592e-08, 
    6.336955e-08, 6.343162e-08, 6.372798e-08, 6.348674e-08, 6.388485e-08, 
    6.35464e-08, 6.413226e-08, 6.307957e-08, 6.353643e-08, 6.27087e-08, 
    6.279787e-08, 6.295917e-08, 6.332909e-08, 6.312938e-08, 6.336294e-08, 
    6.284711e-08, 6.25795e-08, 6.251025e-08, 6.238105e-08, 6.251319e-08, 
    6.250245e-08, 6.262889e-08, 6.258826e-08, 6.289185e-08, 6.272878e-08, 
    6.319203e-08, 6.336109e-08, 6.38385e-08, 6.413116e-08, 6.442907e-08, 
    6.456059e-08, 6.460062e-08, 6.461735e-08 ;

 SOIL1_HR_S3 =
  7.286273e-10, 7.318323e-10, 7.312092e-10, 7.337944e-10, 7.323603e-10, 
    7.34053e-10, 7.29277e-10, 7.319596e-10, 7.302471e-10, 7.289158e-10, 
    7.388112e-10, 7.339097e-10, 7.439023e-10, 7.407763e-10, 7.486288e-10, 
    7.434159e-10, 7.496798e-10, 7.484783e-10, 7.520945e-10, 7.510585e-10, 
    7.556841e-10, 7.525727e-10, 7.580818e-10, 7.54941e-10, 7.554324e-10, 
    7.5247e-10, 7.34896e-10, 7.38201e-10, 7.347002e-10, 7.351715e-10, 
    7.3496e-10, 7.323899e-10, 7.310949e-10, 7.283823e-10, 7.288747e-10, 
    7.30867e-10, 7.353834e-10, 7.338502e-10, 7.37714e-10, 7.376267e-10, 
    7.419283e-10, 7.399888e-10, 7.472187e-10, 7.451638e-10, 7.511017e-10, 
    7.496084e-10, 7.510316e-10, 7.506001e-10, 7.510372e-10, 7.488471e-10, 
    7.497855e-10, 7.478583e-10, 7.403521e-10, 7.425581e-10, 7.359786e-10, 
    7.320226e-10, 7.293947e-10, 7.2753e-10, 7.277937e-10, 7.282962e-10, 
    7.308787e-10, 7.333066e-10, 7.351569e-10, 7.363947e-10, 7.376142e-10, 
    7.413059e-10, 7.432596e-10, 7.476342e-10, 7.468446e-10, 7.481822e-10, 
    7.494599e-10, 7.516051e-10, 7.512519e-10, 7.521971e-10, 7.481468e-10, 
    7.508387e-10, 7.463949e-10, 7.476104e-10, 7.379461e-10, 7.342638e-10, 
    7.32699e-10, 7.31329e-10, 7.279963e-10, 7.302978e-10, 7.293905e-10, 
    7.315489e-10, 7.329204e-10, 7.322421e-10, 7.364285e-10, 7.348009e-10, 
    7.433754e-10, 7.396821e-10, 7.493108e-10, 7.470067e-10, 7.498631e-10, 
    7.484055e-10, 7.50903e-10, 7.486553e-10, 7.525489e-10, 7.533967e-10, 
    7.528173e-10, 7.550429e-10, 7.485307e-10, 7.510316e-10, 7.322231e-10, 
    7.323337e-10, 7.328491e-10, 7.305836e-10, 7.30445e-10, 7.283688e-10, 
    7.302162e-10, 7.310029e-10, 7.329999e-10, 7.341812e-10, 7.353041e-10, 
    7.377731e-10, 7.405305e-10, 7.443861e-10, 7.471561e-10, 7.490129e-10, 
    7.478743e-10, 7.488795e-10, 7.477558e-10, 7.472291e-10, 7.53079e-10, 
    7.497942e-10, 7.547228e-10, 7.544501e-10, 7.522196e-10, 7.544808e-10, 
    7.324114e-10, 7.317748e-10, 7.295645e-10, 7.312942e-10, 7.281427e-10, 
    7.299068e-10, 7.309212e-10, 7.34835e-10, 7.356948e-10, 7.364923e-10, 
    7.380671e-10, 7.400881e-10, 7.436335e-10, 7.467182e-10, 7.495342e-10, 
    7.493278e-10, 7.494005e-10, 7.500296e-10, 7.484713e-10, 7.502854e-10, 
    7.505899e-10, 7.497938e-10, 7.544135e-10, 7.530937e-10, 7.544442e-10, 
    7.535849e-10, 7.319817e-10, 7.33053e-10, 7.324741e-10, 7.335626e-10, 
    7.327958e-10, 7.362057e-10, 7.372279e-10, 7.420116e-10, 7.400483e-10, 
    7.431729e-10, 7.403657e-10, 7.408631e-10, 7.432749e-10, 7.405174e-10, 
    7.465482e-10, 7.424596e-10, 7.500541e-10, 7.459713e-10, 7.503099e-10, 
    7.49522e-10, 7.508265e-10, 7.519949e-10, 7.534646e-10, 7.561767e-10, 
    7.555487e-10, 7.578167e-10, 7.346499e-10, 7.360393e-10, 7.359169e-10, 
    7.37371e-10, 7.384464e-10, 7.407771e-10, 7.445152e-10, 7.431095e-10, 
    7.456901e-10, 7.462082e-10, 7.422876e-10, 7.446949e-10, 7.369692e-10, 
    7.382175e-10, 7.374742e-10, 7.347595e-10, 7.434335e-10, 7.38982e-10, 
    7.472019e-10, 7.447904e-10, 7.518283e-10, 7.483282e-10, 7.55203e-10, 
    7.58142e-10, 7.609078e-10, 7.641405e-10, 7.367976e-10, 7.358535e-10, 
    7.375439e-10, 7.398828e-10, 7.420526e-10, 7.449375e-10, 7.452326e-10, 
    7.457731e-10, 7.471729e-10, 7.4835e-10, 7.45944e-10, 7.48645e-10, 
    7.385071e-10, 7.438198e-10, 7.354966e-10, 7.38003e-10, 7.397448e-10, 
    7.389807e-10, 7.429488e-10, 7.438841e-10, 7.476846e-10, 7.457199e-10, 
    7.574167e-10, 7.522417e-10, 7.666016e-10, 7.625887e-10, 7.355236e-10, 
    7.367943e-10, 7.412168e-10, 7.391125e-10, 7.451301e-10, 7.466112e-10, 
    7.478153e-10, 7.493546e-10, 7.495207e-10, 7.504327e-10, 7.489382e-10, 
    7.503737e-10, 7.449437e-10, 7.473702e-10, 7.407112e-10, 7.42332e-10, 
    7.415863e-10, 7.407685e-10, 7.432926e-10, 7.459819e-10, 7.460393e-10, 
    7.469016e-10, 7.493319e-10, 7.451544e-10, 7.580848e-10, 7.500995e-10, 
    7.381799e-10, 7.406276e-10, 7.409771e-10, 7.400289e-10, 7.464627e-10, 
    7.441316e-10, 7.504105e-10, 7.487135e-10, 7.51494e-10, 7.501123e-10, 
    7.49909e-10, 7.481344e-10, 7.470297e-10, 7.442384e-10, 7.419674e-10, 
    7.401664e-10, 7.405851e-10, 7.425635e-10, 7.461464e-10, 7.495358e-10, 
    7.487934e-10, 7.512826e-10, 7.446938e-10, 7.474567e-10, 7.463888e-10, 
    7.491731e-10, 7.430722e-10, 7.482678e-10, 7.417441e-10, 7.423161e-10, 
    7.440853e-10, 7.476441e-10, 7.484313e-10, 7.49272e-10, 7.487532e-10, 
    7.462373e-10, 7.458251e-10, 7.440423e-10, 7.435501e-10, 7.421915e-10, 
    7.410669e-10, 7.420945e-10, 7.431736e-10, 7.462383e-10, 7.490003e-10, 
    7.520115e-10, 7.527484e-10, 7.562669e-10, 7.534028e-10, 7.581293e-10, 
    7.541111e-10, 7.610668e-10, 7.485687e-10, 7.539928e-10, 7.441657e-10, 
    7.452244e-10, 7.471393e-10, 7.515311e-10, 7.4916e-10, 7.51933e-10, 
    7.45809e-10, 7.426318e-10, 7.418097e-10, 7.40276e-10, 7.418447e-10, 
    7.417171e-10, 7.432183e-10, 7.427359e-10, 7.463401e-10, 7.444041e-10, 
    7.49904e-10, 7.51911e-10, 7.575791e-10, 7.610538e-10, 7.645907e-10, 
    7.661523e-10, 7.666275e-10, 7.668262e-10 ;

 SOIL2C =
  5.784044, 5.784051, 5.78405, 5.784055, 5.784052, 5.784055, 5.784046, 
    5.784051, 5.784048, 5.784045, 5.784065, 5.784055, 5.784075, 5.784069, 
    5.784084, 5.784074, 5.784086, 5.784084, 5.784091, 5.784089, 5.784098, 
    5.784092, 5.784102, 5.784096, 5.784097, 5.784091, 5.784057, 5.784063, 
    5.784057, 5.784058, 5.784057, 5.784052, 5.78405, 5.784044, 5.784045, 
    5.784049, 5.784058, 5.784055, 5.784062, 5.784062, 5.784071, 5.784067, 
    5.784081, 5.784077, 5.784089, 5.784086, 5.784089, 5.784088, 5.784089, 
    5.784084, 5.784086, 5.784082, 5.784068, 5.784072, 5.784059, 5.784051, 
    5.784046, 5.784042, 5.784043, 5.784044, 5.784049, 5.784054, 5.784058, 
    5.78406, 5.784062, 5.78407, 5.784073, 5.784082, 5.784081, 5.784083, 
    5.784086, 5.78409, 5.784089, 5.784091, 5.784083, 5.784088, 5.78408, 
    5.784082, 5.784063, 5.784056, 5.784052, 5.78405, 5.784043, 5.784048, 
    5.784046, 5.78405, 5.784053, 5.784051, 5.78406, 5.784057, 5.784074, 
    5.784066, 5.784085, 5.784081, 5.784086, 5.784083, 5.784089, 5.784084, 
    5.784092, 5.784093, 5.784092, 5.784097, 5.784084, 5.784089, 5.784051, 
    5.784052, 5.784053, 5.784049, 5.784048, 5.784044, 5.784048, 5.784049, 
    5.784053, 5.784055, 5.784058, 5.784062, 5.784068, 5.784076, 5.784081, 
    5.784085, 5.784082, 5.784084, 5.784082, 5.784081, 5.784093, 5.784086, 
    5.784096, 5.784095, 5.784091, 5.784096, 5.784052, 5.78405, 5.784046, 
    5.78405, 5.784043, 5.784047, 5.784049, 5.784057, 5.784059, 5.78406, 
    5.784063, 5.784067, 5.784074, 5.78408, 5.784086, 5.784085, 5.784085, 
    5.784087, 5.784084, 5.784087, 5.784088, 5.784086, 5.784095, 5.784093, 
    5.784095, 5.784094, 5.784051, 5.784053, 5.784052, 5.784054, 5.784053, 
    5.78406, 5.784061, 5.784071, 5.784067, 5.784073, 5.784068, 5.784069, 
    5.784073, 5.784068, 5.78408, 5.784072, 5.784087, 5.784079, 5.784087, 
    5.784086, 5.784088, 5.784091, 5.784093, 5.784099, 5.784098, 5.784102, 
    5.784056, 5.784059, 5.784059, 5.784062, 5.784064, 5.784069, 5.784076, 
    5.784073, 5.784078, 5.784079, 5.784071, 5.784076, 5.784061, 5.784063, 
    5.784062, 5.784057, 5.784074, 5.784065, 5.784081, 5.784076, 5.784091, 
    5.784083, 5.784097, 5.784103, 5.784108, 5.784114, 5.78406, 5.784059, 
    5.784062, 5.784067, 5.784071, 5.784077, 5.784077, 5.784078, 5.784081, 
    5.784083, 5.784079, 5.784084, 5.784064, 5.784074, 5.784058, 5.784063, 
    5.784067, 5.784065, 5.784073, 5.784075, 5.784082, 5.784078, 5.784101, 
    5.784091, 5.78412, 5.784111, 5.784058, 5.78406, 5.78407, 5.784065, 
    5.784077, 5.78408, 5.784082, 5.784085, 5.784086, 5.784088, 5.784085, 
    5.784088, 5.784077, 5.784081, 5.784069, 5.784071, 5.78407, 5.784069, 
    5.784073, 5.784079, 5.784079, 5.784081, 5.784085, 5.784077, 5.784102, 
    5.784087, 5.784063, 5.784068, 5.784069, 5.784067, 5.78408, 5.784075, 
    5.784088, 5.784084, 5.78409, 5.784087, 5.784087, 5.784083, 5.784081, 
    5.784075, 5.784071, 5.784067, 5.784068, 5.784072, 5.784079, 5.784086, 
    5.784084, 5.784089, 5.784076, 5.784081, 5.78408, 5.784085, 5.784073, 
    5.784083, 5.78407, 5.784071, 5.784075, 5.784082, 5.784083, 5.784085, 
    5.784084, 5.784079, 5.784079, 5.784075, 5.784074, 5.784071, 5.784069, 
    5.784071, 5.784073, 5.784079, 5.784085, 5.784091, 5.784092, 5.784099, 
    5.784093, 5.784103, 5.784095, 5.784109, 5.784084, 5.784095, 5.784075, 
    5.784077, 5.784081, 5.78409, 5.784085, 5.784091, 5.784079, 5.784072, 
    5.78407, 5.784068, 5.78407, 5.78407, 5.784073, 5.784072, 5.78408, 
    5.784076, 5.784087, 5.784091, 5.784101, 5.784109, 5.784115, 5.784119, 
    5.78412, 5.78412 ;

 SOIL2C_TO_SOIL1C =
  1.086284e-09, 1.091064e-09, 1.090134e-09, 1.09399e-09, 1.091851e-09, 
    1.094376e-09, 1.087253e-09, 1.091253e-09, 1.088699e-09, 1.086714e-09, 
    1.101472e-09, 1.094162e-09, 1.109065e-09, 1.104403e-09, 1.116113e-09, 
    1.108339e-09, 1.117681e-09, 1.115889e-09, 1.121282e-09, 1.119737e-09, 
    1.126635e-09, 1.121995e-09, 1.130211e-09, 1.125527e-09, 1.12626e-09, 
    1.121842e-09, 1.095633e-09, 1.100562e-09, 1.095341e-09, 1.096044e-09, 
    1.095728e-09, 1.091895e-09, 1.089964e-09, 1.085918e-09, 1.086653e-09, 
    1.089624e-09, 1.09636e-09, 1.094073e-09, 1.099835e-09, 1.099705e-09, 
    1.106121e-09, 1.103228e-09, 1.11401e-09, 1.110946e-09, 1.119801e-09, 
    1.117574e-09, 1.119697e-09, 1.119053e-09, 1.119705e-09, 1.116439e-09, 
    1.117838e-09, 1.114964e-09, 1.10377e-09, 1.10706e-09, 1.097247e-09, 
    1.091347e-09, 1.087428e-09, 1.084647e-09, 1.08504e-09, 1.08579e-09, 
    1.089641e-09, 1.093262e-09, 1.096022e-09, 1.097868e-09, 1.099687e-09, 
    1.105192e-09, 1.108106e-09, 1.11463e-09, 1.113453e-09, 1.115447e-09, 
    1.117353e-09, 1.120552e-09, 1.120026e-09, 1.121435e-09, 1.115395e-09, 
    1.119409e-09, 1.112782e-09, 1.114595e-09, 1.100182e-09, 1.09469e-09, 
    1.092356e-09, 1.090313e-09, 1.085343e-09, 1.088775e-09, 1.087422e-09, 
    1.090641e-09, 1.092686e-09, 1.091675e-09, 1.097918e-09, 1.095491e-09, 
    1.108279e-09, 1.102771e-09, 1.117131e-09, 1.113694e-09, 1.117954e-09, 
    1.11578e-09, 1.119505e-09, 1.116153e-09, 1.12196e-09, 1.123224e-09, 
    1.12236e-09, 1.125679e-09, 1.115967e-09, 1.119697e-09, 1.091646e-09, 
    1.091811e-09, 1.09258e-09, 1.089201e-09, 1.088995e-09, 1.085898e-09, 
    1.088653e-09, 1.089827e-09, 1.092805e-09, 1.094567e-09, 1.096241e-09, 
    1.099924e-09, 1.104036e-09, 1.109786e-09, 1.113917e-09, 1.116686e-09, 
    1.114988e-09, 1.116487e-09, 1.114811e-09, 1.114026e-09, 1.12275e-09, 
    1.117851e-09, 1.125202e-09, 1.124795e-09, 1.121469e-09, 1.124841e-09, 
    1.091927e-09, 1.090978e-09, 1.087681e-09, 1.090261e-09, 1.085561e-09, 
    1.088192e-09, 1.089705e-09, 1.095542e-09, 1.096824e-09, 1.098013e-09, 
    1.100362e-09, 1.103376e-09, 1.108664e-09, 1.113264e-09, 1.117464e-09, 
    1.117156e-09, 1.117264e-09, 1.118203e-09, 1.115879e-09, 1.118584e-09, 
    1.119038e-09, 1.117851e-09, 1.12474e-09, 1.122772e-09, 1.124786e-09, 
    1.123505e-09, 1.091286e-09, 1.092884e-09, 1.092021e-09, 1.093644e-09, 
    1.092501e-09, 1.097586e-09, 1.099111e-09, 1.106245e-09, 1.103317e-09, 
    1.107977e-09, 1.10379e-09, 1.104532e-09, 1.108129e-09, 1.104016e-09, 
    1.113011e-09, 1.106913e-09, 1.118239e-09, 1.11215e-09, 1.118621e-09, 
    1.117445e-09, 1.119391e-09, 1.121133e-09, 1.123325e-09, 1.12737e-09, 
    1.126433e-09, 1.129816e-09, 1.095266e-09, 1.097338e-09, 1.097155e-09, 
    1.099324e-09, 1.100928e-09, 1.104404e-09, 1.109979e-09, 1.107882e-09, 
    1.111731e-09, 1.112503e-09, 1.106656e-09, 1.110247e-09, 1.098725e-09, 
    1.100586e-09, 1.099478e-09, 1.095429e-09, 1.108365e-09, 1.101727e-09, 
    1.113985e-09, 1.110389e-09, 1.120885e-09, 1.115665e-09, 1.125918e-09, 
    1.130301e-09, 1.134425e-09, 1.139246e-09, 1.098469e-09, 1.097061e-09, 
    1.099582e-09, 1.10307e-09, 1.106306e-09, 1.110608e-09, 1.111049e-09, 
    1.111855e-09, 1.113942e-09, 1.115698e-09, 1.11211e-09, 1.116138e-09, 
    1.101018e-09, 1.108942e-09, 1.096529e-09, 1.100267e-09, 1.102864e-09, 
    1.101725e-09, 1.107643e-09, 1.109037e-09, 1.114705e-09, 1.111775e-09, 
    1.129219e-09, 1.121501e-09, 1.142916e-09, 1.136932e-09, 1.096569e-09, 
    1.098464e-09, 1.105059e-09, 1.101921e-09, 1.110896e-09, 1.113105e-09, 
    1.1149e-09, 1.117196e-09, 1.117444e-09, 1.118804e-09, 1.116575e-09, 
    1.118716e-09, 1.110618e-09, 1.114236e-09, 1.104305e-09, 1.106723e-09, 
    1.105611e-09, 1.104391e-09, 1.108155e-09, 1.112166e-09, 1.112252e-09, 
    1.113538e-09, 1.117162e-09, 1.110932e-09, 1.130215e-09, 1.118307e-09, 
    1.10053e-09, 1.104181e-09, 1.104702e-09, 1.103288e-09, 1.112883e-09, 
    1.109406e-09, 1.118771e-09, 1.11624e-09, 1.120386e-09, 1.118326e-09, 
    1.118023e-09, 1.115376e-09, 1.113729e-09, 1.109566e-09, 1.106179e-09, 
    1.103493e-09, 1.104118e-09, 1.107068e-09, 1.112411e-09, 1.117466e-09, 
    1.116359e-09, 1.120071e-09, 1.110245e-09, 1.114365e-09, 1.112773e-09, 
    1.116925e-09, 1.107826e-09, 1.115575e-09, 1.105846e-09, 1.106699e-09, 
    1.109338e-09, 1.114645e-09, 1.115819e-09, 1.117073e-09, 1.116299e-09, 
    1.112547e-09, 1.111932e-09, 1.109273e-09, 1.108539e-09, 1.106513e-09, 
    1.104836e-09, 1.106368e-09, 1.107978e-09, 1.112548e-09, 1.116667e-09, 
    1.121158e-09, 1.122257e-09, 1.127504e-09, 1.123233e-09, 1.130282e-09, 
    1.124289e-09, 1.134662e-09, 1.116024e-09, 1.124113e-09, 1.109458e-09, 
    1.111036e-09, 1.113892e-09, 1.120442e-09, 1.116906e-09, 1.121041e-09, 
    1.111908e-09, 1.10717e-09, 1.105944e-09, 1.103656e-09, 1.105996e-09, 
    1.105806e-09, 1.108044e-09, 1.107325e-09, 1.1127e-09, 1.109813e-09, 
    1.118015e-09, 1.121008e-09, 1.129461e-09, 1.134643e-09, 1.139917e-09, 
    1.142246e-09, 1.142955e-09, 1.143251e-09 ;

 SOIL2C_TO_SOIL3C =
  7.759168e-11, 7.793311e-11, 7.786673e-11, 7.814212e-11, 7.798936e-11, 
    7.816969e-11, 7.766091e-11, 7.794667e-11, 7.776424e-11, 7.762242e-11, 
    7.867657e-11, 7.815441e-11, 7.92189e-11, 7.88859e-11, 7.972238e-11, 
    7.916708e-11, 7.983435e-11, 7.970635e-11, 8.009157e-11, 7.998121e-11, 
    8.047395e-11, 8.01425e-11, 8.072935e-11, 8.039479e-11, 8.044713e-11, 
    8.013157e-11, 7.825948e-11, 7.861155e-11, 7.823862e-11, 7.828883e-11, 
    7.82663e-11, 7.799252e-11, 7.785456e-11, 7.756559e-11, 7.761804e-11, 
    7.783028e-11, 7.831141e-11, 7.814808e-11, 7.855968e-11, 7.855038e-11, 
    7.900861e-11, 7.880201e-11, 7.957218e-11, 7.935328e-11, 7.998582e-11, 
    7.982674e-11, 7.997834e-11, 7.993237e-11, 7.997895e-11, 7.974565e-11, 
    7.98456e-11, 7.964031e-11, 7.88407e-11, 7.907571e-11, 7.837481e-11, 
    7.795338e-11, 7.767344e-11, 7.747479e-11, 7.750288e-11, 7.755641e-11, 
    7.783152e-11, 7.809017e-11, 7.828728e-11, 7.841913e-11, 7.854905e-11, 
    7.894231e-11, 7.915043e-11, 7.961645e-11, 7.953233e-11, 7.967482e-11, 
    7.981091e-11, 8.003943e-11, 8.000182e-11, 8.01025e-11, 7.967105e-11, 
    7.99578e-11, 7.948443e-11, 7.96139e-11, 7.85844e-11, 7.819214e-11, 
    7.802544e-11, 7.787949e-11, 7.752447e-11, 7.776964e-11, 7.7673e-11, 
    7.790293e-11, 7.804903e-11, 7.797677e-11, 7.842274e-11, 7.824936e-11, 
    7.916277e-11, 7.876933e-11, 7.979505e-11, 7.95496e-11, 7.985387e-11, 
    7.96986e-11, 7.996465e-11, 7.972521e-11, 8.013997e-11, 8.023029e-11, 
    8.016857e-11, 8.040564e-11, 7.971194e-11, 7.997835e-11, 7.797474e-11, 
    7.798653e-11, 7.804143e-11, 7.780009e-11, 7.778533e-11, 7.756415e-11, 
    7.776095e-11, 7.784476e-11, 7.80575e-11, 7.818333e-11, 7.830296e-11, 
    7.856597e-11, 7.885971e-11, 7.927044e-11, 7.956551e-11, 7.97633e-11, 
    7.964202e-11, 7.97491e-11, 7.962939e-11, 7.957329e-11, 8.019645e-11, 
    7.984654e-11, 8.037154e-11, 8.034249e-11, 8.010489e-11, 8.034576e-11, 
    7.799481e-11, 7.792698e-11, 7.769153e-11, 7.78758e-11, 7.754006e-11, 
    7.772799e-11, 7.783606e-11, 7.825299e-11, 7.834459e-11, 7.842953e-11, 
    7.859729e-11, 7.881259e-11, 7.919027e-11, 7.951886e-11, 7.981883e-11, 
    7.979686e-11, 7.980459e-11, 7.987161e-11, 7.970561e-11, 7.989886e-11, 
    7.99313e-11, 7.984649e-11, 8.03386e-11, 8.019801e-11, 8.034187e-11, 
    8.025033e-11, 7.794903e-11, 7.806315e-11, 7.800148e-11, 7.811744e-11, 
    7.803575e-11, 7.8399e-11, 7.85079e-11, 7.901749e-11, 7.880835e-11, 
    7.914119e-11, 7.884216e-11, 7.889515e-11, 7.915207e-11, 7.885832e-11, 
    7.950075e-11, 7.906521e-11, 7.987421e-11, 7.94393e-11, 7.990147e-11, 
    7.981753e-11, 7.995649e-11, 8.008095e-11, 8.023752e-11, 8.052642e-11, 
    8.045951e-11, 8.070111e-11, 7.823327e-11, 7.838128e-11, 7.836824e-11, 
    7.852314e-11, 7.863769e-11, 7.888597e-11, 7.928419e-11, 7.913444e-11, 
    7.940935e-11, 7.946453e-11, 7.904689e-11, 7.930332e-11, 7.848034e-11, 
    7.861331e-11, 7.853414e-11, 7.824495e-11, 7.916896e-11, 7.869476e-11, 
    7.957039e-11, 7.93135e-11, 8.006321e-11, 7.969037e-11, 8.042269e-11, 
    8.073577e-11, 8.103038e-11, 8.137472e-11, 7.846206e-11, 7.836148e-11, 
    7.854156e-11, 7.879071e-11, 7.902186e-11, 7.932918e-11, 7.936062e-11, 
    7.941819e-11, 7.95673e-11, 7.969269e-11, 7.943639e-11, 7.972412e-11, 
    7.864417e-11, 7.921012e-11, 7.832347e-11, 7.859047e-11, 7.877602e-11, 
    7.869462e-11, 7.911732e-11, 7.921695e-11, 7.962181e-11, 7.941252e-11, 
    8.06585e-11, 8.010725e-11, 8.163688e-11, 8.120942e-11, 7.832635e-11, 
    7.846171e-11, 7.893282e-11, 7.870866e-11, 7.934969e-11, 7.950747e-11, 
    7.963573e-11, 7.97997e-11, 7.98174e-11, 7.991455e-11, 7.975536e-11, 
    7.990826e-11, 7.932983e-11, 7.958832e-11, 7.887896e-11, 7.905162e-11, 
    7.897219e-11, 7.888507e-11, 7.915395e-11, 7.944043e-11, 7.944654e-11, 
    7.95384e-11, 7.979728e-11, 7.935228e-11, 8.072967e-11, 7.987905e-11, 
    7.860931e-11, 7.887006e-11, 7.890728e-11, 7.880628e-11, 7.949165e-11, 
    7.924332e-11, 7.991218e-11, 7.973141e-11, 8.00276e-11, 7.988041e-11, 
    7.985877e-11, 7.966973e-11, 7.955204e-11, 7.925471e-11, 7.901278e-11, 
    7.882093e-11, 7.886554e-11, 7.907628e-11, 7.945795e-11, 7.981901e-11, 
    7.973992e-11, 8.000509e-11, 7.93032e-11, 7.959752e-11, 7.948377e-11, 
    7.978037e-11, 7.913047e-11, 7.968393e-11, 7.8989e-11, 7.904993e-11, 
    7.923839e-11, 7.961749e-11, 7.970135e-11, 7.979091e-11, 7.973564e-11, 
    7.946764e-11, 7.942373e-11, 7.923381e-11, 7.918138e-11, 7.903666e-11, 
    7.891685e-11, 7.902632e-11, 7.914128e-11, 7.946774e-11, 7.976196e-11, 
    8.008273e-11, 8.016122e-11, 8.053603e-11, 8.023093e-11, 8.073441e-11, 
    8.030639e-11, 8.104731e-11, 7.971599e-11, 8.029377e-11, 7.924696e-11, 
    7.935973e-11, 7.956372e-11, 8.003156e-11, 7.977898e-11, 8.007436e-11, 
    7.942201e-11, 7.908356e-11, 7.899598e-11, 7.883259e-11, 7.899971e-11, 
    7.898612e-11, 7.914603e-11, 7.909464e-11, 7.947858e-11, 7.927235e-11, 
    7.985822e-11, 8.007203e-11, 8.067579e-11, 8.104593e-11, 8.142268e-11, 
    8.158901e-11, 8.163964e-11, 8.16608e-11 ;

 SOIL2C_vr =
  20.00644, 20.00646, 20.00646, 20.00647, 20.00646, 20.00647, 20.00644, 
    20.00646, 20.00645, 20.00644, 20.0065, 20.00647, 20.00652, 20.00651, 
    20.00655, 20.00652, 20.00655, 20.00655, 20.00657, 20.00656, 20.00658, 
    20.00657, 20.0066, 20.00658, 20.00658, 20.00657, 20.00648, 20.00649, 
    20.00647, 20.00648, 20.00648, 20.00646, 20.00645, 20.00644, 20.00644, 
    20.00645, 20.00648, 20.00647, 20.00649, 20.00649, 20.00651, 20.0065, 
    20.00654, 20.00653, 20.00656, 20.00655, 20.00656, 20.00656, 20.00656, 
    20.00655, 20.00655, 20.00654, 20.0065, 20.00652, 20.00648, 20.00646, 
    20.00645, 20.00644, 20.00644, 20.00644, 20.00645, 20.00647, 20.00648, 
    20.00648, 20.00649, 20.00651, 20.00652, 20.00654, 20.00654, 20.00654, 
    20.00655, 20.00656, 20.00656, 20.00657, 20.00654, 20.00656, 20.00654, 
    20.00654, 20.00649, 20.00647, 20.00646, 20.00646, 20.00644, 20.00645, 
    20.00645, 20.00646, 20.00647, 20.00646, 20.00648, 20.00648, 20.00652, 
    20.0065, 20.00655, 20.00654, 20.00655, 20.00655, 20.00656, 20.00655, 
    20.00657, 20.00657, 20.00657, 20.00658, 20.00655, 20.00656, 20.00646, 
    20.00646, 20.00646, 20.00645, 20.00645, 20.00644, 20.00645, 20.00645, 
    20.00647, 20.00647, 20.00648, 20.00649, 20.0065, 20.00653, 20.00654, 
    20.00655, 20.00654, 20.00655, 20.00654, 20.00654, 20.00657, 20.00655, 
    20.00658, 20.00658, 20.00657, 20.00658, 20.00646, 20.00646, 20.00645, 
    20.00646, 20.00644, 20.00645, 20.00645, 20.00648, 20.00648, 20.00648, 
    20.00649, 20.0065, 20.00652, 20.00654, 20.00655, 20.00655, 20.00655, 
    20.00655, 20.00655, 20.00656, 20.00656, 20.00655, 20.00658, 20.00657, 
    20.00658, 20.00657, 20.00646, 20.00647, 20.00646, 20.00647, 20.00646, 
    20.00648, 20.00649, 20.00651, 20.0065, 20.00652, 20.0065, 20.00651, 
    20.00652, 20.0065, 20.00654, 20.00652, 20.00656, 20.00653, 20.00656, 
    20.00655, 20.00656, 20.00657, 20.00657, 20.00659, 20.00658, 20.0066, 
    20.00647, 20.00648, 20.00648, 20.00649, 20.00649, 20.00651, 20.00653, 
    20.00652, 20.00653, 20.00653, 20.00651, 20.00653, 20.00649, 20.00649, 
    20.00649, 20.00648, 20.00652, 20.0065, 20.00654, 20.00653, 20.00656, 
    20.00655, 20.00658, 20.0066, 20.00661, 20.00663, 20.00648, 20.00648, 
    20.00649, 20.0065, 20.00651, 20.00653, 20.00653, 20.00653, 20.00654, 
    20.00655, 20.00653, 20.00655, 20.00649, 20.00652, 20.00648, 20.00649, 
    20.0065, 20.0065, 20.00652, 20.00652, 20.00654, 20.00653, 20.00659, 
    20.00657, 20.00664, 20.00662, 20.00648, 20.00648, 20.00651, 20.0065, 
    20.00653, 20.00654, 20.00654, 20.00655, 20.00655, 20.00656, 20.00655, 
    20.00656, 20.00653, 20.00654, 20.00651, 20.00651, 20.00651, 20.00651, 
    20.00652, 20.00653, 20.00653, 20.00654, 20.00655, 20.00653, 20.0066, 
    20.00656, 20.00649, 20.00651, 20.00651, 20.0065, 20.00654, 20.00652, 
    20.00656, 20.00655, 20.00656, 20.00656, 20.00655, 20.00654, 20.00654, 
    20.00653, 20.00651, 20.0065, 20.00651, 20.00652, 20.00653, 20.00655, 
    20.00655, 20.00656, 20.00653, 20.00654, 20.00654, 20.00655, 20.00652, 
    20.00655, 20.00651, 20.00651, 20.00652, 20.00654, 20.00655, 20.00655, 
    20.00655, 20.00653, 20.00653, 20.00652, 20.00652, 20.00651, 20.00651, 
    20.00651, 20.00652, 20.00653, 20.00655, 20.00657, 20.00657, 20.00659, 
    20.00657, 20.0066, 20.00658, 20.00661, 20.00655, 20.00657, 20.00652, 
    20.00653, 20.00654, 20.00656, 20.00655, 20.00657, 20.00653, 20.00652, 
    20.00651, 20.0065, 20.00651, 20.00651, 20.00652, 20.00652, 20.00653, 
    20.00653, 20.00655, 20.00657, 20.00659, 20.00661, 20.00663, 20.00664, 
    20.00664, 20.00664,
  20.00607, 20.00609, 20.00609, 20.00611, 20.0061, 20.00611, 20.00608, 
    20.0061, 20.00608, 20.00607, 20.00614, 20.00611, 20.00618, 20.00616, 
    20.00621, 20.00618, 20.00622, 20.00621, 20.00624, 20.00623, 20.00626, 
    20.00624, 20.00628, 20.00626, 20.00626, 20.00624, 20.00612, 20.00614, 
    20.00611, 20.00612, 20.00612, 20.0061, 20.00609, 20.00607, 20.00607, 
    20.00609, 20.00612, 20.00611, 20.00614, 20.00614, 20.00617, 20.00615, 
    20.0062, 20.00619, 20.00623, 20.00622, 20.00623, 20.00623, 20.00623, 
    20.00621, 20.00622, 20.00621, 20.00616, 20.00617, 20.00612, 20.0061, 
    20.00608, 20.00606, 20.00607, 20.00607, 20.00609, 20.00611, 20.00612, 
    20.00613, 20.00614, 20.00616, 20.00618, 20.00621, 20.0062, 20.00621, 
    20.00622, 20.00623, 20.00623, 20.00624, 20.00621, 20.00623, 20.0062, 
    20.00621, 20.00614, 20.00611, 20.0061, 20.00609, 20.00607, 20.00608, 
    20.00608, 20.00609, 20.0061, 20.0061, 20.00613, 20.00611, 20.00618, 
    20.00615, 20.00622, 20.0062, 20.00622, 20.00621, 20.00623, 20.00621, 
    20.00624, 20.00625, 20.00624, 20.00626, 20.00621, 20.00623, 20.0061, 
    20.0061, 20.0061, 20.00609, 20.00608, 20.00607, 20.00608, 20.00609, 
    20.0061, 20.00611, 20.00612, 20.00614, 20.00616, 20.00618, 20.0062, 
    20.00622, 20.00621, 20.00621, 20.00621, 20.0062, 20.00624, 20.00622, 
    20.00626, 20.00625, 20.00624, 20.00625, 20.0061, 20.00609, 20.00608, 
    20.00609, 20.00607, 20.00608, 20.00609, 20.00611, 20.00612, 20.00613, 
    20.00614, 20.00615, 20.00618, 20.0062, 20.00622, 20.00622, 20.00622, 
    20.00622, 20.00621, 20.00622, 20.00623, 20.00622, 20.00625, 20.00624, 
    20.00625, 20.00625, 20.0061, 20.0061, 20.0061, 20.00611, 20.0061, 
    20.00612, 20.00613, 20.00617, 20.00615, 20.00617, 20.00616, 20.00616, 
    20.00618, 20.00616, 20.0062, 20.00617, 20.00622, 20.0062, 20.00623, 
    20.00622, 20.00623, 20.00624, 20.00625, 20.00627, 20.00626, 20.00628, 
    20.00611, 20.00612, 20.00612, 20.00613, 20.00614, 20.00616, 20.00618, 
    20.00617, 20.00619, 20.0062, 20.00617, 20.00619, 20.00613, 20.00614, 
    20.00613, 20.00611, 20.00618, 20.00615, 20.0062, 20.00619, 20.00624, 
    20.00621, 20.00626, 20.00628, 20.0063, 20.00632, 20.00613, 20.00612, 
    20.00613, 20.00615, 20.00617, 20.00619, 20.00619, 20.00619, 20.0062, 
    20.00621, 20.00619, 20.00621, 20.00614, 20.00618, 20.00612, 20.00614, 
    20.00615, 20.00615, 20.00617, 20.00618, 20.00621, 20.00619, 20.00628, 
    20.00624, 20.00634, 20.00631, 20.00612, 20.00613, 20.00616, 20.00615, 
    20.00619, 20.0062, 20.00621, 20.00622, 20.00622, 20.00623, 20.00621, 
    20.00623, 20.00619, 20.0062, 20.00616, 20.00617, 20.00616, 20.00616, 
    20.00618, 20.0062, 20.0062, 20.0062, 20.00622, 20.00619, 20.00628, 
    20.00622, 20.00614, 20.00616, 20.00616, 20.00615, 20.0062, 20.00618, 
    20.00623, 20.00621, 20.00623, 20.00622, 20.00622, 20.00621, 20.0062, 
    20.00618, 20.00617, 20.00615, 20.00616, 20.00617, 20.0062, 20.00622, 
    20.00621, 20.00623, 20.00619, 20.0062, 20.0062, 20.00622, 20.00617, 
    20.00621, 20.00616, 20.00617, 20.00618, 20.00621, 20.00621, 20.00622, 
    20.00621, 20.0062, 20.00619, 20.00618, 20.00618, 20.00617, 20.00616, 
    20.00617, 20.00617, 20.0062, 20.00622, 20.00624, 20.00624, 20.00627, 
    20.00625, 20.00628, 20.00625, 20.0063, 20.00621, 20.00625, 20.00618, 
    20.00619, 20.0062, 20.00623, 20.00622, 20.00624, 20.00619, 20.00617, 
    20.00616, 20.00615, 20.00616, 20.00616, 20.00617, 20.00617, 20.0062, 
    20.00618, 20.00622, 20.00624, 20.00628, 20.0063, 20.00632, 20.00634, 
    20.00634, 20.00634,
  20.00552, 20.00554, 20.00554, 20.00556, 20.00555, 20.00556, 20.00553, 
    20.00555, 20.00553, 20.00552, 20.0056, 20.00556, 20.00564, 20.00561, 
    20.00567, 20.00563, 20.00568, 20.00567, 20.0057, 20.00569, 20.00573, 
    20.0057, 20.00574, 20.00572, 20.00572, 20.0057, 20.00557, 20.00559, 
    20.00557, 20.00557, 20.00557, 20.00555, 20.00554, 20.00552, 20.00552, 
    20.00554, 20.00557, 20.00556, 20.00559, 20.00559, 20.00562, 20.00561, 
    20.00566, 20.00565, 20.00569, 20.00568, 20.00569, 20.00569, 20.00569, 
    20.00567, 20.00568, 20.00567, 20.00561, 20.00563, 20.00558, 20.00555, 
    20.00553, 20.00551, 20.00551, 20.00552, 20.00554, 20.00556, 20.00557, 
    20.00558, 20.00559, 20.00562, 20.00563, 20.00566, 20.00566, 20.00567, 
    20.00568, 20.00569, 20.00569, 20.0057, 20.00567, 20.00569, 20.00566, 
    20.00566, 20.00559, 20.00556, 20.00555, 20.00554, 20.00552, 20.00553, 
    20.00553, 20.00554, 20.00555, 20.00555, 20.00558, 20.00557, 20.00563, 
    20.0056, 20.00568, 20.00566, 20.00568, 20.00567, 20.00569, 20.00567, 
    20.0057, 20.00571, 20.0057, 20.00572, 20.00567, 20.00569, 20.00555, 
    20.00555, 20.00555, 20.00554, 20.00554, 20.00552, 20.00553, 20.00554, 
    20.00555, 20.00556, 20.00557, 20.00559, 20.00561, 20.00564, 20.00566, 
    20.00567, 20.00567, 20.00567, 20.00566, 20.00566, 20.0057, 20.00568, 
    20.00572, 20.00572, 20.0057, 20.00572, 20.00555, 20.00554, 20.00553, 
    20.00554, 20.00552, 20.00553, 20.00554, 20.00557, 20.00558, 20.00558, 
    20.00559, 20.00561, 20.00563, 20.00566, 20.00568, 20.00568, 20.00568, 
    20.00568, 20.00567, 20.00568, 20.00569, 20.00568, 20.00572, 20.0057, 
    20.00572, 20.00571, 20.00555, 20.00555, 20.00555, 20.00556, 20.00555, 
    20.00558, 20.00559, 20.00562, 20.00561, 20.00563, 20.00561, 20.00561, 
    20.00563, 20.00561, 20.00566, 20.00562, 20.00568, 20.00565, 20.00568, 
    20.00568, 20.00569, 20.0057, 20.00571, 20.00573, 20.00572, 20.00574, 
    20.00557, 20.00558, 20.00558, 20.00559, 20.0056, 20.00561, 20.00564, 
    20.00563, 20.00565, 20.00565, 20.00562, 20.00564, 20.00558, 20.00559, 
    20.00559, 20.00557, 20.00563, 20.0056, 20.00566, 20.00564, 20.0057, 
    20.00567, 20.00572, 20.00574, 20.00576, 20.00579, 20.00558, 20.00558, 
    20.00559, 20.00561, 20.00562, 20.00564, 20.00565, 20.00565, 20.00566, 
    20.00567, 20.00565, 20.00567, 20.0056, 20.00564, 20.00557, 20.00559, 
    20.00561, 20.0056, 20.00563, 20.00564, 20.00566, 20.00565, 20.00574, 
    20.0057, 20.00581, 20.00578, 20.00557, 20.00558, 20.00562, 20.0056, 
    20.00565, 20.00566, 20.00567, 20.00568, 20.00568, 20.00569, 20.00567, 
    20.00569, 20.00564, 20.00566, 20.00561, 20.00562, 20.00562, 20.00561, 
    20.00563, 20.00565, 20.00565, 20.00566, 20.00568, 20.00565, 20.00574, 
    20.00568, 20.00559, 20.00561, 20.00562, 20.00561, 20.00566, 20.00564, 
    20.00569, 20.00567, 20.00569, 20.00568, 20.00568, 20.00567, 20.00566, 
    20.00564, 20.00562, 20.00561, 20.00561, 20.00563, 20.00565, 20.00568, 
    20.00567, 20.00569, 20.00564, 20.00566, 20.00566, 20.00568, 20.00563, 
    20.00567, 20.00562, 20.00562, 20.00564, 20.00566, 20.00567, 20.00568, 
    20.00567, 20.00565, 20.00565, 20.00564, 20.00563, 20.00562, 20.00562, 
    20.00562, 20.00563, 20.00565, 20.00567, 20.0057, 20.0057, 20.00573, 
    20.00571, 20.00574, 20.00571, 20.00577, 20.00567, 20.00571, 20.00564, 
    20.00565, 20.00566, 20.00569, 20.00568, 20.0057, 20.00565, 20.00563, 
    20.00562, 20.00561, 20.00562, 20.00562, 20.00563, 20.00563, 20.00566, 
    20.00564, 20.00568, 20.0057, 20.00574, 20.00577, 20.00579, 20.0058, 
    20.00581, 20.00581,
  20.00508, 20.00511, 20.0051, 20.00512, 20.00511, 20.00512, 20.00509, 
    20.00511, 20.00509, 20.00508, 20.00516, 20.00512, 20.0052, 20.00517, 
    20.00523, 20.00519, 20.00524, 20.00523, 20.00526, 20.00525, 20.00528, 
    20.00526, 20.0053, 20.00528, 20.00528, 20.00526, 20.00513, 20.00515, 
    20.00513, 20.00513, 20.00513, 20.00511, 20.0051, 20.00508, 20.00508, 
    20.0051, 20.00513, 20.00512, 20.00515, 20.00515, 20.00518, 20.00517, 
    20.00522, 20.00521, 20.00525, 20.00524, 20.00525, 20.00525, 20.00525, 
    20.00523, 20.00524, 20.00522, 20.00517, 20.00519, 20.00514, 20.00511, 
    20.00509, 20.00507, 20.00508, 20.00508, 20.0051, 20.00512, 20.00513, 
    20.00514, 20.00515, 20.00518, 20.00519, 20.00522, 20.00522, 20.00523, 
    20.00524, 20.00525, 20.00525, 20.00526, 20.00523, 20.00525, 20.00521, 
    20.00522, 20.00515, 20.00512, 20.00511, 20.0051, 20.00508, 20.00509, 
    20.00509, 20.0051, 20.00511, 20.00511, 20.00514, 20.00513, 20.00519, 
    20.00516, 20.00524, 20.00522, 20.00524, 20.00523, 20.00525, 20.00523, 
    20.00526, 20.00527, 20.00526, 20.00528, 20.00523, 20.00525, 20.00511, 
    20.00511, 20.00511, 20.0051, 20.00509, 20.00508, 20.00509, 20.0051, 
    20.00511, 20.00512, 20.00513, 20.00515, 20.00517, 20.0052, 20.00522, 
    20.00523, 20.00522, 20.00523, 20.00522, 20.00522, 20.00526, 20.00524, 
    20.00528, 20.00527, 20.00526, 20.00527, 20.00511, 20.0051, 20.00509, 
    20.0051, 20.00508, 20.00509, 20.0051, 20.00513, 20.00513, 20.00514, 
    20.00515, 20.00517, 20.00519, 20.00522, 20.00524, 20.00524, 20.00524, 
    20.00524, 20.00523, 20.00524, 20.00525, 20.00524, 20.00527, 20.00526, 
    20.00527, 20.00527, 20.00511, 20.00511, 20.00511, 20.00512, 20.00511, 
    20.00514, 20.00515, 20.00518, 20.00517, 20.00519, 20.00517, 20.00517, 
    20.00519, 20.00517, 20.00521, 20.00518, 20.00524, 20.00521, 20.00524, 
    20.00524, 20.00525, 20.00526, 20.00527, 20.00529, 20.00528, 20.0053, 
    20.00513, 20.00514, 20.00514, 20.00515, 20.00516, 20.00517, 20.0052, 
    20.00519, 20.00521, 20.00521, 20.00518, 20.0052, 20.00514, 20.00515, 
    20.00515, 20.00513, 20.00519, 20.00516, 20.00522, 20.0052, 20.00525, 
    20.00523, 20.00528, 20.0053, 20.00532, 20.00535, 20.00514, 20.00513, 
    20.00515, 20.00517, 20.00518, 20.0052, 20.00521, 20.00521, 20.00522, 
    20.00523, 20.00521, 20.00523, 20.00516, 20.0052, 20.00513, 20.00515, 
    20.00517, 20.00516, 20.00519, 20.0052, 20.00522, 20.00521, 20.0053, 
    20.00526, 20.00537, 20.00533, 20.00513, 20.00514, 20.00517, 20.00516, 
    20.00521, 20.00522, 20.00522, 20.00524, 20.00524, 20.00524, 20.00523, 
    20.00524, 20.0052, 20.00522, 20.00517, 20.00518, 20.00518, 20.00517, 
    20.00519, 20.00521, 20.00521, 20.00522, 20.00524, 20.00521, 20.0053, 
    20.00524, 20.00515, 20.00517, 20.00517, 20.00517, 20.00521, 20.0052, 
    20.00524, 20.00523, 20.00525, 20.00524, 20.00524, 20.00523, 20.00522, 
    20.0052, 20.00518, 20.00517, 20.00517, 20.00519, 20.00521, 20.00524, 
    20.00523, 20.00525, 20.0052, 20.00522, 20.00521, 20.00524, 20.00519, 
    20.00523, 20.00518, 20.00518, 20.0052, 20.00522, 20.00523, 20.00524, 
    20.00523, 20.00521, 20.00521, 20.0052, 20.00519, 20.00518, 20.00517, 
    20.00518, 20.00519, 20.00521, 20.00523, 20.00526, 20.00526, 20.00529, 
    20.00527, 20.0053, 20.00527, 20.00532, 20.00523, 20.00527, 20.0052, 
    20.00521, 20.00522, 20.00525, 20.00524, 20.00525, 20.00521, 20.00519, 
    20.00518, 20.00517, 20.00518, 20.00518, 20.00519, 20.00519, 20.00521, 
    20.0052, 20.00524, 20.00525, 20.0053, 20.00532, 20.00535, 20.00536, 
    20.00537, 20.00537,
  20.00437, 20.00439, 20.00439, 20.0044, 20.00439, 20.00441, 20.00438, 
    20.00439, 20.00438, 20.00437, 20.00444, 20.0044, 20.00447, 20.00445, 
    20.0045, 20.00447, 20.00451, 20.0045, 20.00452, 20.00451, 20.00454, 
    20.00452, 20.00456, 20.00454, 20.00454, 20.00452, 20.00441, 20.00443, 
    20.00441, 20.00441, 20.00441, 20.00439, 20.00439, 20.00437, 20.00437, 
    20.00438, 20.00441, 20.0044, 20.00443, 20.00443, 20.00446, 20.00444, 
    20.00449, 20.00448, 20.00451, 20.00451, 20.00451, 20.00451, 20.00451, 
    20.0045, 20.00451, 20.00449, 20.00445, 20.00446, 20.00442, 20.00439, 
    20.00438, 20.00436, 20.00437, 20.00437, 20.00438, 20.0044, 20.00441, 
    20.00442, 20.00443, 20.00445, 20.00447, 20.00449, 20.00449, 20.0045, 
    20.0045, 20.00452, 20.00451, 20.00452, 20.0045, 20.00451, 20.00448, 
    20.00449, 20.00443, 20.00441, 20.0044, 20.00439, 20.00437, 20.00438, 
    20.00438, 20.00439, 20.0044, 20.00439, 20.00442, 20.00441, 20.00447, 
    20.00444, 20.0045, 20.00449, 20.00451, 20.0045, 20.00451, 20.0045, 
    20.00452, 20.00453, 20.00452, 20.00454, 20.0045, 20.00451, 20.00439, 
    20.00439, 20.0044, 20.00438, 20.00438, 20.00437, 20.00438, 20.00439, 
    20.0044, 20.00441, 20.00441, 20.00443, 20.00445, 20.00447, 20.00449, 
    20.0045, 20.00449, 20.0045, 20.00449, 20.00449, 20.00453, 20.00451, 
    20.00454, 20.00454, 20.00452, 20.00454, 20.00439, 20.00439, 20.00438, 
    20.00439, 20.00437, 20.00438, 20.00439, 20.00441, 20.00442, 20.00442, 
    20.00443, 20.00444, 20.00447, 20.00449, 20.0045, 20.0045, 20.0045, 
    20.00451, 20.0045, 20.00451, 20.00451, 20.00451, 20.00454, 20.00453, 
    20.00454, 20.00453, 20.00439, 20.0044, 20.0044, 20.0044, 20.0044, 
    20.00442, 20.00443, 20.00446, 20.00444, 20.00446, 20.00445, 20.00445, 
    20.00447, 20.00445, 20.00449, 20.00446, 20.00451, 20.00448, 20.00451, 
    20.0045, 20.00451, 20.00452, 20.00453, 20.00455, 20.00454, 20.00456, 
    20.00441, 20.00442, 20.00442, 20.00443, 20.00443, 20.00445, 20.00447, 
    20.00446, 20.00448, 20.00448, 20.00446, 20.00447, 20.00443, 20.00443, 
    20.00443, 20.00441, 20.00447, 20.00444, 20.00449, 20.00447, 20.00452, 
    20.0045, 20.00454, 20.00456, 20.00458, 20.0046, 20.00442, 20.00442, 
    20.00443, 20.00444, 20.00446, 20.00447, 20.00448, 20.00448, 20.00449, 
    20.0045, 20.00448, 20.0045, 20.00443, 20.00447, 20.00442, 20.00443, 
    20.00444, 20.00444, 20.00446, 20.00447, 20.00449, 20.00448, 20.00455, 
    20.00452, 20.00461, 20.00459, 20.00442, 20.00442, 20.00445, 20.00444, 
    20.00448, 20.00449, 20.00449, 20.0045, 20.0045, 20.00451, 20.0045, 
    20.00451, 20.00447, 20.00449, 20.00445, 20.00446, 20.00445, 20.00445, 
    20.00447, 20.00448, 20.00448, 20.00449, 20.0045, 20.00448, 20.00456, 
    20.00451, 20.00443, 20.00445, 20.00445, 20.00444, 20.00448, 20.00447, 
    20.00451, 20.0045, 20.00452, 20.00451, 20.00451, 20.0045, 20.00449, 
    20.00447, 20.00446, 20.00444, 20.00445, 20.00446, 20.00448, 20.0045, 
    20.0045, 20.00451, 20.00447, 20.00449, 20.00448, 20.0045, 20.00446, 
    20.0045, 20.00446, 20.00446, 20.00447, 20.00449, 20.0045, 20.0045, 
    20.0045, 20.00448, 20.00448, 20.00447, 20.00447, 20.00446, 20.00445, 
    20.00446, 20.00446, 20.00448, 20.0045, 20.00452, 20.00452, 20.00455, 
    20.00453, 20.00456, 20.00453, 20.00458, 20.0045, 20.00453, 20.00447, 
    20.00448, 20.00449, 20.00452, 20.0045, 20.00452, 20.00448, 20.00446, 
    20.00446, 20.00445, 20.00446, 20.00445, 20.00446, 20.00446, 20.00448, 
    20.00447, 20.00451, 20.00452, 20.00455, 20.00458, 20.0046, 20.00461, 
    20.00461, 20.00461,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N =
  0.5258222, 0.5258228, 0.5258227, 0.5258232, 0.5258229, 0.5258232, 
    0.5258223, 0.5258228, 0.5258225, 0.5258223, 0.5258241, 0.5258232, 
    0.525825, 0.5258244, 0.5258258, 0.5258249, 0.525826, 0.5258258, 
    0.5258265, 0.5258263, 0.5258271, 0.5258265, 0.5258275, 0.5258269, 
    0.5258271, 0.5258265, 0.5258234, 0.525824, 0.5258233, 0.5258234, 
    0.5258234, 0.5258229, 0.5258226, 0.5258222, 0.5258223, 0.5258226, 
    0.5258234, 0.5258232, 0.5258238, 0.5258238, 0.5258246, 0.5258242, 
    0.5258256, 0.5258252, 0.5258263, 0.525826, 0.5258263, 0.5258262, 
    0.5258263, 0.5258259, 0.525826, 0.5258257, 0.5258243, 0.5258247, 
    0.5258235, 0.5258228, 0.5258223, 0.525822, 0.5258221, 0.5258222, 
    0.5258226, 0.5258231, 0.5258234, 0.5258236, 0.5258238, 0.5258245, 
    0.5258248, 0.5258256, 0.5258255, 0.5258257, 0.525826, 0.5258263, 
    0.5258263, 0.5258265, 0.5258257, 0.5258262, 0.5258254, 0.5258256, 
    0.5258239, 0.5258232, 0.5258229, 0.5258227, 0.5258221, 0.5258225, 
    0.5258223, 0.5258228, 0.525823, 0.5258229, 0.5258237, 0.5258234, 
    0.5258248, 0.5258242, 0.5258259, 0.5258255, 0.525826, 0.5258258, 
    0.5258262, 0.5258258, 0.5258265, 0.5258267, 0.5258266, 0.525827, 
    0.5258258, 0.5258263, 0.5258229, 0.5258229, 0.525823, 0.5258226, 
    0.5258226, 0.5258222, 0.5258225, 0.5258226, 0.525823, 0.5258232, 
    0.5258234, 0.5258239, 0.5258244, 0.5258251, 0.5258256, 0.5258259, 
    0.5258257, 0.5258259, 0.5258257, 0.5258256, 0.5258266, 0.525826, 
    0.5258269, 0.5258269, 0.5258265, 0.5258269, 0.5258229, 0.5258228, 
    0.5258224, 0.5258227, 0.5258222, 0.5258225, 0.5258226, 0.5258234, 
    0.5258235, 0.5258237, 0.5258239, 0.5258243, 0.5258249, 0.5258255, 
    0.525826, 0.5258259, 0.525826, 0.5258261, 0.5258258, 0.5258261, 
    0.5258262, 0.525826, 0.5258269, 0.5258266, 0.5258269, 0.5258267, 
    0.5258228, 0.525823, 0.5258229, 0.5258231, 0.525823, 0.5258236, 
    0.5258238, 0.5258246, 0.5258242, 0.5258248, 0.5258243, 0.5258244, 
    0.5258248, 0.5258244, 0.5258254, 0.5258247, 0.5258261, 0.5258253, 
    0.5258261, 0.525826, 0.5258262, 0.5258264, 0.5258267, 0.5258272, 
    0.5258271, 0.5258275, 0.5258233, 0.5258235, 0.5258235, 0.5258238, 
    0.525824, 0.5258244, 0.5258251, 0.5258248, 0.5258253, 0.5258254, 
    0.5258247, 0.5258251, 0.5258237, 0.525824, 0.5258238, 0.5258234, 
    0.5258249, 0.5258241, 0.5258256, 0.5258251, 0.5258264, 0.5258257, 
    0.525827, 0.5258275, 0.525828, 0.5258286, 0.5258237, 0.5258235, 
    0.5258238, 0.5258242, 0.5258247, 0.5258251, 0.5258252, 0.5258253, 
    0.5258256, 0.5258257, 0.5258253, 0.5258258, 0.525824, 0.525825, 
    0.5258235, 0.5258239, 0.5258242, 0.5258241, 0.5258248, 0.525825, 
    0.5258256, 0.5258253, 0.5258274, 0.5258265, 0.525829, 0.5258283, 
    0.5258235, 0.5258237, 0.5258245, 0.5258241, 0.5258252, 0.5258254, 
    0.5258257, 0.5258259, 0.525826, 0.5258262, 0.5258259, 0.5258262, 
    0.5258251, 0.5258256, 0.5258244, 0.5258247, 0.5258245, 0.5258244, 
    0.5258248, 0.5258253, 0.5258254, 0.5258255, 0.5258259, 0.5258252, 
    0.5258275, 0.5258261, 0.525824, 0.5258244, 0.5258244, 0.5258242, 
    0.5258254, 0.525825, 0.5258262, 0.5258259, 0.5258263, 0.5258261, 
    0.525826, 0.5258257, 0.5258255, 0.525825, 0.5258246, 0.5258243, 
    0.5258244, 0.5258247, 0.5258254, 0.525826, 0.5258259, 0.5258263, 
    0.5258251, 0.5258256, 0.5258254, 0.5258259, 0.5258248, 0.5258257, 
    0.5258246, 0.5258247, 0.525825, 0.5258256, 0.5258258, 0.5258259, 
    0.5258259, 0.5258254, 0.5258253, 0.525825, 0.5258249, 0.5258247, 
    0.5258245, 0.5258247, 0.5258248, 0.5258254, 0.5258259, 0.5258264, 
    0.5258266, 0.5258272, 0.5258267, 0.5258275, 0.5258268, 0.5258281, 
    0.5258258, 0.5258268, 0.525825, 0.5258252, 0.5258256, 0.5258263, 
    0.5258259, 0.5258264, 0.5258253, 0.5258247, 0.5258246, 0.5258243, 
    0.5258246, 0.5258245, 0.5258248, 0.5258248, 0.5258254, 0.5258251, 
    0.525826, 0.5258264, 0.5258274, 0.5258281, 0.5258287, 0.525829, 0.525829, 
    0.5258291 ;

 SOIL2N_TNDNCY_VERT_TRANS =
  -1.003089e-36, -5.139921e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, 
    1.798972e-20, 1.28498e-20, 5.139921e-21, 2.569961e-21, 2.569961e-21, 
    -7.709882e-21, 1.798972e-20, -7.709882e-21, -5.139921e-21, 2.569961e-21, 
    1.28498e-20, -7.709882e-21, 2.569961e-21, -2.569961e-21, -5.139921e-21, 
    7.709882e-21, -1.003089e-36, -5.139921e-21, -1.798972e-20, 1.798972e-20, 
    5.139921e-21, 1.027984e-20, 2.569961e-21, -1.003089e-36, -5.139921e-21, 
    -7.709882e-21, 2.569961e-21, -2.055969e-20, -2.569961e-21, -5.139921e-21, 
    1.28498e-20, -5.139921e-21, -1.541976e-20, 2.569961e-21, 2.569961e-21, 
    2.569961e-21, -2.569961e-21, -1.027984e-20, -1.28498e-20, 7.709882e-21, 
    5.139921e-21, -7.709882e-21, 1.798972e-20, -1.027984e-20, 7.709882e-21, 
    -2.569961e-21, -5.139921e-21, -1.798972e-20, 1.027984e-20, -1.027984e-20, 
    5.139921e-21, -7.709882e-21, -1.798972e-20, 1.541976e-20, -5.139921e-21, 
    2.569961e-21, -2.569961e-21, -2.569961e-21, 5.139921e-21, 7.709882e-21, 
    5.139921e-21, -1.027984e-20, 7.709882e-21, 1.027984e-20, 1.28498e-20, 
    -2.569961e-21, 5.139921e-21, 0, -1.28498e-20, -1.541976e-20, 
    -7.709882e-21, -5.139921e-21, 5.139921e-21, -1.027984e-20, 5.139921e-21, 
    -7.709882e-21, -1.003089e-36, 1.541976e-20, 2.569961e-21, 1.027984e-20, 
    -1.027984e-20, 5.139921e-21, -1.28498e-20, 1.541976e-20, -1.541976e-20, 
    1.28498e-20, 5.139921e-21, 1.28498e-20, 1.541976e-20, -2.569961e-21, 
    -5.139921e-21, 1.027984e-20, -5.139921e-21, -2.569961e-21, -2.569961e-21, 
    2.055969e-20, 1.027984e-20, -2.569961e-21, -1.541976e-20, 2.569961e-21, 
    7.709882e-21, -7.709882e-21, 1.28498e-20, 1.003089e-36, 1.027984e-20, 
    -1.027984e-20, 7.709882e-21, 7.709882e-21, -1.027984e-20, 0, 
    -7.709882e-21, 1.541976e-20, 1.28498e-20, -3.597945e-20, 2.569961e-21, 
    1.28498e-20, 2.569961e-21, -1.28498e-20, 0, 5.139921e-21, -1.003089e-36, 
    1.28498e-20, -2.569961e-21, -5.139921e-21, -7.709882e-21, -1.027984e-20, 
    -5.139921e-21, -1.541976e-20, -5.139921e-21, 7.709882e-21, 5.139921e-21, 
    0, 2.055969e-20, 1.027984e-20, -1.003089e-36, -2.569961e-21, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, 7.709882e-21, 2.569961e-21, 
    -7.709882e-21, 2.055969e-20, -1.28498e-20, -7.709882e-21, 1.003089e-36, 
    -1.798972e-20, -1.003089e-36, 0, 7.709882e-21, 5.139921e-21, 
    -5.139921e-21, -1.541976e-20, 5.139921e-21, 1.28498e-20, -7.709882e-21, 
    1.28498e-20, -1.003089e-36, 0, 1.003089e-36, 1.003089e-36, 1.28498e-20, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, 0, 2.569961e-21, 
    -5.139921e-21, 7.709882e-21, 1.28498e-20, -1.28498e-20, -1.003089e-36, 
    1.28498e-20, 7.709882e-21, -5.139921e-21, -1.003089e-36, 0, 
    -2.569961e-21, 5.139921e-21, 2.569961e-21, 1.003089e-36, -1.027984e-20, 
    -5.139921e-21, -1.003089e-36, -1.027984e-20, -2.569961e-21, 
    -2.569961e-21, -1.003089e-36, 2.569961e-21, 1.027984e-20, -2.569961e-21, 
    -1.541976e-20, 5.139921e-21, -5.139921e-21, 5.139921e-21, 1.027984e-20, 
    5.139921e-21, -1.003089e-36, -7.709882e-21, -1.027984e-20, -1.541976e-20, 
    -1.28498e-20, 1.027984e-20, -7.709882e-21, -5.139921e-21, -1.798972e-20, 
    1.28498e-20, -2.569961e-21, -5.139921e-21, -7.709882e-21, 1.027984e-20, 
    -7.709882e-21, 2.569961e-21, -2.569961e-21, -2.055969e-20, 2.055969e-20, 
    -2.569961e-21, -7.709882e-21, 1.541976e-20, 5.139921e-21, 0, 
    -7.709882e-21, -2.569961e-21, 5.139921e-21, 1.541976e-20, -7.709882e-21, 
    -1.28498e-20, -2.569961e-21, -2.312965e-20, -7.709882e-21, 5.139921e-21, 
    7.709882e-21, 7.709882e-21, 1.003089e-36, 1.027984e-20, -5.139921e-21, 
    7.709882e-21, 1.027984e-20, 5.139921e-21, 5.139921e-21, 2.569961e-21, 
    5.139921e-21, 5.139921e-21, 1.798972e-20, -5.139921e-21, 1.027984e-20, 
    -2.569961e-21, 2.569961e-21, -7.709882e-21, -7.709882e-21, 2.569961e-21, 
    -1.027984e-20, 1.027984e-20, 7.709882e-21, 5.139921e-21, 1.28498e-20, 
    1.28498e-20, 1.541976e-20, -1.28498e-20, 2.569961e-21, 2.312965e-20, 
    2.569961e-21, -2.569961e-21, 7.709882e-21, -7.709882e-21, -1.28498e-20, 
    -7.709882e-21, 7.709882e-21, -1.027984e-20, -1.28498e-20, -5.139921e-21, 
    2.569961e-21, -2.569961e-21, -5.139921e-21, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, 5.139921e-21, -1.027984e-20, 2.569961e-21, 5.139921e-21, 
    -1.541976e-20, 2.569961e-21, 0, 0, -2.569961e-21, -1.003089e-36, 
    -1.798972e-20, 1.003089e-36, 5.139921e-21, -1.541976e-20, 1.027984e-20, 
    5.139921e-21, -7.709882e-21, -1.541976e-20, -1.541976e-20, -7.709882e-21, 
    1.027984e-20, 1.003089e-36, 1.027984e-20, 2.569961e-21, 1.798972e-20, 
    -7.709882e-21, -5.139921e-21, 5.139921e-21, -2.569961e-21, -1.541976e-20, 
    5.139921e-21, 2.569961e-21, 1.541976e-20, 1.003089e-36, -2.569961e-21, 
    1.027984e-20, -1.28498e-20, 7.709882e-21, 2.569961e-21, 5.139921e-21, 
    1.027984e-20, 0, 7.709882e-21, 1.003089e-36, -7.709882e-21, 
    -5.139921e-21, 1.003089e-36, -1.28498e-20, -1.003089e-36, 1.027984e-20, 
    -5.139921e-21, 5.139921e-21, -7.709882e-21, -7.709882e-21, 1.541976e-20,
  -5.139921e-21, 2.569961e-21, -2.569961e-21, 2.569961e-21, 7.709882e-21, 
    -2.569961e-21, -2.569961e-21, -1.027984e-20, 2.569961e-21, 2.569961e-21, 
    1.003089e-36, 1.003089e-36, 7.709882e-21, -2.569961e-21, 7.709882e-21, 
    1.798972e-20, -2.569961e-21, -7.709882e-21, -7.709882e-21, 5.139921e-21, 
    5.139921e-21, 1.027984e-20, -2.569961e-21, -5.139921e-21, -7.709882e-21, 
    7.709882e-21, -2.569961e-21, 0, -1.003089e-36, -1.027984e-20, 
    -1.28498e-20, 5.139921e-21, 2.569961e-21, -1.003089e-36, 0, 2.569961e-21, 
    7.709882e-21, -7.709882e-21, 1.027984e-20, -5.139921e-21, 5.139921e-21, 
    -7.709882e-21, 2.569961e-21, -1.28498e-20, 5.139921e-21, -1.28498e-20, 
    -2.569961e-21, 0, -7.709882e-21, -5.139921e-21, 1.027984e-20, 
    -5.139921e-21, -2.569961e-21, 1.003089e-36, 1.003089e-36, -7.709882e-21, 
    2.569961e-21, -5.139921e-21, 1.027984e-20, 5.139921e-21, -1.027984e-20, 
    2.569961e-21, 0, -5.139921e-21, 0, -2.569961e-21, -5.139921e-21, 
    -5.139921e-21, -1.003089e-36, -1.003089e-36, -2.569961e-21, 
    -5.139921e-21, 2.569961e-21, -1.003089e-36, 5.139921e-21, 2.569961e-21, 
    -2.569961e-21, -2.569961e-21, -2.569961e-21, -1.28498e-20, 1.798972e-20, 
    -5.139921e-21, -1.541976e-20, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    5.139921e-21, -2.569961e-21, 1.027984e-20, -7.709882e-21, -1.027984e-20, 
    7.709882e-21, 5.139921e-21, 0, 0, 1.003089e-36, 5.139921e-21, 
    -5.139921e-21, 0, 7.709882e-21, 2.569961e-21, -1.027984e-20, 
    7.709882e-21, 0, 5.139921e-21, 7.709882e-21, -1.027984e-20, 5.139921e-21, 
    -2.569961e-21, 5.139921e-21, 2.569961e-21, -7.709882e-21, -1.027984e-20, 
    1.798972e-20, 1.28498e-20, -1.541976e-20, 7.709882e-21, -7.709882e-21, 
    7.709882e-21, 0, 7.709882e-21, -7.709882e-21, -2.569961e-21, 
    -5.139921e-21, 1.027984e-20, -1.027984e-20, -5.139921e-21, 2.569961e-21, 
    -5.139921e-21, 2.569961e-21, 5.139921e-21, -2.569961e-21, -7.709882e-21, 
    1.027984e-20, -1.027984e-20, -5.139921e-21, 2.569961e-21, 0, 
    1.798972e-20, -1.28498e-20, 2.569961e-21, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, -1.027984e-20, -1.003089e-36, 2.569961e-21, 1.28498e-20, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, -7.709882e-21, -2.569961e-21, 
    -1.027984e-20, 7.709882e-21, 0, 1.003089e-36, 1.28498e-20, -2.569961e-21, 
    5.139921e-21, 5.139921e-21, -7.709882e-21, -2.569961e-21, -2.569961e-21, 
    -1.027984e-20, -2.569961e-21, -5.139921e-21, -7.709882e-21, 0, 
    -7.709882e-21, 5.139921e-21, 5.139921e-21, 5.139921e-21, 0, 
    -5.139921e-21, -2.569961e-21, -2.569961e-21, 0, 2.569961e-21, 
    -1.541976e-20, -1.003089e-36, -5.139921e-21, 7.709882e-21, 2.569961e-21, 
    5.139921e-21, -5.139921e-21, 2.569961e-21, 0, -1.28498e-20, 2.569961e-21, 
    -7.709882e-21, 1.541976e-20, 5.139921e-21, -5.139921e-21, 7.709882e-21, 
    1.003089e-36, 7.709882e-21, 0, 5.139921e-21, -1.027984e-20, 
    -1.027984e-20, 0, -7.709882e-21, -2.569961e-21, -2.569961e-21, 
    1.027984e-20, 5.139921e-21, -1.798972e-20, 0, 7.709882e-21, 
    -2.569961e-21, 7.709882e-21, 1.027984e-20, 5.139921e-21, -2.569961e-21, 
    5.139921e-21, 2.569961e-21, 7.709882e-21, -1.003089e-36, 2.569961e-21, 
    -7.709882e-21, -2.569961e-21, -5.139921e-21, 1.027984e-20, -1.027984e-20, 
    5.139921e-21, -5.139921e-21, 2.569961e-21, -1.28498e-20, 1.027984e-20, 
    5.139921e-21, 2.569961e-21, -1.28498e-20, 2.569961e-21, 2.569961e-21, 
    -5.139921e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, 
    1.28498e-20, 1.027984e-20, 5.139921e-21, 1.027984e-20, 2.569961e-21, 
    -2.569961e-21, 7.709882e-21, 2.569961e-21, -2.569961e-21, 1.28498e-20, 
    7.709882e-21, 1.28498e-20, -1.28498e-20, 1.003089e-36, -2.569961e-21, 0, 
    -7.709882e-21, -5.139921e-21, 2.569961e-21, -2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 2.569961e-21, 5.139921e-21, 1.027984e-20, -2.569961e-21, 
    5.139921e-21, 7.709882e-21, 2.569961e-21, -2.569961e-21, -1.003089e-36, 
    -5.139921e-21, 0, -2.569961e-21, -5.139921e-21, -1.027984e-20, 
    -7.709882e-21, 5.139921e-21, 0, 1.003089e-36, -2.569961e-21, 
    -2.569961e-21, 5.139921e-21, -7.709882e-21, -1.28498e-20, -5.139921e-21, 
    -1.28498e-20, -5.139921e-21, 5.139921e-21, -1.28498e-20, 0, 
    -2.569961e-21, 7.709882e-21, -7.709882e-21, -7.709882e-21, -5.139921e-21, 
    -7.709882e-21, 7.709882e-21, -5.139921e-21, 2.569961e-21, 2.569961e-21, 
    0, 0, 7.709882e-21, -7.709882e-21, 5.139921e-21, 1.027984e-20, 
    2.569961e-21, 5.139921e-21, -5.139921e-21, 7.709882e-21, 0, 1.027984e-20, 
    5.139921e-21, 0, 2.569961e-21, 1.003089e-36, -1.027984e-20, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, -7.709882e-21, -2.569961e-21, 
    5.139921e-21, 1.027984e-20, 1.798972e-20, 7.709882e-21, 1.027984e-20, 
    -7.709882e-21, -2.569961e-21, 2.569961e-21, -1.28498e-20, -1.027984e-20, 
    5.139921e-21, 2.569961e-21, 5.139921e-21, 2.569961e-21,
  2.569961e-21, -1.027984e-20, -1.28498e-20, -5.139921e-21, 7.709882e-21, 
    -1.28498e-20, -1.541976e-20, -7.709882e-21, 2.569961e-21, 1.28498e-20, 
    -2.569961e-21, 5.139921e-21, 1.28498e-20, 7.709882e-21, 1.28498e-20, 
    1.027984e-20, 7.709882e-21, 2.569961e-21, 5.139921e-21, 1.003089e-36, 
    1.541976e-20, 2.569961e-21, 1.798972e-20, -2.569961e-21, 2.569961e-21, 
    1.003089e-36, -1.027984e-20, 0, 0, -7.709882e-21, 1.003089e-36, 
    -2.569961e-21, 1.027984e-20, 7.709882e-21, 1.003089e-36, -5.139921e-21, 
    2.569961e-21, 7.709882e-21, 2.569961e-21, 1.003089e-36, -1.027984e-20, 
    -7.709882e-21, 2.569961e-21, 7.709882e-21, -5.139921e-21, 2.569961e-21, 
    -5.139921e-21, 5.139921e-21, -2.569961e-21, -2.569961e-21, -7.709882e-21, 
    7.709882e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, -2.569961e-21, 
    -2.569961e-21, -5.139921e-21, 7.709882e-21, 2.569961e-21, 5.139921e-21, 
    2.569961e-21, 0, -5.139921e-21, -1.027984e-20, 1.798972e-20, 
    -2.569961e-21, 1.027984e-20, 7.709882e-21, 2.569961e-21, -7.709882e-21, 
    7.709882e-21, 2.569961e-21, -2.312965e-20, 7.709882e-21, -2.569961e-21, 
    -5.139921e-21, 5.139921e-21, -5.139921e-21, 7.709882e-21, 5.139921e-21, 
    -5.139921e-21, -2.569961e-21, 2.569961e-21, -1.003089e-36, 1.003089e-36, 
    2.569961e-21, 0, -2.569961e-21, 2.569961e-21, 5.139921e-21, 
    -5.139921e-21, -2.569961e-21, 1.027984e-20, 1.28498e-20, 2.569961e-21, 
    -2.569961e-21, 7.709882e-21, -1.027984e-20, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 1.541976e-20, -2.569961e-21, 1.28498e-20, 7.709882e-21, 
    -7.709882e-21, -5.139921e-21, 1.798972e-20, -2.569961e-21, -5.139921e-21, 
    5.139921e-21, -1.003089e-36, 0, 5.139921e-21, 7.709882e-21, 
    -1.027984e-20, 0, -1.027984e-20, 1.027984e-20, 2.569961e-21, 
    5.139921e-21, -7.709882e-21, -1.027984e-20, -1.28498e-20, 2.569961e-21, 
    1.027984e-20, 7.709882e-21, -1.28498e-20, -5.139921e-21, 1.798972e-20, 
    2.569961e-21, -7.709882e-21, 2.569961e-21, 1.541976e-20, 2.569961e-21, 
    -1.027984e-20, 5.139921e-21, 1.027984e-20, -2.569961e-21, -2.569961e-21, 
    2.569961e-21, 1.28498e-20, -1.798972e-20, -7.709882e-21, 5.139921e-21, 
    -2.569961e-21, -7.709882e-21, -2.569961e-21, 7.709882e-21, 0, 
    1.027984e-20, -1.003089e-36, -1.798972e-20, -1.28498e-20, -1.027984e-20, 
    -2.569961e-21, 1.027984e-20, 0, -2.569961e-21, 5.139921e-21, 
    2.569961e-21, -1.003089e-36, -1.003089e-36, 1.027984e-20, 5.139921e-21, 
    1.027984e-20, -7.709882e-21, -5.139921e-21, 1.541976e-20, -1.28498e-20, 
    -1.027984e-20, 1.027984e-20, -1.027984e-20, -2.569961e-21, 1.28498e-20, 
    -1.027984e-20, -1.003089e-36, 2.569961e-21, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, -5.139921e-21, -5.139921e-21, -1.28498e-20, 2.569961e-21, 
    1.541976e-20, -7.709882e-21, -2.569961e-21, 5.139921e-21, 1.798972e-20, 
    7.709882e-21, -5.139921e-21, -7.709882e-21, 0, 1.027984e-20, 
    7.709882e-21, -5.139921e-21, 7.709882e-21, 1.003089e-36, -2.569961e-21, 
    1.003089e-36, -7.709882e-21, 2.569961e-21, -5.139921e-21, -1.28498e-20, 
    2.569961e-21, -1.798972e-20, -2.569961e-21, -2.569961e-21, -2.569961e-21, 
    1.798972e-20, -1.027984e-20, 1.027984e-20, -1.003089e-36, 5.139921e-21, 
    -1.003089e-36, -1.541976e-20, 1.027984e-20, -7.709882e-21, -1.798972e-20, 
    -5.139921e-21, 2.569961e-21, 2.569961e-21, 7.709882e-21, -2.569961e-21, 
    2.569961e-21, -7.709882e-21, 7.709882e-21, 7.709882e-21, 7.709882e-21, 
    -2.569961e-21, 1.541976e-20, -1.003089e-36, -7.709882e-21, -2.569961e-21, 
    7.709882e-21, -7.709882e-21, -2.569961e-21, 7.709882e-21, -5.139921e-21, 
    -1.027984e-20, 0, 7.709882e-21, 1.027984e-20, 1.027984e-20, 
    -1.027984e-20, 2.569961e-21, 1.798972e-20, 0, -5.139921e-21, 
    -1.003089e-36, -7.709882e-21, -2.569961e-21, 1.027984e-20, 0, 
    1.027984e-20, -1.541976e-20, 2.569961e-21, 1.798972e-20, 1.027984e-20, 
    -2.569961e-21, 5.139921e-21, -7.709882e-21, 1.003089e-36, 1.28498e-20, 
    1.798972e-20, 0, 1.541976e-20, 1.027984e-20, -1.027984e-20, 
    -5.139921e-21, 7.709882e-21, 5.139921e-21, 5.139921e-21, 0, 
    -5.139921e-21, -2.569961e-21, 1.28498e-20, 7.709882e-21, 1.798972e-20, 
    2.055969e-20, -2.569961e-21, -5.139921e-21, 0, 7.709882e-21, 
    -2.569961e-21, 1.027984e-20, 7.709882e-21, -1.28498e-20, 2.569961e-21, 
    5.139921e-21, 7.709882e-21, 7.709882e-21, 1.027984e-20, 1.798972e-20, 0, 
    5.139921e-21, 2.569961e-21, -1.003089e-36, 2.569961e-21, -7.709882e-21, 
    7.709882e-21, -2.569961e-21, -5.139921e-21, 0, 7.709882e-21, 
    -1.28498e-20, -2.569961e-21, -5.139921e-21, -5.139921e-21, -7.709882e-21, 
    -5.139921e-21, 0, -7.709882e-21, -2.569961e-20, -2.569961e-21, 0, 
    2.569961e-21, -5.139921e-21, 5.139921e-21, -1.003089e-36, -5.139921e-21, 
    7.709882e-21, 1.798972e-20, 2.569961e-21, 7.709882e-21, -1.28498e-20, 
    -1.28498e-20, -5.139921e-21, -5.139921e-21, -1.798972e-20, 0, 
    -7.709882e-21, 1.28498e-20, -7.709882e-21, -2.569961e-21, 2.569961e-21,
  1.027984e-20, -7.709882e-21, -5.139921e-21, -7.709882e-21, 1.541976e-20, 
    5.139921e-21, -2.569961e-21, 2.569961e-21, -1.003089e-36, -1.003089e-36, 
    -7.709882e-21, -2.569961e-21, 2.569961e-21, 0, 2.569961e-21, 0, 
    2.569961e-21, -2.569961e-21, -5.139921e-21, -1.798972e-20, 1.28498e-20, 
    -1.003089e-36, 7.709882e-21, 2.312965e-20, 1.541976e-20, 1.027984e-20, 
    1.027984e-20, 2.055969e-20, 0, 5.139921e-21, 2.569961e-21, -1.003089e-36, 
    -1.027984e-20, -7.709882e-21, -2.569961e-21, -1.027984e-20, 
    -7.709882e-21, -2.569961e-21, -7.709882e-21, 2.055969e-20, -1.28498e-20, 
    1.28498e-20, -1.003089e-36, 2.312965e-20, -5.139921e-21, -1.027984e-20, 
    5.139921e-21, -1.28498e-20, 2.569961e-21, -5.139921e-21, -1.28498e-20, 
    1.003089e-36, 0, 1.027984e-20, 1.027984e-20, -2.569961e-21, 
    -1.027984e-20, 7.709882e-21, -1.28498e-20, 0, -2.569961e-21, 
    -5.015443e-37, -5.139921e-21, -1.798972e-20, 1.027984e-20, -2.569961e-21, 
    5.139921e-21, -1.541976e-20, 5.139921e-21, 1.541976e-20, 0, -1.28498e-20, 
    7.709882e-21, -2.569961e-21, -2.569961e-21, -2.569961e-21, 1.541976e-20, 
    -1.541976e-20, 2.569961e-21, -2.569961e-21, -1.003089e-36, 1.28498e-20, 
    -2.569961e-21, 1.28498e-20, 0, 5.139921e-21, 2.569961e-21, 0, 
    -2.569961e-21, 2.569961e-21, 1.798972e-20, 5.139921e-21, -1.28498e-20, 
    -1.003089e-36, -7.709882e-21, -7.709882e-21, -2.569961e-21, 1.541976e-20, 
    0, 5.139921e-21, -2.569961e-21, -7.709882e-21, 7.709882e-21, 
    1.541976e-20, 2.569961e-21, 5.139921e-21, 1.027984e-20, 1.003089e-36, 
    -1.28498e-20, -2.569961e-21, -5.139921e-21, -1.541976e-20, -7.709882e-21, 
    -2.569961e-21, 2.569961e-21, -1.28498e-20, -1.003089e-36, 2.055969e-20, 
    -5.139921e-21, -2.569961e-21, 2.055969e-20, -1.28498e-20, -2.569961e-21, 
    -2.569961e-21, 7.709882e-21, -1.541976e-20, 5.139921e-21, -7.709882e-21, 
    -1.28498e-20, -1.798972e-20, -1.798972e-20, 1.003089e-36, -2.569961e-21, 
    0, 1.28498e-20, 7.709882e-21, 5.139921e-21, -5.139921e-21, 1.798972e-20, 
    -1.027984e-20, 2.569961e-21, 1.027984e-20, -7.709882e-21, -1.28498e-20, 
    -5.139921e-21, -1.003089e-36, 2.569961e-21, 1.28498e-20, 5.139921e-21, 
    -1.28498e-20, -1.798972e-20, 1.28498e-20, -2.569961e-21, -1.027984e-20, 
    2.569961e-21, -1.003089e-36, 2.569961e-21, 1.28498e-20, -1.541976e-20, 
    1.28498e-20, 7.709882e-21, 1.027984e-20, -7.709882e-21, 1.541976e-20, 
    2.312965e-20, 5.139921e-21, -1.027984e-20, -1.28498e-20, 5.139921e-21, 
    5.139921e-21, 7.709882e-21, 1.28498e-20, 1.28498e-20, -1.28498e-20, 
    1.28498e-20, 2.569961e-21, -2.312965e-20, 1.003089e-36, -7.709882e-21, 
    -2.569961e-21, -2.569961e-21, 0, -1.027984e-20, -5.139921e-21, 
    7.709882e-21, 7.709882e-21, 2.569961e-21, -2.569961e-21, -5.139921e-21, 
    -1.541976e-20, 5.139921e-21, 2.569961e-21, 1.003089e-36, -7.709882e-21, 
    2.569961e-21, 7.709882e-21, -1.027984e-20, 7.709882e-21, 7.709882e-21, 
    -1.027984e-20, 1.003089e-36, -1.798972e-20, 1.28498e-20, -7.709882e-21, 
    7.709882e-21, -5.139921e-21, 1.003089e-36, -2.569961e-21, 5.139921e-21, 
    -5.139921e-21, -5.139921e-21, -1.28498e-20, 5.139921e-21, 2.055969e-20, 
    -1.027984e-20, -2.569961e-21, 2.569961e-21, 5.139921e-21, -2.569961e-21, 
    2.569961e-20, 1.027984e-20, 5.139921e-21, -1.541976e-20, -5.139921e-21, 
    -7.709882e-21, 0, -1.28498e-20, 1.28498e-20, -1.28498e-20, 1.541976e-20, 
    2.569961e-20, 5.139921e-21, 5.139921e-21, -7.709882e-21, -1.28498e-20, 
    -5.139921e-21, 5.139921e-21, 7.709882e-21, -2.569961e-21, 5.139921e-21, 
    -1.28498e-20, 5.139921e-21, 2.569961e-21, 2.569961e-21, 1.027984e-20, 
    7.709882e-21, 7.709882e-21, 2.569961e-21, -2.569961e-21, 7.709882e-21, 
    1.027984e-20, -1.003089e-36, -1.003089e-36, 1.28498e-20, 1.027984e-20, 
    1.027984e-20, 1.541976e-20, 1.003089e-36, -2.569961e-21, -1.027984e-20, 
    -5.139921e-21, -1.003089e-36, -2.569961e-21, -5.139921e-21, 2.569961e-21, 
    2.569961e-21, -1.003089e-36, -2.569961e-21, -1.28498e-20, 1.541976e-20, 
    -1.541976e-20, 0, 7.709882e-21, -5.139921e-21, -5.139921e-21, 
    -1.027984e-20, -1.027984e-20, 5.139921e-21, -1.541976e-20, -2.312965e-20, 
    2.569961e-21, 2.569961e-21, 7.709882e-21, 7.709882e-21, 0, 1.541976e-20, 
    7.709882e-21, 5.139921e-21, 7.709882e-21, -2.569961e-21, 2.312965e-20, 
    -1.28498e-20, -1.027984e-20, 2.569961e-21, -1.541976e-20, 1.027984e-20, 
    1.798972e-20, -2.569961e-21, 5.139921e-21, -1.28498e-20, -1.003089e-36, 
    5.139921e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, -2.569961e-21, 
    -5.139921e-21, -7.709882e-21, 1.003089e-36, 7.709882e-21, -1.541976e-20, 
    1.003089e-36, 1.027984e-20, 7.709882e-21, 0, 1.28498e-20, 1.003089e-36, 
    2.569961e-21, 1.28498e-20, -2.569961e-21, 1.28498e-20, 7.709882e-21, 
    5.139921e-21, 5.139921e-21, -1.798972e-20, 1.003089e-36, 1.027984e-20, 
    2.569961e-21, 5.139921e-21, 1.28498e-20, -7.709882e-21, -5.139921e-21, 
    -1.798972e-20, 7.709882e-21, 5.139921e-21, -1.541976e-20, -5.139921e-21, 
    -1.027984e-20,
  2.055969e-20, -2.055969e-20, -7.709882e-21, 5.139921e-21, 2.569961e-21, 
    -1.003089e-36, 2.055969e-20, 2.569961e-21, -5.139921e-21, 7.709882e-21, 
    -1.027984e-20, 2.569961e-21, -1.027984e-20, 5.139921e-21, -1.027984e-20, 
    -2.569961e-21, 7.709882e-21, 2.569961e-21, 1.541976e-20, -1.027984e-20, 
    1.027984e-20, 1.003089e-36, -5.139921e-21, -1.003089e-36, 1.027984e-20, 
    2.569961e-21, -2.569961e-21, -7.709882e-21, 1.541976e-20, 1.28498e-20, 
    1.027984e-20, 5.139921e-21, 2.055969e-20, 0, -5.139921e-21, 2.312965e-20, 
    2.569961e-21, -1.798972e-20, 0, 1.28498e-20, 2.569961e-21, 1.027984e-20, 
    5.139921e-21, 1.798972e-20, -2.569961e-21, 7.709882e-21, 2.569961e-21, 
    -1.027984e-20, 5.139921e-21, 2.569961e-21, -2.569961e-21, 0, 
    1.027984e-20, -5.139921e-21, -5.139921e-21, -2.569961e-21, -2.055969e-20, 
    -1.027984e-20, 1.003089e-36, 1.541976e-20, 5.139921e-21, -1.003089e-36, 
    -1.541976e-20, -5.139921e-21, -2.569961e-21, 0, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, 2.569961e-21, 7.709882e-21, 2.569961e-21, 
    1.027984e-20, -1.28498e-20, -5.139921e-21, 1.027984e-20, 5.139921e-21, 
    1.28498e-20, 5.139921e-21, -2.569961e-20, 2.569961e-21, -1.027984e-20, 
    5.139921e-21, -2.569961e-21, -7.709882e-21, 1.798972e-20, 1.541976e-20, 
    7.709882e-21, -7.709882e-21, 1.027984e-20, -2.569961e-21, 1.541976e-20, 
    5.139921e-21, -1.027984e-20, 1.027984e-20, -1.027984e-20, 1.28498e-20, 
    7.709882e-21, -7.709882e-21, 5.139921e-21, -2.312965e-20, 2.569961e-21, 
    1.027984e-20, -1.28498e-20, -2.569961e-21, -5.139921e-21, -5.139921e-21, 
    1.003089e-36, -2.055969e-20, -1.027984e-20, -2.055969e-20, 1.027984e-20, 
    -2.569961e-21, 5.139921e-21, -1.027984e-20, 2.055969e-20, 5.139921e-21, 
    2.312965e-20, 7.709882e-21, 1.28498e-20, -7.709882e-21, 2.569961e-21, 
    7.709882e-21, -7.709882e-21, 1.798972e-20, 1.003089e-36, -5.015443e-37, 
    1.28498e-20, 1.798972e-20, -1.027984e-20, 7.709882e-21, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, 2.569961e-21, -1.027984e-20, -2.569961e-21, 
    -7.709882e-21, -1.798972e-20, -1.541976e-20, -1.28498e-20, -2.569961e-21, 
    2.569961e-21, 1.541976e-20, 7.709882e-21, 7.709882e-21, 5.139921e-21, 
    1.28498e-20, -1.003089e-36, 1.003089e-36, -2.569961e-21, 7.709882e-21, 
    1.28498e-20, -1.003089e-36, -2.569961e-21, 7.709882e-21, 0, 
    -1.541976e-20, -2.055969e-20, -5.139921e-21, 1.541976e-20, -1.003089e-36, 
    1.541976e-20, 1.28498e-20, -1.003089e-36, -2.569961e-21, 7.709882e-21, 
    1.798972e-20, -1.003089e-36, -2.569961e-21, -1.28498e-20, 7.709882e-21, 
    2.569961e-21, 1.003089e-36, 1.798972e-20, 1.28498e-20, -5.139921e-21, 
    1.28498e-20, 7.709882e-21, 2.055969e-20, 2.569961e-21, -5.139921e-21, 
    2.569961e-21, -2.055969e-20, -5.139921e-21, -5.139921e-21, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, 5.139921e-21, -2.569961e-21, 5.139921e-21, 
    2.569961e-21, 1.798972e-20, 3.009266e-36, -2.569961e-21, 2.569961e-21, 
    -7.709882e-21, -1.003089e-36, -1.541976e-20, -1.027984e-20, 1.027984e-20, 
    5.139921e-21, 7.709882e-21, 1.28498e-20, 2.569961e-21, 1.003089e-36, 
    -7.709882e-21, 7.709882e-21, 1.28498e-20, 1.798972e-20, -1.541976e-20, 
    1.28498e-20, -7.709882e-21, 7.709882e-21, -1.541976e-20, -1.28498e-20, 
    -2.569961e-21, -5.139921e-21, 7.709882e-21, -1.027984e-20, -1.28498e-20, 
    -2.569961e-21, 1.798972e-20, 7.709882e-21, -2.055969e-20, 1.027984e-20, 
    -7.709882e-21, -1.541976e-20, 0, 1.003089e-36, -1.027984e-20, 
    1.027984e-20, 1.28498e-20, 7.709882e-21, 2.569961e-21, 2.569961e-21, 
    5.139921e-21, -5.139921e-21, 1.027984e-20, 1.541976e-20, 1.027984e-20, 
    1.798972e-20, -2.569961e-21, -2.569961e-21, 2.055969e-20, 2.055969e-20, 
    5.139921e-21, 0, 2.569961e-21, -2.055969e-20, -2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 1.28498e-20, -5.139921e-21, -7.709882e-21, 
    0, -2.569961e-21, -2.569961e-21, 5.139921e-21, -2.569961e-21, 
    -1.027984e-20, 2.569961e-20, -2.569961e-21, 0, 1.541976e-20, 1.28498e-20, 
    -2.055969e-20, 5.139921e-21, 1.027984e-20, 2.569961e-21, 2.569961e-21, 
    -1.027984e-20, -1.003089e-36, 1.28498e-20, -7.709882e-21, 2.826957e-20, 
    1.28498e-20, 5.139921e-21, -2.312965e-20, 2.569961e-21, -1.027984e-20, 
    -1.027984e-20, -1.541976e-20, -5.139921e-21, -2.055969e-20, 7.709882e-21, 
    5.139921e-21, -2.569961e-21, 5.139921e-21, 2.569961e-21, 2.569961e-21, 
    1.027984e-20, 1.027984e-20, 7.709882e-21, 1.798972e-20, 1.798972e-20, 
    1.027984e-20, -2.569961e-21, 1.541976e-20, 7.709882e-21, -7.709882e-21, 
    7.709882e-21, -7.709882e-21, -7.709882e-21, -5.139921e-21, -5.139921e-21, 
    5.139921e-21, 5.015443e-37, 1.003089e-36, 1.541976e-20, 1.027984e-20, 
    1.027984e-20, 1.541976e-20, -7.709882e-21, -1.28498e-20, -2.569961e-21, 
    -5.139921e-21, 2.569961e-21, -5.139921e-21, -2.569961e-21, -7.709882e-21, 
    -5.139921e-21, 5.139921e-21, 1.027984e-20, -1.541976e-20, 7.709882e-21, 
    2.569961e-21, -2.569961e-21, 2.312965e-20, -5.139921e-21, 5.139921e-21, 
    2.569961e-21, -2.569961e-21, 5.139921e-21, -1.003089e-36, 1.003089e-36,
  6.259414e-29, 6.25942e-29, 6.259419e-29, 6.259425e-29, 6.259422e-29, 
    6.259425e-29, 6.259416e-29, 6.259421e-29, 6.259417e-29, 6.259415e-29, 
    6.259434e-29, 6.259425e-29, 6.259444e-29, 6.259438e-29, 6.259454e-29, 
    6.259443e-29, 6.259456e-29, 6.259453e-29, 6.259461e-29, 6.259459e-29, 
    6.259468e-29, 6.259462e-29, 6.259473e-29, 6.259467e-29, 6.259467e-29, 
    6.259461e-29, 6.259426e-29, 6.259433e-29, 6.259426e-29, 6.259427e-29, 
    6.259427e-29, 6.259422e-29, 6.259419e-29, 6.259414e-29, 6.259414e-29, 
    6.259419e-29, 6.259428e-29, 6.259425e-29, 6.259432e-29, 6.259432e-29, 
    6.259441e-29, 6.259437e-29, 6.259451e-29, 6.259447e-29, 6.259459e-29, 
    6.259456e-29, 6.259459e-29, 6.259458e-29, 6.259459e-29, 6.259454e-29, 
    6.259456e-29, 6.259452e-29, 6.259437e-29, 6.259442e-29, 6.259429e-29, 
    6.259421e-29, 6.259416e-29, 6.259412e-29, 6.259413e-29, 6.259414e-29, 
    6.259419e-29, 6.259423e-29, 6.259427e-29, 6.259429e-29, 6.259432e-29, 
    6.259439e-29, 6.259443e-29, 6.259452e-29, 6.25945e-29, 6.259453e-29, 
    6.259455e-29, 6.25946e-29, 6.259459e-29, 6.259461e-29, 6.259453e-29, 
    6.259458e-29, 6.259449e-29, 6.259452e-29, 6.259432e-29, 6.259425e-29, 
    6.259422e-29, 6.25942e-29, 6.259413e-29, 6.259417e-29, 6.259416e-29, 
    6.25942e-29, 6.259423e-29, 6.259422e-29, 6.259429e-29, 6.259426e-29, 
    6.259443e-29, 6.259436e-29, 6.259455e-29, 6.25945e-29, 6.259456e-29, 
    6.259453e-29, 6.259458e-29, 6.259454e-29, 6.259462e-29, 6.259463e-29, 
    6.259463e-29, 6.259467e-29, 6.259453e-29, 6.259459e-29, 6.259422e-29, 
    6.259422e-29, 6.259423e-29, 6.259418e-29, 6.259418e-29, 6.259414e-29, 
    6.259417e-29, 6.259419e-29, 6.259423e-29, 6.259425e-29, 6.259428e-29, 
    6.259432e-29, 6.259438e-29, 6.259446e-29, 6.259451e-29, 6.259455e-29, 
    6.259452e-29, 6.259455e-29, 6.259452e-29, 6.259451e-29, 6.259463e-29, 
    6.259456e-29, 6.259466e-29, 6.259466e-29, 6.259461e-29, 6.259466e-29, 
    6.259422e-29, 6.25942e-29, 6.259416e-29, 6.259419e-29, 6.259413e-29, 
    6.259417e-29, 6.259419e-29, 6.259426e-29, 6.259428e-29, 6.25943e-29, 
    6.259433e-29, 6.259437e-29, 6.259444e-29, 6.25945e-29, 6.259456e-29, 
    6.259455e-29, 6.259455e-29, 6.259456e-29, 6.259453e-29, 6.259457e-29, 
    6.259458e-29, 6.259456e-29, 6.259466e-29, 6.259463e-29, 6.259466e-29, 
    6.259464e-29, 6.259421e-29, 6.259423e-29, 6.259422e-29, 6.259424e-29, 
    6.259422e-29, 6.259429e-29, 6.259431e-29, 6.259441e-29, 6.259437e-29, 
    6.259443e-29, 6.259437e-29, 6.259438e-29, 6.259443e-29, 6.259438e-29, 
    6.25945e-29, 6.259441e-29, 6.259456e-29, 6.259449e-29, 6.259457e-29, 
    6.259456e-29, 6.259458e-29, 6.259461e-29, 6.259464e-29, 6.259469e-29, 
    6.259468e-29, 6.259472e-29, 6.259426e-29, 6.259429e-29, 6.259429e-29, 
    6.259432e-29, 6.259434e-29, 6.259438e-29, 6.259446e-29, 6.259443e-29, 
    6.259448e-29, 6.259449e-29, 6.259441e-29, 6.259446e-29, 6.259431e-29, 
    6.259433e-29, 6.259432e-29, 6.259426e-29, 6.259444e-29, 6.259435e-29, 
    6.259451e-29, 6.259446e-29, 6.25946e-29, 6.259453e-29, 6.259467e-29, 
    6.259473e-29, 6.259478e-29, 6.259485e-29, 6.259431e-29, 6.259428e-29, 
    6.259432e-29, 6.259437e-29, 6.259441e-29, 6.259446e-29, 6.259447e-29, 
    6.259448e-29, 6.259451e-29, 6.259453e-29, 6.259449e-29, 6.259454e-29, 
    6.259434e-29, 6.259444e-29, 6.259428e-29, 6.259433e-29, 6.259436e-29, 
    6.259435e-29, 6.259443e-29, 6.259444e-29, 6.259452e-29, 6.259448e-29, 
    6.259472e-29, 6.259461e-29, 6.25949e-29, 6.259482e-29, 6.259428e-29, 
    6.259431e-29, 6.259439e-29, 6.259435e-29, 6.259447e-29, 6.25945e-29, 
    6.259452e-29, 6.259455e-29, 6.259456e-29, 6.259458e-29, 6.259455e-29, 
    6.259457e-29, 6.259447e-29, 6.259452e-29, 6.259438e-29, 6.259441e-29, 
    6.25944e-29, 6.259438e-29, 6.259443e-29, 6.259449e-29, 6.259449e-29, 
    6.25945e-29, 6.259455e-29, 6.259447e-29, 6.259473e-29, 6.259457e-29, 
    6.259433e-29, 6.259438e-29, 6.259438e-29, 6.259437e-29, 6.25945e-29, 
    6.259445e-29, 6.259458e-29, 6.259454e-29, 6.259459e-29, 6.259457e-29, 
    6.259456e-29, 6.259453e-29, 6.25945e-29, 6.259445e-29, 6.259441e-29, 
    6.259437e-29, 6.259438e-29, 6.259442e-29, 6.259449e-29, 6.259456e-29, 
    6.259454e-29, 6.259459e-29, 6.259446e-29, 6.259452e-29, 6.259449e-29, 
    6.259455e-29, 6.259443e-29, 6.259453e-29, 6.25944e-29, 6.259441e-29, 
    6.259445e-29, 6.259452e-29, 6.259453e-29, 6.259455e-29, 6.259454e-29, 
    6.259449e-29, 6.259448e-29, 6.259445e-29, 6.259444e-29, 6.259441e-29, 
    6.259439e-29, 6.259441e-29, 6.259443e-29, 6.259449e-29, 6.259455e-29, 
    6.259461e-29, 6.259462e-29, 6.259469e-29, 6.259463e-29, 6.259473e-29, 
    6.259465e-29, 6.259479e-29, 6.259454e-29, 6.259464e-29, 6.259445e-29, 
    6.259447e-29, 6.259451e-29, 6.259459e-29, 6.259455e-29, 6.259461e-29, 
    6.259448e-29, 6.259442e-29, 6.25944e-29, 6.259437e-29, 6.25944e-29, 
    6.25944e-29, 6.259443e-29, 6.259442e-29, 6.259449e-29, 6.259446e-29, 
    6.259456e-29, 6.259461e-29, 6.259472e-29, 6.259479e-29, 6.259486e-29, 
    6.259489e-29, 6.25949e-29, 6.25949e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N_TO_SOIL1N =
  2.194512e-10, 2.204169e-10, 2.202292e-10, 2.21008e-10, 2.20576e-10, 
    2.21086e-10, 2.19647e-10, 2.204552e-10, 2.199393e-10, 2.195382e-10, 
    2.225196e-10, 2.210428e-10, 2.240534e-10, 2.231116e-10, 2.254774e-10, 
    2.239069e-10, 2.257941e-10, 2.254321e-10, 2.265216e-10, 2.262095e-10, 
    2.276031e-10, 2.266657e-10, 2.283254e-10, 2.273792e-10, 2.275272e-10, 
    2.266347e-10, 2.213399e-10, 2.223357e-10, 2.21281e-10, 2.214229e-10, 
    2.213592e-10, 2.205849e-10, 2.201947e-10, 2.193774e-10, 2.195258e-10, 
    2.20126e-10, 2.214868e-10, 2.210249e-10, 2.22189e-10, 2.221627e-10, 
    2.234587e-10, 2.228744e-10, 2.250526e-10, 2.244335e-10, 2.262225e-10, 
    2.257726e-10, 2.262014e-10, 2.260714e-10, 2.262031e-10, 2.255432e-10, 
    2.25826e-10, 2.252453e-10, 2.229838e-10, 2.236485e-10, 2.216661e-10, 
    2.204742e-10, 2.196825e-10, 2.191206e-10, 2.192001e-10, 2.193515e-10, 
    2.201296e-10, 2.208611e-10, 2.214186e-10, 2.217915e-10, 2.221589e-10, 
    2.232712e-10, 2.238598e-10, 2.251778e-10, 2.249399e-10, 2.253429e-10, 
    2.257279e-10, 2.263742e-10, 2.262678e-10, 2.265525e-10, 2.253323e-10, 
    2.261433e-10, 2.248044e-10, 2.251706e-10, 2.222589e-10, 2.211495e-10, 
    2.20678e-10, 2.202653e-10, 2.192611e-10, 2.199546e-10, 2.196812e-10, 
    2.203315e-10, 2.207447e-10, 2.205403e-10, 2.218017e-10, 2.213113e-10, 
    2.238947e-10, 2.22782e-10, 2.256829e-10, 2.249888e-10, 2.258493e-10, 
    2.254102e-10, 2.261626e-10, 2.254854e-10, 2.266585e-10, 2.269139e-10, 
    2.267394e-10, 2.274099e-10, 2.254479e-10, 2.262014e-10, 2.205346e-10, 
    2.20568e-10, 2.207232e-10, 2.200407e-10, 2.199989e-10, 2.193734e-10, 
    2.1993e-10, 2.20167e-10, 2.207687e-10, 2.211246e-10, 2.214629e-10, 
    2.222068e-10, 2.230376e-10, 2.241992e-10, 2.250338e-10, 2.255932e-10, 
    2.252501e-10, 2.25553e-10, 2.252144e-10, 2.250558e-10, 2.268182e-10, 
    2.258286e-10, 2.273134e-10, 2.272313e-10, 2.265593e-10, 2.272405e-10, 
    2.205914e-10, 2.203995e-10, 2.197336e-10, 2.202548e-10, 2.193052e-10, 
    2.198367e-10, 2.201424e-10, 2.213216e-10, 2.215806e-10, 2.218209e-10, 
    2.222954e-10, 2.229043e-10, 2.239725e-10, 2.249018e-10, 2.257502e-10, 
    2.256881e-10, 2.2571e-10, 2.258995e-10, 2.2543e-10, 2.259766e-10, 
    2.260683e-10, 2.258285e-10, 2.272203e-10, 2.268226e-10, 2.272295e-10, 
    2.269706e-10, 2.204619e-10, 2.207847e-10, 2.206103e-10, 2.209382e-10, 
    2.207072e-10, 2.217345e-10, 2.220426e-10, 2.234838e-10, 2.228923e-10, 
    2.238337e-10, 2.229879e-10, 2.231378e-10, 2.238644e-10, 2.230336e-10, 
    2.248506e-10, 2.236188e-10, 2.259069e-10, 2.246768e-10, 2.25984e-10, 
    2.257466e-10, 2.261396e-10, 2.264916e-10, 2.269344e-10, 2.277515e-10, 
    2.275623e-10, 2.282456e-10, 2.212658e-10, 2.216844e-10, 2.216476e-10, 
    2.220856e-10, 2.224096e-10, 2.231118e-10, 2.242381e-10, 2.238146e-10, 
    2.245921e-10, 2.247482e-10, 2.235669e-10, 2.242922e-10, 2.219646e-10, 
    2.223407e-10, 2.221167e-10, 2.212988e-10, 2.239122e-10, 2.22571e-10, 
    2.250476e-10, 2.24321e-10, 2.264414e-10, 2.253869e-10, 2.274581e-10, 
    2.283436e-10, 2.291768e-10, 2.301507e-10, 2.219129e-10, 2.216284e-10, 
    2.221377e-10, 2.228424e-10, 2.234962e-10, 2.243653e-10, 2.244543e-10, 
    2.246171e-10, 2.250388e-10, 2.253935e-10, 2.246686e-10, 2.254824e-10, 
    2.224279e-10, 2.240286e-10, 2.215209e-10, 2.222761e-10, 2.228009e-10, 
    2.225706e-10, 2.237662e-10, 2.240479e-10, 2.25193e-10, 2.246011e-10, 
    2.281251e-10, 2.26566e-10, 2.308922e-10, 2.296832e-10, 2.215291e-10, 
    2.219119e-10, 2.232443e-10, 2.226104e-10, 2.244234e-10, 2.248696e-10, 
    2.252324e-10, 2.256961e-10, 2.257462e-10, 2.26021e-10, 2.255707e-10, 
    2.260032e-10, 2.243672e-10, 2.250983e-10, 2.23092e-10, 2.235803e-10, 
    2.233557e-10, 2.231093e-10, 2.238698e-10, 2.2468e-10, 2.246973e-10, 
    2.249571e-10, 2.256893e-10, 2.244307e-10, 2.283263e-10, 2.259205e-10, 
    2.223294e-10, 2.230668e-10, 2.231721e-10, 2.228865e-10, 2.248249e-10, 
    2.241225e-10, 2.260142e-10, 2.25503e-10, 2.263407e-10, 2.259244e-10, 
    2.258632e-10, 2.253285e-10, 2.249957e-10, 2.241547e-10, 2.234705e-10, 
    2.229279e-10, 2.23054e-10, 2.236501e-10, 2.247296e-10, 2.257507e-10, 
    2.25527e-10, 2.26277e-10, 2.242919e-10, 2.251243e-10, 2.248026e-10, 
    2.256414e-10, 2.238033e-10, 2.253687e-10, 2.234032e-10, 2.235755e-10, 
    2.241086e-10, 2.251808e-10, 2.25418e-10, 2.256712e-10, 2.25515e-10, 
    2.247569e-10, 2.246328e-10, 2.240956e-10, 2.239473e-10, 2.23538e-10, 
    2.231992e-10, 2.235088e-10, 2.238339e-10, 2.247573e-10, 2.255894e-10, 
    2.264966e-10, 2.267186e-10, 2.277787e-10, 2.269158e-10, 2.283397e-10, 
    2.271292e-10, 2.292247e-10, 2.254594e-10, 2.270935e-10, 2.241328e-10, 
    2.244518e-10, 2.250287e-10, 2.263519e-10, 2.256375e-10, 2.264729e-10, 
    2.246279e-10, 2.236707e-10, 2.23423e-10, 2.229609e-10, 2.234335e-10, 
    2.233951e-10, 2.238474e-10, 2.23702e-10, 2.247879e-10, 2.242046e-10, 
    2.258616e-10, 2.264663e-10, 2.28174e-10, 2.292208e-10, 2.302864e-10, 
    2.307568e-10, 2.309e-10, 2.309598e-10 ;

 SOIL2N_TO_SOIL3N =
  1.567509e-11, 1.574406e-11, 1.573065e-11, 1.578629e-11, 1.575543e-11, 
    1.579186e-11, 1.568907e-11, 1.57468e-11, 1.570995e-11, 1.56813e-11, 
    1.589425e-11, 1.578877e-11, 1.600382e-11, 1.593655e-11, 1.610553e-11, 
    1.599335e-11, 1.612815e-11, 1.610229e-11, 1.618011e-11, 1.615782e-11, 
    1.625736e-11, 1.61904e-11, 1.630896e-11, 1.624137e-11, 1.625195e-11, 
    1.61882e-11, 1.581e-11, 1.588112e-11, 1.580578e-11, 1.581592e-11, 
    1.581137e-11, 1.575606e-11, 1.572819e-11, 1.566981e-11, 1.568041e-11, 
    1.572329e-11, 1.582049e-11, 1.578749e-11, 1.587064e-11, 1.586876e-11, 
    1.596134e-11, 1.59196e-11, 1.607519e-11, 1.603097e-11, 1.615875e-11, 
    1.612661e-11, 1.615724e-11, 1.614795e-11, 1.615736e-11, 1.611023e-11, 
    1.613043e-11, 1.608895e-11, 1.592742e-11, 1.597489e-11, 1.58333e-11, 
    1.574816e-11, 1.56916e-11, 1.565147e-11, 1.565715e-11, 1.566796e-11, 
    1.572354e-11, 1.577579e-11, 1.581561e-11, 1.584225e-11, 1.586849e-11, 
    1.594794e-11, 1.598999e-11, 1.608413e-11, 1.606714e-11, 1.609592e-11, 
    1.612342e-11, 1.616958e-11, 1.616198e-11, 1.618232e-11, 1.609516e-11, 
    1.615309e-11, 1.605746e-11, 1.608362e-11, 1.587564e-11, 1.579639e-11, 
    1.576271e-11, 1.573323e-11, 1.566151e-11, 1.571104e-11, 1.569151e-11, 
    1.573796e-11, 1.576748e-11, 1.575288e-11, 1.584298e-11, 1.580795e-11, 
    1.599248e-11, 1.5913e-11, 1.612021e-11, 1.607063e-11, 1.61321e-11, 
    1.610073e-11, 1.615447e-11, 1.61061e-11, 1.618989e-11, 1.620814e-11, 
    1.619567e-11, 1.624356e-11, 1.610342e-11, 1.615724e-11, 1.575247e-11, 
    1.575485e-11, 1.576595e-11, 1.571719e-11, 1.571421e-11, 1.566952e-11, 
    1.570928e-11, 1.572621e-11, 1.576919e-11, 1.579461e-11, 1.581878e-11, 
    1.587191e-11, 1.593125e-11, 1.601423e-11, 1.607384e-11, 1.61138e-11, 
    1.60893e-11, 1.611093e-11, 1.608675e-11, 1.607541e-11, 1.62013e-11, 
    1.613061e-11, 1.623668e-11, 1.62308e-11, 1.618281e-11, 1.623147e-11, 
    1.575653e-11, 1.574283e-11, 1.569526e-11, 1.573248e-11, 1.566466e-11, 
    1.570262e-11, 1.572445e-11, 1.580868e-11, 1.582719e-11, 1.584435e-11, 
    1.587824e-11, 1.592173e-11, 1.599803e-11, 1.606442e-11, 1.612502e-11, 
    1.612058e-11, 1.612214e-11, 1.613568e-11, 1.610214e-11, 1.614118e-11, 
    1.614774e-11, 1.61306e-11, 1.623002e-11, 1.620162e-11, 1.623068e-11, 
    1.621219e-11, 1.574728e-11, 1.577033e-11, 1.575788e-11, 1.57813e-11, 
    1.57648e-11, 1.583818e-11, 1.586018e-11, 1.596313e-11, 1.592088e-11, 
    1.598812e-11, 1.592771e-11, 1.593841e-11, 1.599032e-11, 1.593097e-11, 
    1.606076e-11, 1.597277e-11, 1.613621e-11, 1.604834e-11, 1.614171e-11, 
    1.612475e-11, 1.615283e-11, 1.617797e-11, 1.62096e-11, 1.626796e-11, 
    1.625445e-11, 1.630326e-11, 1.58047e-11, 1.58346e-11, 1.583197e-11, 
    1.586326e-11, 1.58864e-11, 1.593656e-11, 1.601701e-11, 1.598676e-11, 
    1.604229e-11, 1.605344e-11, 1.596907e-11, 1.602087e-11, 1.585461e-11, 
    1.588148e-11, 1.586548e-11, 1.580706e-11, 1.599373e-11, 1.589793e-11, 
    1.607483e-11, 1.602293e-11, 1.617438e-11, 1.609906e-11, 1.624701e-11, 
    1.631026e-11, 1.636978e-11, 1.643934e-11, 1.585092e-11, 1.58306e-11, 
    1.586698e-11, 1.591731e-11, 1.596401e-11, 1.60261e-11, 1.603245e-11, 
    1.604408e-11, 1.60742e-11, 1.609953e-11, 1.604776e-11, 1.610588e-11, 
    1.588771e-11, 1.600204e-11, 1.582292e-11, 1.587686e-11, 1.591435e-11, 
    1.58979e-11, 1.59833e-11, 1.600343e-11, 1.608521e-11, 1.604293e-11, 
    1.629465e-11, 1.618328e-11, 1.64923e-11, 1.640594e-11, 1.58235e-11, 
    1.585085e-11, 1.594602e-11, 1.590074e-11, 1.603024e-11, 1.606212e-11, 
    1.608803e-11, 1.612115e-11, 1.612473e-11, 1.614435e-11, 1.611219e-11, 
    1.614308e-11, 1.602623e-11, 1.607845e-11, 1.593514e-11, 1.597002e-11, 
    1.595398e-11, 1.593638e-11, 1.59907e-11, 1.604857e-11, 1.604981e-11, 
    1.606836e-11, 1.612066e-11, 1.603076e-11, 1.630903e-11, 1.613718e-11, 
    1.588067e-11, 1.593334e-11, 1.594086e-11, 1.592046e-11, 1.605892e-11, 
    1.600875e-11, 1.614387e-11, 1.610736e-11, 1.616719e-11, 1.613746e-11, 
    1.613308e-11, 1.609489e-11, 1.607112e-11, 1.601105e-11, 1.596218e-11, 
    1.592342e-11, 1.593243e-11, 1.597501e-11, 1.605211e-11, 1.612505e-11, 
    1.610907e-11, 1.616264e-11, 1.602085e-11, 1.608031e-11, 1.605733e-11, 
    1.611725e-11, 1.598595e-11, 1.609776e-11, 1.595737e-11, 1.596968e-11, 
    1.600776e-11, 1.608434e-11, 1.610128e-11, 1.611937e-11, 1.610821e-11, 
    1.605407e-11, 1.60452e-11, 1.600683e-11, 1.599624e-11, 1.5967e-11, 
    1.59428e-11, 1.596491e-11, 1.598814e-11, 1.605409e-11, 1.611353e-11, 
    1.617833e-11, 1.619418e-11, 1.62699e-11, 1.620827e-11, 1.630998e-11, 
    1.622351e-11, 1.637319e-11, 1.610424e-11, 1.622096e-11, 1.600949e-11, 
    1.603227e-11, 1.607348e-11, 1.616799e-11, 1.611697e-11, 1.617664e-11, 
    1.604485e-11, 1.597648e-11, 1.595878e-11, 1.592578e-11, 1.595954e-11, 
    1.595679e-11, 1.59891e-11, 1.597872e-11, 1.605628e-11, 1.601462e-11, 
    1.613298e-11, 1.617617e-11, 1.629814e-11, 1.637292e-11, 1.644903e-11, 
    1.648263e-11, 1.649286e-11, 1.649713e-11 ;

 SOIL2N_vr =
  1.818768, 1.818769, 1.818769, 1.81877, 1.818769, 1.81877, 1.818768, 
    1.818769, 1.818768, 1.818768, 1.818772, 1.81877, 1.818775, 1.818773, 
    1.818777, 1.818775, 1.818778, 1.818777, 1.818779, 1.818778, 1.81878, 
    1.818779, 1.818781, 1.81878, 1.81878, 1.818779, 1.818771, 1.818772, 
    1.81877, 1.818771, 1.818771, 1.818769, 1.818769, 1.818767, 1.818768, 
    1.818769, 1.818771, 1.81877, 1.818772, 1.818772, 1.818774, 1.818773, 
    1.818776, 1.818775, 1.818778, 1.818777, 1.818778, 1.818778, 1.818778, 
    1.818777, 1.818778, 1.818777, 1.818773, 1.818774, 1.818771, 1.818769, 
    1.818768, 1.818767, 1.818767, 1.818767, 1.818769, 1.81877, 1.818771, 
    1.818771, 1.818772, 1.818774, 1.818774, 1.818777, 1.818776, 1.818777, 
    1.818777, 1.818778, 1.818778, 1.818779, 1.818777, 1.818778, 1.818776, 
    1.818776, 1.818772, 1.81877, 1.818769, 1.818769, 1.818767, 1.818768, 
    1.818768, 1.818769, 1.81877, 1.818769, 1.818771, 1.81877, 1.818775, 
    1.818773, 1.818777, 1.818776, 1.818778, 1.818777, 1.818778, 1.818777, 
    1.818779, 1.818779, 1.818779, 1.81878, 1.818777, 1.818778, 1.818769, 
    1.818769, 1.818769, 1.818768, 1.818768, 1.818767, 1.818768, 1.818769, 
    1.81877, 1.81877, 1.818771, 1.818772, 1.818773, 1.818775, 1.818776, 
    1.818777, 1.818777, 1.818777, 1.818777, 1.818776, 1.818779, 1.818778, 
    1.81878, 1.81878, 1.818779, 1.81878, 1.818769, 1.818769, 1.818768, 
    1.818769, 1.818767, 1.818768, 1.818769, 1.81877, 1.818771, 1.818771, 
    1.818772, 1.818773, 1.818775, 1.818776, 1.818777, 1.818777, 1.818777, 
    1.818778, 1.818777, 1.818778, 1.818778, 1.818778, 1.81878, 1.818779, 
    1.81878, 1.818779, 1.818769, 1.81877, 1.818769, 1.81877, 1.818769, 
    1.818771, 1.818772, 1.818774, 1.818773, 1.818774, 1.818773, 1.818773, 
    1.818774, 1.818773, 1.818776, 1.818774, 1.818778, 1.818776, 1.818778, 
    1.818777, 1.818778, 1.818779, 1.818779, 1.818781, 1.81878, 1.818781, 
    1.81877, 1.818771, 1.818771, 1.818772, 1.818772, 1.818773, 1.818775, 
    1.818774, 1.818776, 1.818776, 1.818774, 1.818775, 1.818771, 1.818772, 
    1.818772, 1.81877, 1.818775, 1.818772, 1.818776, 1.818775, 1.818779, 
    1.818777, 1.81878, 1.818781, 1.818783, 1.818784, 1.818771, 1.818771, 
    1.818772, 1.818773, 1.818774, 1.818775, 1.818775, 1.818776, 1.818776, 
    1.818777, 1.818776, 1.818777, 1.818772, 1.818775, 1.818771, 1.818772, 
    1.818773, 1.818772, 1.818774, 1.818775, 1.818777, 1.818776, 1.818781, 
    1.818779, 1.818786, 1.818784, 1.818771, 1.818771, 1.818774, 1.818773, 
    1.818775, 1.818776, 1.818777, 1.818777, 1.818777, 1.818778, 1.818777, 
    1.818778, 1.818775, 1.818776, 1.818773, 1.818774, 1.818774, 1.818773, 
    1.818774, 1.818776, 1.818776, 1.818776, 1.818777, 1.818775, 1.818781, 
    1.818778, 1.818772, 1.818773, 1.818773, 1.818773, 1.818776, 1.818775, 
    1.818778, 1.818777, 1.818778, 1.818778, 1.818778, 1.818777, 1.818776, 
    1.818775, 1.818774, 1.818773, 1.818773, 1.818774, 1.818776, 1.818777, 
    1.818777, 1.818778, 1.818775, 1.818776, 1.818776, 1.818777, 1.818774, 
    1.818777, 1.818774, 1.818774, 1.818775, 1.818777, 1.818777, 1.818777, 
    1.818777, 1.818776, 1.818776, 1.818775, 1.818775, 1.818774, 1.818773, 
    1.818774, 1.818774, 1.818776, 1.818777, 1.818779, 1.818779, 1.818781, 
    1.818779, 1.818781, 1.81878, 1.818783, 1.818777, 1.81878, 1.818775, 
    1.818775, 1.818776, 1.818778, 1.818777, 1.818779, 1.818776, 1.818774, 
    1.818774, 1.818773, 1.818774, 1.818774, 1.818774, 1.818774, 1.818776, 
    1.818775, 1.818778, 1.818779, 1.818781, 1.818783, 1.818785, 1.818785, 
    1.818786, 1.818786,
  1.818734, 1.818736, 1.818735, 1.818737, 1.818736, 1.818737, 1.818734, 
    1.818736, 1.818735, 1.818734, 1.81874, 1.818737, 1.818744, 1.818742, 
    1.818747, 1.818743, 1.818747, 1.818747, 1.818749, 1.818748, 1.818751, 
    1.818749, 1.818753, 1.818751, 1.818751, 1.818749, 1.818738, 1.81874, 
    1.818738, 1.818738, 1.818738, 1.818736, 1.818735, 1.818734, 1.818734, 
    1.818735, 1.818738, 1.818737, 1.81874, 1.81874, 1.818742, 1.818741, 
    1.818746, 1.818744, 1.818748, 1.818747, 1.818748, 1.818748, 1.818748, 
    1.818747, 1.818747, 1.818746, 1.818741, 1.818743, 1.818738, 1.818736, 
    1.818734, 1.818733, 1.818733, 1.818734, 1.818735, 1.818737, 1.818738, 
    1.818739, 1.81874, 1.818742, 1.818743, 1.818746, 1.818745, 1.818746, 
    1.818747, 1.818748, 1.818748, 1.818749, 1.818746, 1.818748, 1.818745, 
    1.818746, 1.81874, 1.818737, 1.818736, 1.818735, 1.818733, 1.818735, 
    1.818734, 1.818736, 1.818737, 1.818736, 1.818739, 1.818738, 1.818743, 
    1.818741, 1.818747, 1.818746, 1.818747, 1.818746, 1.818748, 1.818747, 
    1.818749, 1.81875, 1.818749, 1.818751, 1.818747, 1.818748, 1.818736, 
    1.818736, 1.818737, 1.818735, 1.818735, 1.818734, 1.818735, 1.818735, 
    1.818737, 1.818737, 1.818738, 1.81874, 1.818741, 1.818744, 1.818746, 
    1.818747, 1.818746, 1.818747, 1.818746, 1.818746, 1.818749, 1.818747, 
    1.818751, 1.81875, 1.818749, 1.81875, 1.818736, 1.818736, 1.818734, 
    1.818735, 1.818733, 1.818735, 1.818735, 1.818738, 1.818738, 1.818739, 
    1.81874, 1.818741, 1.818743, 1.818745, 1.818747, 1.818747, 1.818747, 
    1.818748, 1.818747, 1.818748, 1.818748, 1.818747, 1.81875, 1.818749, 
    1.81875, 1.81875, 1.818736, 1.818737, 1.818736, 1.818737, 1.818736, 
    1.818739, 1.818739, 1.818742, 1.818741, 1.818743, 1.818741, 1.818742, 
    1.818743, 1.818741, 1.818745, 1.818743, 1.818748, 1.818745, 1.818748, 
    1.818747, 1.818748, 1.818749, 1.81875, 1.818751, 1.818751, 1.818753, 
    1.818738, 1.818739, 1.818738, 1.818739, 1.81874, 1.818742, 1.818744, 
    1.818743, 1.818745, 1.818745, 1.818743, 1.818744, 1.818739, 1.81874, 
    1.81874, 1.818738, 1.818743, 1.81874, 1.818746, 1.818744, 1.818749, 
    1.818746, 1.818751, 1.818753, 1.818754, 1.818756, 1.818739, 1.818738, 
    1.81874, 1.818741, 1.818742, 1.818744, 1.818744, 1.818745, 1.818746, 
    1.818746, 1.818745, 1.818747, 1.81874, 1.818744, 1.818738, 1.81874, 
    1.818741, 1.81874, 1.818743, 1.818744, 1.818746, 1.818745, 1.818752, 
    1.818749, 1.818758, 1.818756, 1.818738, 1.818739, 1.818742, 1.81874, 
    1.818744, 1.818745, 1.818746, 1.818747, 1.818747, 1.818748, 1.818747, 
    1.818748, 1.818744, 1.818746, 1.818742, 1.818743, 1.818742, 1.818742, 
    1.818743, 1.818745, 1.818745, 1.818745, 1.818747, 1.818744, 1.818753, 
    1.818748, 1.81874, 1.818741, 1.818742, 1.818741, 1.818745, 1.818744, 
    1.818748, 1.818747, 1.818748, 1.818748, 1.818747, 1.818746, 1.818746, 
    1.818744, 1.818742, 1.818741, 1.818741, 1.818743, 1.818745, 1.818747, 
    1.818747, 1.818748, 1.818744, 1.818746, 1.818745, 1.818747, 1.818743, 
    1.818746, 1.818742, 1.818743, 1.818744, 1.818746, 1.818746, 1.818747, 
    1.818747, 1.818745, 1.818745, 1.818744, 1.818743, 1.818743, 1.818742, 
    1.818742, 1.818743, 1.818745, 1.818747, 1.818749, 1.818749, 1.818751, 
    1.81875, 1.818753, 1.81875, 1.818755, 1.818747, 1.81875, 1.818744, 
    1.818744, 1.818746, 1.818748, 1.818747, 1.818749, 1.818745, 1.818743, 
    1.818742, 1.818741, 1.818742, 1.818742, 1.818743, 1.818743, 1.818745, 
    1.818744, 1.818747, 1.818749, 1.818752, 1.818755, 1.818757, 1.818758, 
    1.818758, 1.818758,
  1.818684, 1.818686, 1.818686, 1.818687, 1.818686, 1.818687, 1.818684, 
    1.818686, 1.818685, 1.818684, 1.818691, 1.818687, 1.818694, 1.818692, 
    1.818697, 1.818694, 1.818698, 1.818697, 1.8187, 1.818699, 1.818702, 
    1.8187, 1.818704, 1.818702, 1.818702, 1.8187, 1.818688, 1.81869, 
    1.818688, 1.818688, 1.818688, 1.818686, 1.818685, 1.818684, 1.818684, 
    1.818685, 1.818688, 1.818687, 1.81869, 1.81869, 1.818693, 1.818691, 
    1.818696, 1.818695, 1.818699, 1.818698, 1.818699, 1.818699, 1.818699, 
    1.818698, 1.818698, 1.818697, 1.818692, 1.818693, 1.818689, 1.818686, 
    1.818684, 1.818683, 1.818683, 1.818684, 1.818685, 1.818687, 1.818688, 
    1.818689, 1.81869, 1.818692, 1.818694, 1.818697, 1.818696, 1.818697, 
    1.818698, 1.818699, 1.818699, 1.8187, 1.818697, 1.818699, 1.818696, 
    1.818697, 1.81869, 1.818688, 1.818686, 1.818686, 1.818683, 1.818685, 
    1.818684, 1.818686, 1.818687, 1.818686, 1.818689, 1.818688, 1.818694, 
    1.818691, 1.818698, 1.818696, 1.818698, 1.818697, 1.818699, 1.818697, 
    1.8187, 1.818701, 1.8187, 1.818702, 1.818697, 1.818699, 1.818686, 
    1.818686, 1.818687, 1.818685, 1.818685, 1.818684, 1.818685, 1.818685, 
    1.818687, 1.818688, 1.818688, 1.81869, 1.818692, 1.818695, 1.818696, 
    1.818698, 1.818697, 1.818698, 1.818697, 1.818696, 1.818701, 1.818698, 
    1.818702, 1.818701, 1.8187, 1.818702, 1.818686, 1.818686, 1.818684, 
    1.818686, 1.818683, 1.818685, 1.818685, 1.818688, 1.818689, 1.818689, 
    1.81869, 1.818692, 1.818694, 1.818696, 1.818698, 1.818698, 1.818698, 
    1.818698, 1.818697, 1.818699, 1.818699, 1.818698, 1.818701, 1.818701, 
    1.818701, 1.818701, 1.818686, 1.818687, 1.818686, 1.818687, 1.818687, 
    1.818689, 1.81869, 1.818693, 1.818692, 1.818694, 1.818692, 1.818692, 
    1.818694, 1.818692, 1.818696, 1.818693, 1.818698, 1.818696, 1.818699, 
    1.818698, 1.818699, 1.8187, 1.818701, 1.818703, 1.818702, 1.818704, 
    1.818688, 1.818689, 1.818689, 1.81869, 1.818691, 1.818692, 1.818695, 
    1.818694, 1.818695, 1.818696, 1.818693, 1.818695, 1.818689, 1.81869, 
    1.81869, 1.818688, 1.818694, 1.818691, 1.818696, 1.818695, 1.8187, 
    1.818697, 1.818702, 1.818704, 1.818706, 1.818708, 1.818689, 1.818689, 
    1.81869, 1.818691, 1.818693, 1.818695, 1.818695, 1.818696, 1.818696, 
    1.818697, 1.818696, 1.818697, 1.818691, 1.818694, 1.818689, 1.81869, 
    1.818691, 1.818691, 1.818694, 1.818694, 1.818697, 1.818695, 1.818703, 
    1.8187, 1.81871, 1.818707, 1.818689, 1.818689, 1.818692, 1.818691, 
    1.818695, 1.818696, 1.818697, 1.818698, 1.818698, 1.818699, 1.818698, 
    1.818699, 1.818695, 1.818697, 1.818692, 1.818693, 1.818693, 1.818692, 
    1.818694, 1.818696, 1.818696, 1.818696, 1.818698, 1.818695, 1.818704, 
    1.818698, 1.81869, 1.818692, 1.818692, 1.818692, 1.818696, 1.818694, 
    1.818699, 1.818697, 1.818699, 1.818699, 1.818698, 1.818697, 1.818696, 
    1.818694, 1.818693, 1.818692, 1.818692, 1.818693, 1.818696, 1.818698, 
    1.818698, 1.818699, 1.818695, 1.818697, 1.818696, 1.818698, 1.818694, 
    1.818697, 1.818693, 1.818693, 1.818694, 1.818697, 1.818697, 1.818698, 
    1.818698, 1.818696, 1.818696, 1.818694, 1.818694, 1.818693, 1.818692, 
    1.818693, 1.818694, 1.818696, 1.818698, 1.8187, 1.8187, 1.818703, 
    1.818701, 1.818704, 1.818701, 1.818706, 1.818697, 1.818701, 1.818694, 
    1.818695, 1.818696, 1.818699, 1.818698, 1.8187, 1.818696, 1.818693, 
    1.818693, 1.818692, 1.818693, 1.818693, 1.818694, 1.818693, 1.818696, 
    1.818695, 1.818698, 1.8187, 1.818704, 1.818706, 1.818708, 1.818709, 
    1.81871, 1.81871,
  1.818644, 1.818646, 1.818645, 1.818647, 1.818646, 1.818647, 1.818644, 
    1.818646, 1.818645, 1.818644, 1.818651, 1.818647, 1.818654, 1.818652, 
    1.818657, 1.818654, 1.818658, 1.818657, 1.81866, 1.818659, 1.818662, 
    1.81866, 1.818664, 1.818662, 1.818662, 1.81866, 1.818648, 1.81865, 
    1.818648, 1.818648, 1.818648, 1.818646, 1.818645, 1.818644, 1.818644, 
    1.818645, 1.818648, 1.818647, 1.81865, 1.81865, 1.818653, 1.818651, 
    1.818656, 1.818655, 1.818659, 1.818658, 1.818659, 1.818659, 1.818659, 
    1.818658, 1.818658, 1.818657, 1.818652, 1.818653, 1.818649, 1.818646, 
    1.818644, 1.818643, 1.818643, 1.818644, 1.818645, 1.818647, 1.818648, 
    1.818649, 1.81865, 1.818652, 1.818654, 1.818657, 1.818656, 1.818657, 
    1.818658, 1.818659, 1.818659, 1.81866, 1.818657, 1.818659, 1.818656, 
    1.818657, 1.81865, 1.818648, 1.818647, 1.818646, 1.818643, 1.818645, 
    1.818644, 1.818646, 1.818647, 1.818646, 1.818649, 1.818648, 1.818654, 
    1.818651, 1.818658, 1.818656, 1.818658, 1.818657, 1.818659, 1.818657, 
    1.81866, 1.818661, 1.81866, 1.818662, 1.818657, 1.818659, 1.818646, 
    1.818646, 1.818647, 1.818645, 1.818645, 1.818644, 1.818645, 1.818645, 
    1.818647, 1.818648, 1.818648, 1.81865, 1.818652, 1.818654, 1.818656, 
    1.818658, 1.818657, 1.818658, 1.818657, 1.818656, 1.81866, 1.818658, 
    1.818661, 1.818661, 1.81866, 1.818661, 1.818646, 1.818646, 1.818644, 
    1.818646, 1.818643, 1.818645, 1.818645, 1.818648, 1.818649, 1.818649, 
    1.81865, 1.818652, 1.818654, 1.818656, 1.818658, 1.818658, 1.818658, 
    1.818658, 1.818657, 1.818658, 1.818659, 1.818658, 1.818661, 1.81866, 
    1.818661, 1.818661, 1.818646, 1.818647, 1.818646, 1.818647, 1.818647, 
    1.818649, 1.81865, 1.818653, 1.818652, 1.818654, 1.818652, 1.818652, 
    1.818654, 1.818652, 1.818656, 1.818653, 1.818658, 1.818655, 1.818658, 
    1.818658, 1.818659, 1.81866, 1.818661, 1.818663, 1.818662, 1.818664, 
    1.818648, 1.818649, 1.818649, 1.81865, 1.81865, 1.818652, 1.818655, 
    1.818654, 1.818655, 1.818656, 1.818653, 1.818655, 1.818649, 1.81865, 
    1.81865, 1.818648, 1.818654, 1.818651, 1.818656, 1.818655, 1.81866, 
    1.818657, 1.818662, 1.818664, 1.818666, 1.818668, 1.818649, 1.818649, 
    1.81865, 1.818651, 1.818653, 1.818655, 1.818655, 1.818655, 1.818656, 
    1.818657, 1.818655, 1.818657, 1.81865, 1.818654, 1.818648, 1.81865, 
    1.818651, 1.818651, 1.818653, 1.818654, 1.818657, 1.818655, 1.818663, 
    1.81866, 1.81867, 1.818667, 1.818648, 1.818649, 1.818652, 1.818651, 
    1.818655, 1.818656, 1.818657, 1.818658, 1.818658, 1.818659, 1.818658, 
    1.818658, 1.818655, 1.818656, 1.818652, 1.818653, 1.818653, 1.818652, 
    1.818654, 1.818655, 1.818656, 1.818656, 1.818658, 1.818655, 1.818664, 
    1.818658, 1.81865, 1.818652, 1.818652, 1.818652, 1.818656, 1.818654, 
    1.818659, 1.818657, 1.818659, 1.818658, 1.818658, 1.818657, 1.818656, 
    1.818654, 1.818653, 1.818652, 1.818652, 1.818653, 1.818656, 1.818658, 
    1.818657, 1.818659, 1.818655, 1.818657, 1.818656, 1.818658, 1.818654, 
    1.818657, 1.818653, 1.818653, 1.818654, 1.818657, 1.818657, 1.818658, 
    1.818657, 1.818656, 1.818655, 1.818654, 1.818654, 1.818653, 1.818652, 
    1.818653, 1.818654, 1.818656, 1.818658, 1.81866, 1.81866, 1.818663, 
    1.818661, 1.818664, 1.818661, 1.818666, 1.818657, 1.818661, 1.818654, 
    1.818655, 1.818656, 1.818659, 1.818658, 1.81866, 1.818655, 1.818653, 
    1.818653, 1.818652, 1.818653, 1.818653, 1.818654, 1.818653, 1.818656, 
    1.818654, 1.818658, 1.81866, 1.818663, 1.818666, 1.818668, 1.818669, 
    1.81867, 1.81867,
  1.818579, 1.818581, 1.818581, 1.818582, 1.818581, 1.818582, 1.81858, 
    1.818581, 1.81858, 1.818579, 1.818585, 1.818582, 1.818588, 1.818586, 
    1.818591, 1.818588, 1.818591, 1.818591, 1.818593, 1.818592, 1.818595, 
    1.818593, 1.818596, 1.818594, 1.818595, 1.818593, 1.818583, 1.818585, 
    1.818583, 1.818583, 1.818583, 1.818581, 1.818581, 1.818579, 1.818579, 
    1.818581, 1.818583, 1.818582, 1.818584, 1.818584, 1.818587, 1.818586, 
    1.81859, 1.818589, 1.818592, 1.818591, 1.818592, 1.818592, 1.818592, 
    1.818591, 1.818591, 1.81859, 1.818586, 1.818587, 1.818583, 1.818581, 
    1.81858, 1.818579, 1.818579, 1.818579, 1.818581, 1.818582, 1.818583, 
    1.818584, 1.818584, 1.818587, 1.818588, 1.81859, 1.81859, 1.818591, 
    1.818591, 1.818592, 1.818592, 1.818593, 1.818591, 1.818592, 1.818589, 
    1.81859, 1.818585, 1.818582, 1.818582, 1.818581, 1.818579, 1.81858, 
    1.81858, 1.818581, 1.818582, 1.818581, 1.818584, 1.818583, 1.818588, 
    1.818586, 1.818591, 1.81859, 1.818591, 1.818591, 1.818592, 1.818591, 
    1.818593, 1.818594, 1.818593, 1.818594, 1.818591, 1.818592, 1.818581, 
    1.818581, 1.818582, 1.81858, 1.81858, 1.818579, 1.81858, 1.818581, 
    1.818582, 1.818582, 1.818583, 1.818584, 1.818586, 1.818588, 1.81859, 
    1.818591, 1.81859, 1.818591, 1.81859, 1.81859, 1.818593, 1.818591, 
    1.818594, 1.818594, 1.818593, 1.818594, 1.818581, 1.818581, 1.81858, 
    1.818581, 1.818579, 1.81858, 1.818581, 1.818583, 1.818583, 1.818584, 
    1.818585, 1.818586, 1.818588, 1.81859, 1.818591, 1.818591, 1.818591, 
    1.818592, 1.818591, 1.818592, 1.818592, 1.818591, 1.818594, 1.818593, 
    1.818594, 1.818594, 1.818581, 1.818582, 1.818581, 1.818582, 1.818582, 
    1.818584, 1.818584, 1.818587, 1.818586, 1.818588, 1.818586, 1.818586, 
    1.818588, 1.818586, 1.81859, 1.818587, 1.818592, 1.818589, 1.818592, 
    1.818591, 1.818592, 1.818593, 1.818594, 1.818595, 1.818595, 1.818596, 
    1.818583, 1.818583, 1.818583, 1.818584, 1.818585, 1.818586, 1.818588, 
    1.818588, 1.818589, 1.818589, 1.818587, 1.818588, 1.818584, 1.818585, 
    1.818584, 1.818583, 1.818588, 1.818585, 1.81859, 1.818588, 1.818593, 
    1.818591, 1.818595, 1.818596, 1.818598, 1.8186, 1.818584, 1.818583, 
    1.818584, 1.818586, 1.818587, 1.818589, 1.818589, 1.818589, 1.81859, 
    1.818591, 1.818589, 1.818591, 1.818585, 1.818588, 1.818583, 1.818585, 
    1.818586, 1.818585, 1.818588, 1.818588, 1.81859, 1.818589, 1.818596, 
    1.818593, 1.818601, 1.818599, 1.818583, 1.818584, 1.818586, 1.818585, 
    1.818589, 1.81859, 1.81859, 1.818591, 1.818591, 1.818592, 1.818591, 
    1.818592, 1.818589, 1.81859, 1.818586, 1.818587, 1.818587, 1.818586, 
    1.818588, 1.818589, 1.818589, 1.81859, 1.818591, 1.818589, 1.818596, 
    1.818592, 1.818585, 1.818586, 1.818586, 1.818586, 1.81859, 1.818588, 
    1.818592, 1.818591, 1.818592, 1.818592, 1.818591, 1.818591, 1.81859, 
    1.818588, 1.818587, 1.818586, 1.818586, 1.818587, 1.818589, 1.818591, 
    1.818591, 1.818592, 1.818588, 1.81859, 1.818589, 1.818591, 1.818588, 
    1.818591, 1.818587, 1.818587, 1.818588, 1.81859, 1.818591, 1.818591, 
    1.818591, 1.818589, 1.818589, 1.818588, 1.818588, 1.818587, 1.818586, 
    1.818587, 1.818588, 1.818589, 1.818591, 1.818593, 1.818593, 1.818595, 
    1.818594, 1.818596, 1.818594, 1.818598, 1.818591, 1.818594, 1.818588, 
    1.818589, 1.81859, 1.818592, 1.818591, 1.818593, 1.818589, 1.818587, 
    1.818587, 1.818586, 1.818587, 1.818587, 1.818588, 1.818587, 1.818589, 
    1.818588, 1.818591, 1.818593, 1.818596, 1.818598, 1.8186, 1.818601, 
    1.818601, 1.818601,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2_HR_S1 =
  1.32768e-09, 1.333522e-09, 1.332386e-09, 1.337099e-09, 1.334485e-09, 
    1.33757e-09, 1.328864e-09, 1.333754e-09, 1.330633e-09, 1.328206e-09, 
    1.346243e-09, 1.337309e-09, 1.355523e-09, 1.349825e-09, 1.364139e-09, 
    1.354637e-09, 1.366054e-09, 1.363864e-09, 1.370456e-09, 1.368567e-09, 
    1.376999e-09, 1.371327e-09, 1.381369e-09, 1.375644e-09, 1.37654e-09, 
    1.37114e-09, 1.339107e-09, 1.345131e-09, 1.33875e-09, 1.339609e-09, 
    1.339223e-09, 1.334539e-09, 1.332178e-09, 1.327233e-09, 1.328131e-09, 
    1.331763e-09, 1.339995e-09, 1.3372e-09, 1.344243e-09, 1.344084e-09, 
    1.351925e-09, 1.34839e-09, 1.361568e-09, 1.357823e-09, 1.368646e-09, 
    1.365924e-09, 1.368518e-09, 1.367732e-09, 1.368529e-09, 1.364537e-09, 
    1.366247e-09, 1.362734e-09, 1.349052e-09, 1.353073e-09, 1.34108e-09, 
    1.333869e-09, 1.329079e-09, 1.32568e-09, 1.32616e-09, 1.327076e-09, 
    1.331784e-09, 1.33621e-09, 1.339582e-09, 1.341839e-09, 1.344061e-09, 
    1.350791e-09, 1.354352e-09, 1.362326e-09, 1.360887e-09, 1.363325e-09, 
    1.365653e-09, 1.369564e-09, 1.36892e-09, 1.370643e-09, 1.36326e-09, 
    1.368167e-09, 1.360067e-09, 1.362282e-09, 1.344666e-09, 1.337954e-09, 
    1.335102e-09, 1.332605e-09, 1.32653e-09, 1.330725e-09, 1.329071e-09, 
    1.333006e-09, 1.335506e-09, 1.334269e-09, 1.3419e-09, 1.338934e-09, 
    1.354563e-09, 1.347831e-09, 1.365382e-09, 1.361182e-09, 1.366388e-09, 
    1.363732e-09, 1.368284e-09, 1.364187e-09, 1.371284e-09, 1.372829e-09, 
    1.371773e-09, 1.37583e-09, 1.36396e-09, 1.368518e-09, 1.334235e-09, 
    1.334436e-09, 1.335376e-09, 1.331246e-09, 1.330993e-09, 1.327209e-09, 
    1.330576e-09, 1.33201e-09, 1.33565e-09, 1.337804e-09, 1.339851e-09, 
    1.344351e-09, 1.349377e-09, 1.356405e-09, 1.361454e-09, 1.364839e-09, 
    1.362763e-09, 1.364596e-09, 1.362547e-09, 1.361587e-09, 1.37225e-09, 
    1.366263e-09, 1.375246e-09, 1.374749e-09, 1.370684e-09, 1.374805e-09, 
    1.334578e-09, 1.333417e-09, 1.329388e-09, 1.332541e-09, 1.326797e-09, 
    1.330012e-09, 1.331861e-09, 1.338996e-09, 1.340563e-09, 1.342016e-09, 
    1.344887e-09, 1.348571e-09, 1.355033e-09, 1.360656e-09, 1.365789e-09, 
    1.365413e-09, 1.365545e-09, 1.366692e-09, 1.363852e-09, 1.367158e-09, 
    1.367713e-09, 1.366262e-09, 1.374683e-09, 1.372277e-09, 1.374739e-09, 
    1.373172e-09, 1.333795e-09, 1.335747e-09, 1.334692e-09, 1.336676e-09, 
    1.335278e-09, 1.341494e-09, 1.343357e-09, 1.352077e-09, 1.348498e-09, 
    1.354194e-09, 1.349077e-09, 1.349984e-09, 1.35438e-09, 1.349353e-09, 
    1.360346e-09, 1.352894e-09, 1.366737e-09, 1.359295e-09, 1.367203e-09, 
    1.365767e-09, 1.368144e-09, 1.370274e-09, 1.372953e-09, 1.377896e-09, 
    1.376752e-09, 1.380886e-09, 1.338658e-09, 1.341191e-09, 1.340968e-09, 
    1.343618e-09, 1.345578e-09, 1.349827e-09, 1.356641e-09, 1.354078e-09, 
    1.358782e-09, 1.359726e-09, 1.35258e-09, 1.356968e-09, 1.342886e-09, 
    1.345161e-09, 1.343806e-09, 1.338858e-09, 1.354669e-09, 1.346555e-09, 
    1.361538e-09, 1.357142e-09, 1.36997e-09, 1.363591e-09, 1.376122e-09, 
    1.381479e-09, 1.38652e-09, 1.392412e-09, 1.342573e-09, 1.340852e-09, 
    1.343933e-09, 1.348197e-09, 1.352152e-09, 1.35741e-09, 1.357948e-09, 
    1.358933e-09, 1.361485e-09, 1.36363e-09, 1.359245e-09, 1.364168e-09, 
    1.345689e-09, 1.355373e-09, 1.340202e-09, 1.34477e-09, 1.347945e-09, 
    1.346552e-09, 1.353785e-09, 1.35549e-09, 1.362418e-09, 1.358836e-09, 
    1.380157e-09, 1.370724e-09, 1.396898e-09, 1.389583e-09, 1.340251e-09, 
    1.342567e-09, 1.350628e-09, 1.346793e-09, 1.357761e-09, 1.360461e-09, 
    1.362656e-09, 1.365462e-09, 1.365764e-09, 1.367427e-09, 1.364703e-09, 
    1.367319e-09, 1.357422e-09, 1.361845e-09, 1.349707e-09, 1.352661e-09, 
    1.351302e-09, 1.349811e-09, 1.354412e-09, 1.359314e-09, 1.359419e-09, 
    1.36099e-09, 1.36542e-09, 1.357806e-09, 1.381374e-09, 1.366819e-09, 
    1.345093e-09, 1.349554e-09, 1.350191e-09, 1.348463e-09, 1.36019e-09, 
    1.355941e-09, 1.367386e-09, 1.364293e-09, 1.369361e-09, 1.366843e-09, 
    1.366472e-09, 1.363238e-09, 1.361224e-09, 1.356136e-09, 1.351996e-09, 
    1.348714e-09, 1.349477e-09, 1.353083e-09, 1.359614e-09, 1.365792e-09, 
    1.364439e-09, 1.368976e-09, 1.356966e-09, 1.362002e-09, 1.360056e-09, 
    1.365131e-09, 1.35401e-09, 1.363481e-09, 1.35159e-09, 1.352632e-09, 
    1.355857e-09, 1.362344e-09, 1.363779e-09, 1.365311e-09, 1.364365e-09, 
    1.35978e-09, 1.359028e-09, 1.355778e-09, 1.354881e-09, 1.352405e-09, 
    1.350355e-09, 1.352228e-09, 1.354195e-09, 1.359781e-09, 1.364816e-09, 
    1.370304e-09, 1.371647e-09, 1.378061e-09, 1.37284e-09, 1.381456e-09, 
    1.374131e-09, 1.38681e-09, 1.364029e-09, 1.373916e-09, 1.356004e-09, 
    1.357933e-09, 1.361424e-09, 1.369429e-09, 1.365107e-09, 1.370161e-09, 
    1.358999e-09, 1.353208e-09, 1.351709e-09, 1.348913e-09, 1.351773e-09, 
    1.35154e-09, 1.354277e-09, 1.353397e-09, 1.359967e-09, 1.356438e-09, 
    1.366463e-09, 1.370121e-09, 1.380453e-09, 1.386786e-09, 1.393233e-09, 
    1.396079e-09, 1.396945e-09, 1.397307e-09 ;

 SOIL2_HR_S3 =
  9.483429e-11, 9.525158e-11, 9.517045e-11, 9.550704e-11, 9.532033e-11, 
    9.554073e-11, 9.491888e-11, 9.526815e-11, 9.504519e-11, 9.487185e-11, 
    9.616025e-11, 9.552206e-11, 9.682309e-11, 9.64161e-11, 9.743847e-11, 
    9.675977e-11, 9.757532e-11, 9.741888e-11, 9.78897e-11, 9.775481e-11, 
    9.835704e-11, 9.795195e-11, 9.86692e-11, 9.82603e-11, 9.832427e-11, 
    9.793859e-11, 9.565047e-11, 9.60808e-11, 9.562498e-11, 9.568635e-11, 
    9.565881e-11, 9.532419e-11, 9.515556e-11, 9.480238e-11, 9.48665e-11, 
    9.51259e-11, 9.571394e-11, 9.551432e-11, 9.601738e-11, 9.600602e-11, 
    9.656609e-11, 9.631357e-11, 9.725488e-11, 9.698734e-11, 9.776045e-11, 
    9.756602e-11, 9.775131e-11, 9.769512e-11, 9.775204e-11, 9.74669e-11, 
    9.758907e-11, 9.733815e-11, 9.636086e-11, 9.664809e-11, 9.579144e-11, 
    9.527636e-11, 9.49342e-11, 9.469141e-11, 9.472574e-11, 9.479117e-11, 
    9.512741e-11, 9.544354e-11, 9.568445e-11, 9.584561e-11, 9.600439e-11, 
    9.648505e-11, 9.673942e-11, 9.730899e-11, 9.720619e-11, 9.738033e-11, 
    9.754668e-11, 9.782598e-11, 9.778e-11, 9.790305e-11, 9.737573e-11, 
    9.77262e-11, 9.714763e-11, 9.730588e-11, 9.60476e-11, 9.556817e-11, 
    9.536442e-11, 9.518605e-11, 9.475213e-11, 9.505179e-11, 9.493367e-11, 
    9.521469e-11, 9.539326e-11, 9.530494e-11, 9.585002e-11, 9.56381e-11, 
    9.675449e-11, 9.627363e-11, 9.752728e-11, 9.722728e-11, 9.759918e-11, 
    9.740941e-11, 9.773457e-11, 9.744192e-11, 9.794885e-11, 9.805923e-11, 
    9.79838e-11, 9.827356e-11, 9.742571e-11, 9.775131e-11, 9.530247e-11, 
    9.531687e-11, 9.538397e-11, 9.5089e-11, 9.507096e-11, 9.480063e-11, 
    9.504116e-11, 9.514359e-11, 9.540361e-11, 9.555741e-11, 9.570362e-11, 
    9.602508e-11, 9.638409e-11, 9.688609e-11, 9.724673e-11, 9.748848e-11, 
    9.734024e-11, 9.747111e-11, 9.732481e-11, 9.725624e-11, 9.801788e-11, 
    9.759021e-11, 9.823188e-11, 9.819637e-11, 9.790598e-11, 9.820038e-11, 
    9.532698e-11, 9.524409e-11, 9.495631e-11, 9.518152e-11, 9.477118e-11, 
    9.500088e-11, 9.513296e-11, 9.564254e-11, 9.575449e-11, 9.585831e-11, 
    9.606335e-11, 9.63265e-11, 9.67881e-11, 9.718972e-11, 9.755635e-11, 
    9.752949e-11, 9.753895e-11, 9.762086e-11, 9.741797e-11, 9.765416e-11, 
    9.76938e-11, 9.759016e-11, 9.819162e-11, 9.801979e-11, 9.819562e-11, 
    9.808374e-11, 9.527103e-11, 9.541051e-11, 9.533514e-11, 9.547687e-11, 
    9.537703e-11, 9.5821e-11, 9.595411e-11, 9.657693e-11, 9.632131e-11, 
    9.672813e-11, 9.636263e-11, 9.64274e-11, 9.674141e-11, 9.638238e-11, 
    9.716759e-11, 9.663526e-11, 9.762404e-11, 9.709248e-11, 9.765735e-11, 
    9.755477e-11, 9.772461e-11, 9.787672e-11, 9.806807e-11, 9.842117e-11, 
    9.833941e-11, 9.863469e-11, 9.561844e-11, 9.579935e-11, 9.578341e-11, 
    9.597272e-11, 9.611274e-11, 9.641619e-11, 9.69029e-11, 9.671988e-11, 
    9.705587e-11, 9.712332e-11, 9.661286e-11, 9.692629e-11, 9.592041e-11, 
    9.608294e-11, 9.598616e-11, 9.563271e-11, 9.676206e-11, 9.618249e-11, 
    9.725269e-11, 9.693873e-11, 9.785503e-11, 9.739935e-11, 9.82944e-11, 
    9.867705e-11, 9.903714e-11, 9.9458e-11, 9.589807e-11, 9.577514e-11, 
    9.599524e-11, 9.629975e-11, 9.658227e-11, 9.695788e-11, 9.699631e-11, 
    9.706667e-11, 9.724893e-11, 9.740218e-11, 9.708893e-11, 9.744059e-11, 
    9.612065e-11, 9.681236e-11, 9.572868e-11, 9.605502e-11, 9.62818e-11, 
    9.618231e-11, 9.669895e-11, 9.682073e-11, 9.731554e-11, 9.705975e-11, 
    9.858261e-11, 9.790886e-11, 9.977841e-11, 9.925596e-11, 9.57322e-11, 
    9.589764e-11, 9.647345e-11, 9.619948e-11, 9.698295e-11, 9.71758e-11, 
    9.733256e-11, 9.753297e-11, 9.75546e-11, 9.767334e-11, 9.747876e-11, 
    9.766565e-11, 9.695868e-11, 9.727461e-11, 9.640762e-11, 9.661864e-11, 
    9.652156e-11, 9.641508e-11, 9.674372e-11, 9.709386e-11, 9.710133e-11, 
    9.72136e-11, 9.753001e-11, 9.698612e-11, 9.86696e-11, 9.762995e-11, 
    9.607805e-11, 9.639673e-11, 9.644224e-11, 9.631879e-11, 9.715646e-11, 
    9.685295e-11, 9.767044e-11, 9.74495e-11, 9.781151e-11, 9.763163e-11, 
    9.760516e-11, 9.737412e-11, 9.723027e-11, 9.686687e-11, 9.657117e-11, 
    9.633669e-11, 9.639121e-11, 9.664879e-11, 9.711527e-11, 9.755657e-11, 
    9.74599e-11, 9.7784e-11, 9.692614e-11, 9.728586e-11, 9.714683e-11, 
    9.750934e-11, 9.671501e-11, 9.739148e-11, 9.654211e-11, 9.661658e-11, 
    9.684692e-11, 9.731027e-11, 9.741276e-11, 9.752222e-11, 9.745468e-11, 
    9.712711e-11, 9.707345e-11, 9.684132e-11, 9.677724e-11, 9.660036e-11, 
    9.645393e-11, 9.658772e-11, 9.672823e-11, 9.712724e-11, 9.748684e-11, 
    9.787889e-11, 9.797482e-11, 9.843292e-11, 9.806003e-11, 9.867539e-11, 
    9.815225e-11, 9.905782e-11, 9.743065e-11, 9.813683e-11, 9.68574e-11, 
    9.699523e-11, 9.724455e-11, 9.781635e-11, 9.750764e-11, 9.786866e-11, 
    9.707134e-11, 9.665768e-11, 9.655064e-11, 9.635095e-11, 9.65552e-11, 
    9.653859e-11, 9.673404e-11, 9.667123e-11, 9.714049e-11, 9.688843e-11, 
    9.760449e-11, 9.786581e-11, 9.860375e-11, 9.905614e-11, 9.951661e-11, 
    9.971991e-11, 9.978179e-11, 9.980766e-11 ;

 SOIL3C =
  5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782611, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782613, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782613, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 
    5.782612, 5.782612, 5.782612, 5.782612, 5.782612, 5.782613, 5.782613, 
    5.782613, 5.782613 ;

 SOIL3C_TO_SOIL1C =
  2.618136e-11, 2.629654e-11, 2.627415e-11, 2.636705e-11, 2.631552e-11, 
    2.637635e-11, 2.620471e-11, 2.630112e-11, 2.623957e-11, 2.619173e-11, 
    2.654735e-11, 2.63712e-11, 2.67303e-11, 2.661796e-11, 2.690015e-11, 
    2.671282e-11, 2.693792e-11, 2.689475e-11, 2.70247e-11, 2.698747e-11, 
    2.715369e-11, 2.704188e-11, 2.723985e-11, 2.712698e-11, 2.714464e-11, 
    2.703819e-11, 2.640664e-11, 2.652542e-11, 2.639961e-11, 2.641654e-11, 
    2.640894e-11, 2.631658e-11, 2.627004e-11, 2.617256e-11, 2.619025e-11, 
    2.626185e-11, 2.642416e-11, 2.636906e-11, 2.650792e-11, 2.650478e-11, 
    2.665936e-11, 2.658967e-11, 2.684948e-11, 2.677564e-11, 2.698902e-11, 
    2.693536e-11, 2.69865e-11, 2.697099e-11, 2.69867e-11, 2.6908e-11, 
    2.694172e-11, 2.687246e-11, 2.660272e-11, 2.6682e-11, 2.644555e-11, 
    2.630338e-11, 2.620894e-11, 2.614193e-11, 2.61514e-11, 2.616946e-11, 
    2.626227e-11, 2.634953e-11, 2.641602e-11, 2.64605e-11, 2.650433e-11, 
    2.6637e-11, 2.670721e-11, 2.686441e-11, 2.683604e-11, 2.68841e-11, 
    2.693002e-11, 2.700711e-11, 2.699442e-11, 2.702838e-11, 2.688283e-11, 
    2.697957e-11, 2.681988e-11, 2.686355e-11, 2.651626e-11, 2.638393e-11, 
    2.632769e-11, 2.627846e-11, 2.615869e-11, 2.62414e-11, 2.620879e-11, 
    2.628636e-11, 2.633565e-11, 2.631127e-11, 2.646172e-11, 2.640323e-11, 
    2.671137e-11, 2.657864e-11, 2.692466e-11, 2.684186e-11, 2.694451e-11, 
    2.689213e-11, 2.698188e-11, 2.690111e-11, 2.704102e-11, 2.707149e-11, 
    2.705067e-11, 2.713064e-11, 2.689663e-11, 2.69865e-11, 2.631059e-11, 
    2.631456e-11, 2.633309e-11, 2.625167e-11, 2.624669e-11, 2.617207e-11, 
    2.623846e-11, 2.626674e-11, 2.63385e-11, 2.638096e-11, 2.642131e-11, 
    2.651004e-11, 2.660913e-11, 2.674769e-11, 2.684723e-11, 2.691396e-11, 
    2.687304e-11, 2.690916e-11, 2.686878e-11, 2.684985e-11, 2.706008e-11, 
    2.694204e-11, 2.711914e-11, 2.710934e-11, 2.702919e-11, 2.711045e-11, 
    2.631736e-11, 2.629448e-11, 2.621504e-11, 2.627721e-11, 2.616395e-11, 
    2.622735e-11, 2.62638e-11, 2.640446e-11, 2.643535e-11, 2.646401e-11, 
    2.65206e-11, 2.659323e-11, 2.672064e-11, 2.68315e-11, 2.693269e-11, 
    2.692527e-11, 2.692789e-11, 2.695049e-11, 2.68945e-11, 2.695969e-11, 
    2.697063e-11, 2.694202e-11, 2.710803e-11, 2.70606e-11, 2.710913e-11, 
    2.707825e-11, 2.630191e-11, 2.634041e-11, 2.631961e-11, 2.635873e-11, 
    2.633117e-11, 2.645371e-11, 2.649045e-11, 2.666236e-11, 2.659181e-11, 
    2.670409e-11, 2.660321e-11, 2.662109e-11, 2.670776e-11, 2.660866e-11, 
    2.682539e-11, 2.667846e-11, 2.695137e-11, 2.680465e-11, 2.696057e-11, 
    2.693225e-11, 2.697913e-11, 2.702111e-11, 2.707393e-11, 2.717139e-11, 
    2.714882e-11, 2.723032e-11, 2.63978e-11, 2.644773e-11, 2.644334e-11, 
    2.649559e-11, 2.653423e-11, 2.661799e-11, 2.675233e-11, 2.670181e-11, 
    2.679455e-11, 2.681317e-11, 2.667227e-11, 2.675878e-11, 2.648115e-11, 
    2.652601e-11, 2.64993e-11, 2.640174e-11, 2.671346e-11, 2.655349e-11, 
    2.684888e-11, 2.676222e-11, 2.701513e-11, 2.688935e-11, 2.71364e-11, 
    2.724201e-11, 2.73414e-11, 2.745756e-11, 2.647498e-11, 2.644105e-11, 
    2.65018e-11, 2.658585e-11, 2.666383e-11, 2.67675e-11, 2.677811e-11, 
    2.679753e-11, 2.684784e-11, 2.689013e-11, 2.680368e-11, 2.690074e-11, 
    2.653642e-11, 2.672734e-11, 2.642823e-11, 2.65183e-11, 2.65809e-11, 
    2.655344e-11, 2.669604e-11, 2.672965e-11, 2.686622e-11, 2.679562e-11, 
    2.721595e-11, 2.702999e-11, 2.7546e-11, 2.74018e-11, 2.64292e-11, 
    2.647487e-11, 2.663379e-11, 2.655818e-11, 2.677442e-11, 2.682765e-11, 
    2.687092e-11, 2.692624e-11, 2.693221e-11, 2.696498e-11, 2.691127e-11, 
    2.696286e-11, 2.676773e-11, 2.685492e-11, 2.661562e-11, 2.667387e-11, 
    2.664708e-11, 2.661768e-11, 2.670839e-11, 2.680504e-11, 2.68071e-11, 
    2.683809e-11, 2.692542e-11, 2.67753e-11, 2.723996e-11, 2.6953e-11, 
    2.652466e-11, 2.661262e-11, 2.662518e-11, 2.659111e-11, 2.682232e-11, 
    2.673854e-11, 2.696418e-11, 2.69032e-11, 2.700312e-11, 2.695346e-11, 
    2.694616e-11, 2.688239e-11, 2.684269e-11, 2.674238e-11, 2.666077e-11, 
    2.659605e-11, 2.66111e-11, 2.668219e-11, 2.681095e-11, 2.693275e-11, 
    2.690607e-11, 2.699552e-11, 2.675874e-11, 2.685803e-11, 2.681966e-11, 
    2.691971e-11, 2.670047e-11, 2.688718e-11, 2.665275e-11, 2.66733e-11, 
    2.673688e-11, 2.686477e-11, 2.689306e-11, 2.692327e-11, 2.690463e-11, 
    2.681421e-11, 2.67994e-11, 2.673533e-11, 2.671765e-11, 2.666883e-11, 
    2.662841e-11, 2.666534e-11, 2.670412e-11, 2.681425e-11, 2.69135e-11, 
    2.702171e-11, 2.704819e-11, 2.717463e-11, 2.707171e-11, 2.724156e-11, 
    2.709716e-11, 2.734711e-11, 2.689799e-11, 2.709291e-11, 2.673977e-11, 
    2.677781e-11, 2.684663e-11, 2.700445e-11, 2.691924e-11, 2.701889e-11, 
    2.679882e-11, 2.668465e-11, 2.66551e-11, 2.659998e-11, 2.665636e-11, 
    2.665177e-11, 2.670572e-11, 2.668839e-11, 2.681791e-11, 2.674833e-11, 
    2.694598e-11, 2.70181e-11, 2.722178e-11, 2.734665e-11, 2.747374e-11, 
    2.752985e-11, 2.754693e-11, 2.755407e-11 ;

 SOIL3C_vr =
  20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009,
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00008, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00008, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 
    20.00008, 20.00007, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00007, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00007, 20.00008, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 
    20.00008, 20.00008, 20.00007, 20.00008, 20.00007, 20.00008, 20.00007, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N =
  0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 0.525692, 
    0.525692, 0.525692 ;

 SOIL3N_TNDNCY_VERT_TRANS =
  -1.28498e-20, 1.28498e-20, 1.28498e-20, 0, -7.709882e-21, -1.027984e-20, 
    5.139921e-21, -1.798972e-20, -5.139921e-21, 5.139921e-21, -2.569961e-21, 
    2.569961e-21, 1.003089e-36, 2.569961e-21, 1.027984e-20, 1.003089e-36, 
    -5.139921e-21, -1.28498e-20, -1.798972e-20, 1.28498e-20, 1.027984e-20, 
    5.139921e-21, 5.139921e-21, 7.709882e-21, -1.28498e-20, 1.541976e-20, 
    -1.28498e-20, -2.569961e-21, -5.139921e-21, 1.798972e-20, 2.569961e-21, 
    -1.28498e-20, -2.569961e-21, -2.569961e-21, 1.027984e-20, 5.139921e-21, 
    5.139921e-21, 2.569961e-21, -2.569961e-21, -1.541976e-20, 1.027984e-20, 
    -5.139921e-21, 1.28498e-20, 1.28498e-20, -7.709882e-21, 5.139921e-21, 
    -5.139921e-21, 1.003089e-36, -2.569961e-21, 2.055969e-20, -1.027984e-20, 
    1.798972e-20, 7.709882e-21, -1.027984e-20, 1.003089e-36, -1.28498e-20, 
    -1.027984e-20, 5.139921e-21, 2.569961e-21, -1.027984e-20, -1.027984e-20, 
    -2.569961e-21, 1.027984e-20, -1.798972e-20, -2.569961e-21, 2.569961e-21, 
    1.28498e-20, 5.139921e-21, 1.28498e-20, 2.569961e-21, 2.569961e-21, 
    7.709882e-21, -1.003089e-36, 2.569961e-21, 7.709882e-21, 5.139921e-21, 
    1.027984e-20, 1.28498e-20, 1.027984e-20, 1.28498e-20, 2.569961e-21, 
    5.139921e-21, 5.139921e-21, 7.709882e-21, 2.569961e-20, -2.569961e-21, 
    7.709882e-21, 5.139921e-21, 1.28498e-20, 1.003089e-36, 0, -1.003089e-36, 
    -1.28498e-20, -1.027984e-20, 7.709882e-21, -7.709882e-21, -2.569961e-21, 
    5.139921e-21, 5.139921e-21, -2.569961e-21, -1.28498e-20, -1.027984e-20, 
    7.709882e-21, -2.569961e-21, -2.569961e-21, 7.709882e-21, -7.709882e-21, 
    2.569961e-21, 2.569961e-21, 1.027984e-20, 2.569961e-21, 0, 7.709882e-21, 
    -5.139921e-21, 1.003089e-36, -2.569961e-21, 2.569961e-21, -2.569961e-21, 
    -1.541976e-20, 0, 2.569961e-21, 2.569961e-21, 1.027984e-20, 1.541976e-20, 
    -2.569961e-21, -1.541976e-20, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -1.28498e-20, -1.541976e-20, 2.569961e-21, 7.709882e-21, 
    -7.709882e-21, -1.027984e-20, -7.709882e-21, 2.312965e-20, -1.027984e-20, 
    7.709882e-21, 5.139921e-21, 1.027984e-20, 2.569961e-21, -2.569961e-21, 
    2.569961e-21, -5.139921e-21, -7.709882e-21, -2.569961e-21, 1.027984e-20, 
    1.027984e-20, -2.569961e-21, 2.569961e-21, -1.541976e-20, 5.139921e-21, 
    -1.027984e-20, 0, -5.139921e-21, 5.139921e-21, 2.569961e-21, 
    -2.569961e-21, -1.003089e-36, -1.28498e-20, 3.340949e-20, 1.003089e-36, 
    -2.569961e-21, 5.139921e-21, 7.709882e-21, -2.569961e-21, 7.709882e-21, 
    1.798972e-20, 1.28498e-20, -7.709882e-21, 1.28498e-20, -1.541976e-20, 
    5.139921e-21, -5.139921e-21, 2.569961e-21, -1.003089e-36, 7.709882e-21, 
    -2.055969e-20, 7.709882e-21, 1.28498e-20, -1.027984e-20, 5.139921e-21, 
    1.798972e-20, 1.798972e-20, 1.027984e-20, 5.139921e-21, 5.139921e-21, 
    2.569961e-21, 2.569961e-21, 7.709882e-21, -2.312965e-20, -5.139921e-21, 
    -1.28498e-20, 5.139921e-21, -2.569961e-21, 5.139921e-21, -1.027984e-20, 
    3.340949e-20, 0, -1.798972e-20, -1.027984e-20, -5.139921e-21, 
    -2.569961e-21, -7.709882e-21, -1.027984e-20, 5.139921e-21, 2.569961e-21, 
    1.027984e-20, -5.139921e-21, -1.798972e-20, 1.003089e-36, -2.569961e-21, 
    -1.003089e-36, -7.709882e-21, 2.569961e-21, 7.709882e-21, 1.027984e-20, 
    1.28498e-20, -2.569961e-21, -1.541976e-20, -5.139921e-21, -1.541976e-20, 
    1.28498e-20, 2.569961e-21, -2.569961e-21, -2.569961e-21, 5.139921e-21, 
    5.139921e-21, 5.139921e-21, -7.709882e-21, -1.027984e-20, 2.569961e-21, 
    -1.027984e-20, 1.28498e-20, -1.28498e-20, 2.569961e-21, 7.709882e-21, 
    7.709882e-21, -7.709882e-21, -2.569961e-21, -1.28498e-20, 5.139921e-21, 
    2.569961e-21, 1.28498e-20, -5.139921e-21, -2.569961e-21, -1.027984e-20, 
    0, -1.003089e-36, -1.027984e-20, -1.798972e-20, 7.709882e-21, 
    -7.709882e-21, -1.027984e-20, 7.709882e-21, 1.027984e-20, 1.541976e-20, 
    7.709882e-21, 2.569961e-21, 0, -5.139921e-21, -1.027984e-20, 1.28498e-20, 
    1.541976e-20, -1.541976e-20, 5.139921e-21, -2.569961e-21, 1.28498e-20, 
    -2.569961e-21, 7.709882e-21, -5.139921e-21, 1.28498e-20, 2.569961e-21, 
    2.569961e-21, 0, 2.569961e-21, 2.569961e-21, 1.28498e-20, -2.055969e-20, 
    5.139921e-21, 0, 2.569961e-21, 0, 0, 1.027984e-20, -5.139921e-21, 
    -2.569961e-21, 1.28498e-20, 5.139921e-21, 1.003089e-36, -2.569961e-21, 0, 
    1.003089e-36, 2.569961e-21, -5.139921e-21, -1.28498e-20, 1.003089e-36, 
    -5.139921e-21, -1.003089e-36, -1.003089e-36, 2.569961e-21, -7.709882e-21, 
    1.798972e-20, 5.139921e-21, 1.541976e-20, -7.709882e-21, -7.709882e-21, 
    1.798972e-20, -1.798972e-20, -1.027984e-20, -2.569961e-21, 0, 
    1.28498e-20, -5.139921e-21, 1.28498e-20, -1.027984e-20, -7.709882e-21, 
    1.28498e-20, -1.28498e-20, 1.003089e-36, -1.28498e-20, -1.003089e-36, 
    5.139921e-21, -1.28498e-20, -2.569961e-21, -5.139921e-21, -1.28498e-20, 
    -5.139921e-21, 1.027984e-20, -5.139921e-21, -5.139921e-21, 1.798972e-20, 
    5.139921e-21, 5.139921e-21, -1.027984e-20, 2.569961e-21, -7.709882e-21,
  -1.027984e-20, 1.027984e-20, 7.709882e-21, 2.569961e-21, 2.569961e-21, 
    -5.139921e-21, 7.709882e-21, -2.569961e-21, -2.569961e-21, -2.055969e-20, 
    -2.569961e-21, 1.541976e-20, -2.569961e-21, -1.003089e-36, 0, 
    -1.003089e-36, -7.709882e-21, 1.027984e-20, 7.709882e-21, 2.569961e-21, 
    -7.709882e-21, -2.569961e-21, 5.139921e-21, -2.569961e-21, 2.569961e-21, 
    1.28498e-20, 1.003089e-36, 1.027984e-20, -1.027984e-20, -7.709882e-21, 
    -7.709882e-21, -7.709882e-21, 5.139921e-21, -2.569961e-21, 7.709882e-21, 
    -1.027984e-20, 7.709882e-21, -5.139921e-21, 2.569961e-21, 0, 
    2.826957e-20, 1.003089e-36, 0, -1.027984e-20, 2.569961e-21, 
    -7.709882e-21, 0, 2.569961e-21, 2.569961e-21, 0, -5.139921e-21, 
    5.139921e-21, 1.027984e-20, 0, -2.569961e-21, -2.569961e-21, 
    7.709882e-21, -2.569961e-21, 0, -2.569961e-21, -5.139921e-21, 
    -5.139921e-21, 0, 2.569961e-21, 5.139921e-21, -1.28498e-20, 
    -7.709882e-21, -1.28498e-20, 2.569961e-21, 2.569961e-21, 2.055969e-20, 0, 
    -5.139921e-21, 7.709882e-21, -1.027984e-20, 1.027984e-20, 2.569961e-21, 
    0, -7.709882e-21, -7.709882e-21, 0, -2.569961e-21, 2.569961e-21, 
    7.709882e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, 2.569961e-21, 
    -7.709882e-21, -1.003089e-36, 2.569961e-21, 1.027984e-20, -5.139921e-21, 
    -7.709882e-21, -2.569961e-21, 1.541976e-20, -5.139921e-21, 2.569961e-21, 
    -7.709882e-21, -5.139921e-21, 1.027984e-20, -2.569961e-21, -1.541976e-20, 
    -7.709882e-21, -2.569961e-21, 2.569961e-21, -5.139921e-21, -2.569961e-21, 
    -2.569961e-21, 7.709882e-21, -2.569961e-21, 1.541976e-20, 2.569961e-21, 
    -1.541976e-20, -1.541976e-20, 2.569961e-21, 0, 1.798972e-20, 
    -2.569961e-21, -2.569961e-21, -5.139921e-21, -5.139921e-21, -1.28498e-20, 
    -1.027984e-20, 2.569961e-21, -7.709882e-21, -1.027984e-20, -2.569961e-21, 
    2.569961e-21, 0, -2.569961e-21, 1.027984e-20, 1.28498e-20, 2.569961e-21, 
    0, -7.709882e-21, 5.139921e-21, 5.139921e-21, 7.709882e-21, 
    -2.569961e-21, 1.28498e-20, -2.569961e-21, 1.003089e-36, 2.569961e-21, 
    -1.027984e-20, -1.027984e-20, -5.139921e-21, 7.709882e-21, 1.027984e-20, 
    0, 1.027984e-20, -5.139921e-21, 1.027984e-20, 2.569961e-21, 
    -1.027984e-20, 0, 5.139921e-21, -7.709882e-21, 0, 1.28498e-20, 
    -5.139921e-21, -7.709882e-21, 7.709882e-21, 7.709882e-21, -5.139921e-21, 
    1.28498e-20, -2.569961e-21, -2.569961e-21, -1.027984e-20, -5.139921e-21, 
    1.027984e-20, -7.709882e-21, 2.569961e-21, 5.139921e-21, -1.027984e-20, 
    -1.28498e-20, -1.027984e-20, -2.569961e-21, -5.139921e-21, 1.027984e-20, 
    7.709882e-21, 2.569961e-21, -1.027984e-20, 2.569961e-21, -2.569961e-21, 
    0, 0, 7.709882e-21, 2.569961e-21, -7.709882e-21, -1.003089e-36, 
    2.569961e-21, -1.541976e-20, 5.139921e-21, 7.709882e-21, 5.139921e-21, 
    2.569961e-21, -5.139921e-21, -5.139921e-21, 0, 7.709882e-21, 
    -7.709882e-21, 7.709882e-21, -1.027984e-20, -5.139921e-21, -7.709882e-21, 
    2.569961e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, 5.139921e-21, 
    -1.027984e-20, -1.28498e-20, 1.027984e-20, 5.139921e-21, -1.28498e-20, 
    -1.28498e-20, 1.027984e-20, 1.027984e-20, -1.027984e-20, 2.569961e-21, 
    2.569961e-21, -2.569961e-21, 2.569961e-21, -5.139921e-21, -2.569961e-21, 
    2.569961e-21, 2.569961e-21, -5.139921e-21, 1.027984e-20, -2.569961e-21, 
    -5.139921e-21, 5.139921e-21, -2.569961e-21, -1.027984e-20, -1.28498e-20, 
    -2.569961e-21, -2.569961e-21, 1.027984e-20, 0, 5.139921e-21, 
    1.027984e-20, 1.027984e-20, 1.027984e-20, -7.709882e-21, 5.139921e-21, 
    -1.027984e-20, -1.027984e-20, -7.709882e-21, 7.709882e-21, 0, 
    5.139921e-21, -1.027984e-20, -2.569961e-21, -5.139921e-21, 5.139921e-21, 
    0, -2.569961e-21, -7.709882e-21, -1.28498e-20, 1.027984e-20, 
    1.003089e-36, -1.027984e-20, -1.003089e-36, 5.139921e-21, 2.569961e-21, 
    2.569961e-21, -5.139921e-21, -7.709882e-21, 1.027984e-20, 1.003089e-36, 
    -1.003089e-36, -7.709882e-21, 5.139921e-21, -7.709882e-21, -2.569961e-21, 
    0, 1.28498e-20, 2.569961e-21, 2.569961e-21, 5.139921e-21, -7.709882e-21, 
    -2.569961e-21, 0, 2.569961e-21, -1.28498e-20, 1.027984e-20, 
    -7.709882e-21, -2.569961e-21, -2.569961e-21, 2.569961e-21, -5.139921e-21, 
    1.541976e-20, 7.709882e-21, -1.541976e-20, 2.569961e-21, -1.28498e-20, 
    -5.139921e-21, 5.139921e-21, 1.027984e-20, 1.541976e-20, 7.709882e-21, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, 5.139921e-21, -7.709882e-21, 
    -7.709882e-21, 5.139921e-21, -5.139921e-21, 0, 7.709882e-21, 
    -5.139921e-21, -2.569961e-21, -5.139921e-21, -5.139921e-21, 
    -7.709882e-21, 0, -1.28498e-20, 2.569961e-21, -1.541976e-20, 
    -5.139921e-21, 2.569961e-21, -1.28498e-20, 0, 7.709882e-21, 
    -1.003089e-36, 7.709882e-21, 5.139921e-21, 7.709882e-21, 0, 7.709882e-21, 
    1.027984e-20, 5.139921e-21, 1.28498e-20, 0, 0, -1.027984e-20,
  2.569961e-21, -1.28498e-20, 5.139921e-21, -7.709882e-21, 1.28498e-20, 
    -1.027984e-20, 7.709882e-21, 2.569961e-21, -1.28498e-20, 1.28498e-20, 
    -1.027984e-20, 1.027984e-20, -1.027984e-20, -1.28498e-20, 1.28498e-20, 
    -2.312965e-20, 7.709882e-21, -2.569961e-21, -1.28498e-20, 2.569961e-21, 
    -2.569961e-21, -5.139921e-21, 2.569961e-21, -2.569961e-21, -2.569961e-21, 
    1.003089e-36, -1.003089e-36, 2.569961e-21, 1.027984e-20, -2.569961e-21, 
    -5.139921e-21, 2.569961e-21, 5.139921e-21, 7.709882e-21, 1.027984e-20, 
    -1.798972e-20, -1.027984e-20, -2.569961e-21, 2.569961e-21, 2.569961e-21, 
    5.139921e-21, 7.709882e-21, -1.027984e-20, -2.569961e-21, 2.569961e-21, 
    1.003089e-36, 0, 1.28498e-20, 7.709882e-21, 1.28498e-20, -1.027984e-20, 
    1.027984e-20, 1.28498e-20, 0, 5.139921e-21, -2.569961e-21, 2.569961e-21, 
    2.569961e-21, 1.28498e-20, -5.139921e-21, 5.139921e-21, 1.003089e-36, 
    5.139921e-21, -7.709882e-21, 2.569961e-21, -1.027984e-20, 5.139921e-21, 
    -7.709882e-21, -1.027984e-20, 7.709882e-21, -2.569961e-21, -1.027984e-20, 
    5.139921e-21, 5.139921e-21, -1.027984e-20, 2.569961e-21, 1.027984e-20, 
    -2.569961e-21, -1.541976e-20, -5.139921e-21, 1.027984e-20, 0, 
    5.139921e-21, -7.709882e-21, -1.027984e-20, 0, 7.709882e-21, 
    -7.709882e-21, -5.139921e-21, 0, 0, 1.027984e-20, 1.027984e-20, 
    -5.139921e-21, 2.569961e-21, 5.139921e-21, -1.28498e-20, -2.569961e-21, 
    -7.709882e-21, -5.139921e-21, 1.28498e-20, 5.139921e-21, -5.139921e-21, 
    -1.027984e-20, 2.569961e-21, 7.709882e-21, -5.139921e-21, 5.139921e-21, 
    -1.027984e-20, 1.798972e-20, 0, 1.027984e-20, 7.709882e-21, 
    -2.569961e-21, 2.569961e-21, -5.139921e-21, -5.139921e-21, 2.569961e-21, 
    -1.003089e-36, 5.139921e-21, 2.569961e-21, -5.139921e-21, -7.709882e-21, 
    7.709882e-21, 1.027984e-20, 2.569961e-21, 1.28498e-20, 7.709882e-21, 0, 
    1.027984e-20, -5.139921e-21, -1.027984e-20, -5.139921e-21, -1.003089e-36, 
    -1.541976e-20, 0, -1.541976e-20, -1.28498e-20, 1.541976e-20, 
    5.139921e-21, 2.569961e-21, -1.28498e-20, 2.569961e-21, 0, 5.139921e-21, 
    -2.569961e-21, 5.139921e-21, 7.709882e-21, -5.139921e-21, 2.569961e-21, 
    2.569961e-21, -7.709882e-21, 1.027984e-20, 2.569961e-21, 5.139921e-21, 
    2.312965e-20, -1.28498e-20, 1.28498e-20, -5.139921e-21, 2.569961e-21, 0, 
    7.709882e-21, 5.139921e-21, -1.28498e-20, -1.003089e-36, 2.569961e-21, 
    -7.709882e-21, -2.569961e-21, -1.027984e-20, -2.569961e-21, 
    -5.139921e-21, 2.569961e-21, 7.709882e-21, 2.569961e-21, 1.28498e-20, 
    7.709882e-21, -2.569961e-21, 0, -2.569961e-21, -7.709882e-21, 
    1.541976e-20, 7.709882e-21, -7.709882e-21, 1.798972e-20, 0, 
    -2.569961e-21, 2.569961e-21, 1.003089e-36, 5.139921e-21, 1.027984e-20, 
    -1.027984e-20, 1.027984e-20, -2.569961e-21, 2.569961e-21, 1.027984e-20, 
    -1.027984e-20, -2.569961e-21, 1.28498e-20, 5.139921e-21, -1.541976e-20, 
    -5.139921e-21, 1.027984e-20, -2.569961e-21, 0, -1.003089e-36, 
    -1.541976e-20, -7.709882e-21, 2.569961e-21, 2.569961e-21, 1.28498e-20, 
    7.709882e-21, 7.709882e-21, 7.709882e-21, -2.569961e-21, 1.027984e-20, 
    1.28498e-20, 2.569961e-21, 0, 2.569961e-21, -2.569961e-21, 7.709882e-21, 
    5.139921e-21, -5.139921e-21, 1.28498e-20, 7.709882e-21, 1.28498e-20, 
    7.709882e-21, 0, -2.569961e-21, 1.027984e-20, 7.709882e-21, 0, 
    -1.28498e-20, -2.569961e-21, -1.003089e-36, -7.709882e-21, 2.569961e-21, 
    5.139921e-21, 1.027984e-20, 2.569961e-21, -1.003089e-36, 1.28498e-20, 
    -5.139921e-21, -1.541976e-20, -1.28498e-20, 0, 2.569961e-21, 
    7.709882e-21, -5.139921e-21, 0, -2.569961e-21, 1.541976e-20, 
    -7.709882e-21, 1.798972e-20, -7.709882e-21, -5.139921e-21, 1.027984e-20, 
    5.139921e-21, -5.139921e-21, -2.569961e-21, -2.569961e-21, -5.139921e-21, 
    1.027984e-20, 1.027984e-20, -7.709882e-21, 2.569961e-21, 7.709882e-21, 
    2.569961e-21, 5.139921e-21, 5.139921e-21, -1.003089e-36, 5.139921e-21, 
    7.709882e-21, -5.139921e-21, -2.569961e-21, 2.569961e-21, -7.709882e-21, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, -1.003089e-36, 5.139921e-21, 
    -5.139921e-21, 0, 5.139921e-21, -7.709882e-21, 7.709882e-21, 
    5.139921e-21, 1.541976e-20, 5.139921e-21, -2.569961e-21, -1.28498e-20, 
    -1.027984e-20, -1.027984e-20, 2.569961e-21, 2.055969e-20, 7.709882e-21, 
    -7.709882e-21, -7.709882e-21, -5.139921e-21, -2.569961e-21, 2.569961e-21, 
    1.003089e-36, 0, 5.139921e-21, 5.139921e-21, -7.709882e-21, 
    -2.569961e-21, 1.003089e-36, -1.541976e-20, -7.709882e-21, 7.709882e-21, 
    0, 1.541976e-20, -1.541976e-20, 7.709882e-21, 5.139921e-21, 5.139921e-21, 
    1.28498e-20, 5.139921e-21, 0, -1.541976e-20, -7.709882e-21, 5.139921e-21, 
    -2.055969e-20, 2.569961e-21, 5.139921e-21, 7.709882e-21, 5.139921e-21, 
    -5.139921e-21, -1.027984e-20, -2.569961e-21, 2.569961e-21, 2.569961e-21, 
    2.569961e-21, -7.709882e-21, -2.569961e-21, -1.541976e-20,
  -5.139921e-21, 2.569961e-21, -1.541976e-20, -5.139921e-21, 0, -1.28498e-20, 
    -1.003089e-36, -7.709882e-21, -1.28498e-20, -3.340949e-20, -2.569961e-21, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, -1.28498e-20, -2.569961e-21, 
    7.709882e-21, -1.28498e-20, 2.569961e-21, -7.709882e-21, 2.569961e-21, 
    -5.139921e-21, -5.139921e-21, 7.709882e-21, 1.28498e-20, -1.798972e-20, 
    -1.027984e-20, 1.027984e-20, 7.709882e-21, -2.569961e-21, 1.027984e-20, 
    -1.003089e-36, 2.569961e-21, 7.709882e-21, -2.569961e-21, -1.798972e-20, 
    -7.709882e-21, 5.139921e-21, 2.569961e-21, 5.139921e-21, -5.139921e-21, 
    -1.003089e-36, -7.709882e-21, 2.569961e-21, -1.28498e-20, -1.003089e-36, 
    -5.139921e-21, 0, -5.139921e-21, -1.027984e-20, -7.709882e-21, 
    -1.541976e-20, 7.709882e-21, -5.139921e-21, -5.139921e-21, -2.569961e-21, 
    -2.569961e-21, 2.569961e-21, 1.541976e-20, -2.569961e-21, 5.139921e-21, 
    7.709882e-21, 5.139921e-21, 1.28498e-20, -3.009266e-36, 1.003089e-36, 
    -2.055969e-20, -1.541976e-20, -5.139921e-21, 1.541976e-20, -5.139921e-21, 
    1.541976e-20, -5.139921e-21, 1.541976e-20, 5.139921e-21, 1.28498e-20, 
    1.003089e-36, 5.139921e-21, -2.569961e-21, -2.569961e-21, 1.541976e-20, 
    -1.027984e-20, 1.027984e-20, 2.055969e-20, -5.139921e-21, -1.541976e-20, 
    1.28498e-20, 1.027984e-20, 7.709882e-21, -2.569961e-21, 2.569961e-21, 
    -2.312965e-20, 2.055969e-20, -7.709882e-21, 7.709882e-21, 1.28498e-20, 
    1.003089e-36, -5.139921e-21, 2.569961e-21, -2.312965e-20, 1.003089e-36, 
    2.569961e-21, -7.709882e-21, 5.139921e-21, -2.569961e-21, -5.139921e-21, 
    -5.139921e-21, -2.569961e-21, -1.003089e-36, -5.139921e-21, 
    -2.312965e-20, -5.139921e-21, -7.709882e-21, -1.027984e-20, 2.569961e-21, 
    1.003089e-36, -1.027984e-20, 1.027984e-20, 1.003089e-36, 2.569961e-21, 
    7.709882e-21, 7.709882e-21, 0, -2.569961e-21, -2.569961e-21, 
    1.541976e-20, -5.139921e-21, -5.139921e-21, -7.709882e-21, -1.003089e-36, 
    -1.027984e-20, -1.027984e-20, -1.798972e-20, 5.139921e-21, -5.139921e-21, 
    7.709882e-21, 7.709882e-21, 7.709882e-21, 2.569961e-21, 7.709882e-21, 
    5.139921e-21, -1.541976e-20, 2.055969e-20, -2.569961e-21, -5.139921e-21, 
    1.541976e-20, -2.055969e-20, -7.709882e-21, -1.28498e-20, 1.003089e-36, 
    2.569961e-21, -1.28498e-20, 2.569961e-21, 1.28498e-20, -5.139921e-21, 
    -2.569961e-21, -7.709882e-21, 1.027984e-20, 2.569961e-21, -7.709882e-21, 
    0, -7.709882e-21, -2.569961e-21, -7.709882e-21, 7.709882e-21, 0, 
    -1.541976e-20, 1.027984e-20, -5.139921e-21, -1.28498e-20, 1.027984e-20, 
    -2.569961e-21, -7.709882e-21, 1.798972e-20, -7.709882e-21, -1.027984e-20, 
    1.541976e-20, -1.003089e-36, 7.709882e-21, 2.569961e-21, -1.027984e-20, 
    0, 1.28498e-20, -1.027984e-20, 2.569961e-21, -7.709882e-21, 0, 0, 
    -1.28498e-20, -7.709882e-21, 1.027984e-20, 5.139921e-21, 7.709882e-21, 
    2.569961e-21, -5.139921e-21, 1.798972e-20, -1.003089e-36, -5.139921e-21, 
    -2.569961e-21, 0, -1.027984e-20, -5.139921e-21, 5.139921e-21, 
    7.709882e-21, 1.798972e-20, 5.139921e-21, -2.569961e-21, -1.027984e-20, 
    -7.709882e-21, -5.139921e-21, 1.28498e-20, -5.139921e-21, 2.312965e-20, 
    -2.569961e-21, 1.027984e-20, 1.28498e-20, -1.027984e-20, -1.003089e-36, 
    2.569961e-21, 0, 5.139921e-21, -1.541976e-20, 2.569961e-21, 0, 
    7.709882e-21, -1.798972e-20, 0, -1.003089e-36, -2.569961e-21, 
    -2.569961e-21, 7.709882e-21, 1.027984e-20, -7.709882e-21, 5.139921e-21, 
    1.541976e-20, 1.541976e-20, 0, 1.541976e-20, -2.569961e-21, 1.003089e-36, 
    -1.798972e-20, 1.798972e-20, -2.569961e-21, -1.027984e-20, -5.139921e-21, 
    1.003089e-36, 1.28498e-20, -1.541976e-20, -1.003089e-36, -1.027984e-20, 
    -2.569961e-21, 5.139921e-21, 7.709882e-21, -1.027984e-20, 7.709882e-21, 
    1.28498e-20, 1.28498e-20, -1.28498e-20, -5.139921e-21, -2.569961e-21, 
    1.541976e-20, -2.569961e-21, 1.541976e-20, -5.139921e-21, -7.709882e-21, 
    -2.569961e-21, 5.139921e-21, 1.798972e-20, 2.312965e-20, -2.826957e-20, 
    -7.709882e-21, 7.709882e-21, 1.541976e-20, 1.541976e-20, 5.139921e-21, 
    -1.798972e-20, 1.027984e-20, -1.003089e-36, -1.28498e-20, 0, 
    -5.139921e-21, -1.003089e-36, 7.709882e-21, 1.003089e-36, 1.798972e-20, 
    -1.027984e-20, 1.003089e-36, -5.139921e-21, 7.709882e-21, 2.569961e-21, 
    1.28498e-20, 2.569961e-21, 5.139921e-21, 5.139921e-21, 1.027984e-20, 
    7.709882e-21, 7.709882e-21, 7.709882e-21, 2.569961e-21, 0, 1.003089e-36, 
    1.541976e-20, -7.709882e-21, -1.28498e-20, -1.541976e-20, -1.541976e-20, 
    -2.569961e-21, -1.28498e-20, -1.28498e-20, 1.003089e-36, -1.027984e-20, 
    -5.139921e-21, -5.139921e-21, 0, 2.569961e-21, 5.139921e-21, 
    -1.027984e-20, 1.027984e-20, -1.28498e-20, 2.569961e-21, 1.003089e-36, 
    2.569961e-21, -7.709882e-21, 1.798972e-20, 7.709882e-21, -5.139921e-21, 
    -2.055969e-20, -7.709882e-21, -1.541976e-20, 1.28498e-20, 7.709882e-21, 
    -1.027984e-20, 1.798972e-20, -1.798972e-20, 0, -5.139921e-21, 
    -1.027984e-20, 2.569961e-21,
  1.28498e-20, 2.569961e-21, 2.569961e-21, -1.28498e-20, 0, 7.709882e-21, 
    -7.709882e-21, -2.569961e-21, -1.003089e-36, 2.569961e-21, -1.28498e-20, 
    7.709882e-21, -5.139921e-21, 1.003089e-36, 2.569961e-21, -1.541976e-20, 
    1.28498e-20, 2.569961e-21, 2.569961e-21, 7.709882e-21, 1.003089e-36, 
    1.28498e-20, -5.139921e-21, -1.541976e-20, 7.709882e-21, -5.139921e-21, 
    -5.139921e-21, -2.569961e-21, -1.28498e-20, -1.027984e-20, 2.569961e-21, 
    1.28498e-20, -5.139921e-21, 2.569961e-21, -1.798972e-20, -5.139921e-21, 
    -2.569961e-21, -1.027984e-20, 0, 2.055969e-20, -1.798972e-20, 
    5.139921e-21, 0, 2.569961e-21, 7.709882e-21, -2.055969e-20, 2.569961e-21, 
    -1.003089e-36, 2.569961e-21, 2.569961e-21, -1.027984e-20, 1.003089e-36, 
    -2.569961e-21, 5.139921e-21, -5.139921e-21, -1.027984e-20, 7.709882e-21, 
    -5.139921e-21, 1.541976e-20, -1.027984e-20, 1.28498e-20, -2.569961e-21, 
    -5.139921e-21, -1.798972e-20, 1.003089e-36, -1.027984e-20, -5.139921e-21, 
    1.28498e-20, 4.625929e-20, -2.569961e-21, 1.541976e-20, -1.003089e-36, 
    7.709882e-21, 5.139921e-21, -5.139921e-21, -7.709882e-21, 1.027984e-20, 
    0, -2.569961e-21, 5.139921e-21, -2.569961e-21, 1.28498e-20, 5.139921e-21, 
    -2.055969e-20, -1.541976e-20, 2.055969e-20, -7.709882e-21, -2.312965e-20, 
    5.015443e-37, 5.139921e-21, 0, 5.139921e-21, 1.541976e-20, 2.569961e-21, 
    1.541976e-20, -2.569961e-21, -5.139921e-21, 1.003089e-36, 1.798972e-20, 
    -5.139921e-21, -5.139921e-21, 7.709882e-21, -5.139921e-21, -2.569961e-21, 
    -5.139921e-21, 2.569961e-21, 1.027984e-20, -1.28498e-20, 1.027984e-20, 
    1.28498e-20, 1.28498e-20, 5.139921e-21, -1.798972e-20, -2.569961e-21, 
    2.569961e-21, 1.003089e-36, 2.569961e-21, -5.139921e-21, -7.709882e-21, 
    5.139921e-21, 1.003089e-36, -1.28498e-20, -1.28498e-20, -1.027984e-20, 
    1.027984e-20, -5.139921e-21, 2.569961e-20, 2.569961e-21, 1.541976e-20, 
    5.139921e-21, 0, -1.28498e-20, -1.541976e-20, 7.709882e-21, 
    -7.709882e-21, -1.027984e-20, -5.139921e-21, 1.541976e-20, -1.027984e-20, 
    -2.569961e-21, -2.569961e-21, -2.569961e-20, 7.709882e-21, -2.312965e-20, 
    1.28498e-20, -7.709882e-21, -1.28498e-20, 2.569961e-21, 0, 1.798972e-20, 
    1.027984e-20, -1.003089e-36, 1.28498e-20, -5.139921e-21, -1.28498e-20, 
    1.798972e-20, -2.569961e-21, 2.312965e-20, 5.139921e-21, -1.798972e-20, 
    2.569961e-21, -1.28498e-20, -2.569961e-21, -5.139921e-21, 1.28498e-20, 
    1.027984e-20, 5.139921e-21, 5.139921e-21, 2.569961e-21, -1.003089e-36, 
    -1.798972e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, 0, 
    2.569961e-21, -5.139921e-21, -1.003089e-36, 0, 1.28498e-20, 0, 
    2.569961e-21, -2.569961e-21, -2.569961e-21, 1.027984e-20, 5.139921e-21, 
    5.139921e-21, 1.541976e-20, -7.709882e-21, 7.709882e-21, 2.569961e-21, 
    2.569961e-21, 2.569961e-21, -2.569961e-20, -7.709882e-21, 5.139921e-21, 
    1.541976e-20, -5.139921e-21, -5.139921e-21, -1.798972e-20, -5.139921e-21, 
    2.569961e-21, -7.709882e-21, 1.28498e-20, 7.709882e-21, -2.569961e-21, 
    -5.139921e-21, -7.709882e-21, -2.569961e-21, 5.139921e-21, -3.597945e-20, 
    1.027984e-20, -1.28498e-20, -7.709882e-21, 1.027984e-20, 1.027984e-20, 
    1.28498e-20, 5.139921e-21, 1.003089e-36, 7.709882e-21, -1.003089e-36, 
    1.798972e-20, 1.003089e-36, -5.139921e-21, 1.798972e-20, 1.027984e-20, 
    1.027984e-20, -2.569961e-21, 1.541976e-20, -7.709882e-21, -1.027984e-20, 
    -5.139921e-21, -7.709882e-21, 1.798972e-20, -1.027984e-20, -5.139921e-21, 
    5.139921e-21, 2.569961e-21, 7.709882e-21, 7.709882e-21, -1.027984e-20, 
    1.28498e-20, 5.139921e-21, 7.709882e-21, -5.139921e-21, 7.709882e-21, 
    -2.569961e-21, -1.027984e-20, -2.569961e-21, 1.003089e-36, 2.569961e-20, 
    1.28498e-20, -7.709882e-21, 1.027984e-20, 1.003089e-36, 5.139921e-21, 
    -5.139921e-21, 1.798972e-20, -7.709882e-21, -5.139921e-21, 2.569961e-21, 
    2.055969e-20, -2.569961e-21, -2.569961e-21, 7.709882e-21, -1.28498e-20, 
    2.569961e-20, 1.798972e-20, 1.003089e-36, -1.541976e-20, -2.569961e-21, 
    -1.027984e-20, -1.003089e-36, 1.798972e-20, 2.055969e-20, -5.139921e-21, 
    2.569961e-21, 0, 7.709882e-21, -5.139921e-21, -1.798972e-20, 
    -1.027984e-20, -2.569961e-21, 5.139921e-21, 1.027984e-20, 7.709882e-21, 
    -1.798972e-20, 7.709882e-21, 7.709882e-21, 2.055969e-20, -1.541976e-20, 
    -1.003089e-36, 7.709882e-21, -2.055969e-20, 7.709882e-21, -1.027984e-20, 
    -2.569961e-21, -7.709882e-21, 7.709882e-21, -2.569961e-21, -1.541976e-20, 
    -2.569961e-21, 5.139921e-21, 7.709882e-21, 1.027984e-20, 1.027984e-20, 
    2.569961e-21, 5.139921e-21, 1.28498e-20, 7.709882e-21, -7.709882e-21, 
    -1.798972e-20, 1.541976e-20, 2.312965e-20, 1.28498e-20, 7.709882e-21, 
    -1.003089e-36, 2.569961e-21, -1.541976e-20, -1.003089e-36, 1.541976e-20, 
    -5.139921e-21, -1.798972e-20, 0, -1.28498e-20, 2.569961e-21, 
    -5.139921e-21, -1.003089e-36, 2.055969e-20, -7.709882e-21, -5.139921e-21, 
    5.139921e-21, 5.139921e-21, 2.569961e-21, -1.541976e-20, -1.541976e-20, 
    -1.541976e-20, -2.569961e-21,
  6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N_TO_SOIL1N =
  5.289164e-12, 5.312433e-12, 5.307909e-12, 5.326677e-12, 5.316266e-12, 
    5.328556e-12, 5.293882e-12, 5.313357e-12, 5.300924e-12, 5.291259e-12, 
    5.3631e-12, 5.327515e-12, 5.400061e-12, 5.377367e-12, 5.434374e-12, 
    5.39653e-12, 5.442005e-12, 5.433282e-12, 5.459535e-12, 5.452013e-12, 
    5.485594e-12, 5.463006e-12, 5.503e-12, 5.480199e-12, 5.483766e-12, 
    5.462261e-12, 5.334675e-12, 5.35867e-12, 5.333254e-12, 5.336676e-12, 
    5.33514e-12, 5.316482e-12, 5.307079e-12, 5.287386e-12, 5.29096e-12, 
    5.305425e-12, 5.338214e-12, 5.327083e-12, 5.355134e-12, 5.354501e-12, 
    5.38573e-12, 5.37165e-12, 5.424137e-12, 5.40922e-12, 5.452327e-12, 
    5.441486e-12, 5.451818e-12, 5.448685e-12, 5.451859e-12, 5.435959e-12, 
    5.442772e-12, 5.428781e-12, 5.374287e-12, 5.390303e-12, 5.342536e-12, 
    5.313814e-12, 5.294736e-12, 5.281198e-12, 5.283112e-12, 5.28676e-12, 
    5.30551e-12, 5.323137e-12, 5.33657e-12, 5.345556e-12, 5.35441e-12, 
    5.381211e-12, 5.395395e-12, 5.427154e-12, 5.421422e-12, 5.431132e-12, 
    5.440408e-12, 5.455982e-12, 5.453418e-12, 5.460279e-12, 5.430876e-12, 
    5.450418e-12, 5.418157e-12, 5.426981e-12, 5.356819e-12, 5.330086e-12, 
    5.318725e-12, 5.308779e-12, 5.284583e-12, 5.301292e-12, 5.294706e-12, 
    5.310376e-12, 5.320333e-12, 5.315408e-12, 5.345802e-12, 5.333986e-12, 
    5.396236e-12, 5.369423e-12, 5.439326e-12, 5.422599e-12, 5.443335e-12, 
    5.432754e-12, 5.450885e-12, 5.434567e-12, 5.462833e-12, 5.468988e-12, 
    5.464782e-12, 5.480939e-12, 5.433662e-12, 5.451819e-12, 5.31527e-12, 
    5.316074e-12, 5.319815e-12, 5.303368e-12, 5.302361e-12, 5.287288e-12, 
    5.3007e-12, 5.306412e-12, 5.32091e-12, 5.329486e-12, 5.337639e-12, 
    5.355563e-12, 5.375582e-12, 5.403574e-12, 5.423683e-12, 5.437163e-12, 
    5.428897e-12, 5.436194e-12, 5.428037e-12, 5.424213e-12, 5.466682e-12, 
    5.442835e-12, 5.478615e-12, 5.476635e-12, 5.460443e-12, 5.476858e-12, 
    5.316637e-12, 5.312016e-12, 5.295969e-12, 5.308527e-12, 5.285646e-12, 
    5.298454e-12, 5.305818e-12, 5.334233e-12, 5.340475e-12, 5.346265e-12, 
    5.357698e-12, 5.372371e-12, 5.398109e-12, 5.420504e-12, 5.440947e-12, 
    5.43945e-12, 5.439977e-12, 5.444544e-12, 5.433231e-12, 5.446401e-12, 
    5.448612e-12, 5.442832e-12, 5.47637e-12, 5.466788e-12, 5.476593e-12, 
    5.470354e-12, 5.313518e-12, 5.321295e-12, 5.317093e-12, 5.324995e-12, 
    5.319428e-12, 5.344184e-12, 5.351606e-12, 5.386335e-12, 5.372082e-12, 
    5.394765e-12, 5.374386e-12, 5.377997e-12, 5.395507e-12, 5.375487e-12, 
    5.41927e-12, 5.389588e-12, 5.444721e-12, 5.415082e-12, 5.446579e-12, 
    5.440859e-12, 5.450329e-12, 5.458811e-12, 5.469481e-12, 5.489169e-12, 
    5.48461e-12, 5.501075e-12, 5.332889e-12, 5.342976e-12, 5.342088e-12, 
    5.352644e-12, 5.360451e-12, 5.377372e-12, 5.404511e-12, 5.394305e-12, 
    5.41304e-12, 5.416802e-12, 5.388338e-12, 5.405815e-12, 5.349727e-12, 
    5.35879e-12, 5.353394e-12, 5.333685e-12, 5.396658e-12, 5.36434e-12, 
    5.424015e-12, 5.406509e-12, 5.457602e-12, 5.432192e-12, 5.4821e-12, 
    5.503437e-12, 5.523515e-12, 5.546982e-12, 5.348481e-12, 5.341627e-12, 
    5.3539e-12, 5.37088e-12, 5.386633e-12, 5.407577e-12, 5.409719e-12, 
    5.413643e-12, 5.423806e-12, 5.43235e-12, 5.414884e-12, 5.434493e-12, 
    5.360892e-12, 5.399463e-12, 5.339036e-12, 5.357233e-12, 5.369879e-12, 
    5.364331e-12, 5.393139e-12, 5.399929e-12, 5.42752e-12, 5.413257e-12, 
    5.498171e-12, 5.460603e-12, 5.564848e-12, 5.535717e-12, 5.339233e-12, 
    5.348457e-12, 5.380564e-12, 5.365288e-12, 5.408974e-12, 5.419728e-12, 
    5.428469e-12, 5.439644e-12, 5.44085e-12, 5.447471e-12, 5.436621e-12, 
    5.447042e-12, 5.407621e-12, 5.425237e-12, 5.376894e-12, 5.388661e-12, 
    5.383248e-12, 5.37731e-12, 5.395635e-12, 5.415159e-12, 5.415576e-12, 
    5.421836e-12, 5.439478e-12, 5.409151e-12, 5.503022e-12, 5.445051e-12, 
    5.358517e-12, 5.376287e-12, 5.378824e-12, 5.371941e-12, 5.418649e-12, 
    5.401726e-12, 5.447309e-12, 5.434989e-12, 5.455175e-12, 5.445144e-12, 
    5.443669e-12, 5.430786e-12, 5.422765e-12, 5.402502e-12, 5.386014e-12, 
    5.372939e-12, 5.375979e-12, 5.390342e-12, 5.416353e-12, 5.440959e-12, 
    5.435569e-12, 5.453641e-12, 5.405807e-12, 5.425865e-12, 5.418113e-12, 
    5.438326e-12, 5.394034e-12, 5.431754e-12, 5.384393e-12, 5.388546e-12, 
    5.401389e-12, 5.427226e-12, 5.432941e-12, 5.439044e-12, 5.435278e-12, 
    5.417013e-12, 5.41402e-12, 5.401077e-12, 5.397504e-12, 5.387641e-12, 
    5.379476e-12, 5.386937e-12, 5.394771e-12, 5.417021e-12, 5.437071e-12, 
    5.458932e-12, 5.464281e-12, 5.489825e-12, 5.469032e-12, 5.503345e-12, 
    5.474174e-12, 5.524669e-12, 5.433938e-12, 5.473315e-12, 5.401974e-12, 
    5.409659e-12, 5.423561e-12, 5.455445e-12, 5.438231e-12, 5.458362e-12, 
    5.413903e-12, 5.390838e-12, 5.384869e-12, 5.373734e-12, 5.385123e-12, 
    5.384197e-12, 5.395095e-12, 5.391593e-12, 5.417759e-12, 5.403704e-12, 
    5.443632e-12, 5.458202e-12, 5.49935e-12, 5.524575e-12, 5.55025e-12, 
    5.561586e-12, 5.565036e-12, 5.566479e-12 ;

 SOIL3N_vr =
  1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819,
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.81819, 1.81819, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.81819, 1.81819, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.81819, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819,
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 
    1.818187, 1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818187, 1.818188, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818188, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3_HR =
  3.199944e-11, 3.214022e-11, 3.211285e-11, 3.22264e-11, 3.216341e-11, 
    3.223776e-11, 3.202798e-11, 3.214581e-11, 3.207059e-11, 3.201212e-11, 
    3.244676e-11, 3.223146e-11, 3.267037e-11, 3.253307e-11, 3.287796e-11, 
    3.264901e-11, 3.292413e-11, 3.287135e-11, 3.303018e-11, 3.298468e-11, 
    3.318784e-11, 3.305118e-11, 3.329315e-11, 3.31552e-11, 3.317678e-11, 
    3.304668e-11, 3.227479e-11, 3.241996e-11, 3.226619e-11, 3.228689e-11, 
    3.22776e-11, 3.216471e-11, 3.210783e-11, 3.198868e-11, 3.201031e-11, 
    3.209782e-11, 3.22962e-11, 3.222886e-11, 3.239856e-11, 3.239473e-11, 
    3.258367e-11, 3.249848e-11, 3.281603e-11, 3.272578e-11, 3.298658e-11, 
    3.292099e-11, 3.29835e-11, 3.296455e-11, 3.298375e-11, 3.288755e-11, 
    3.292877e-11, 3.284412e-11, 3.251444e-11, 3.261133e-11, 3.232234e-11, 
    3.214858e-11, 3.203315e-11, 3.195125e-11, 3.196282e-11, 3.19849e-11, 
    3.209833e-11, 3.220498e-11, 3.228625e-11, 3.234061e-11, 3.239418e-11, 
    3.255633e-11, 3.264214e-11, 3.283428e-11, 3.27996e-11, 3.285835e-11, 
    3.291447e-11, 3.300869e-11, 3.299318e-11, 3.303469e-11, 3.28568e-11, 
    3.297503e-11, 3.277985e-11, 3.283323e-11, 3.240876e-11, 3.224702e-11, 
    3.217829e-11, 3.211811e-11, 3.197173e-11, 3.207282e-11, 3.203297e-11, 
    3.212777e-11, 3.218802e-11, 3.215822e-11, 3.23421e-11, 3.227061e-11, 
    3.264723e-11, 3.248501e-11, 3.290792e-11, 3.280672e-11, 3.293218e-11, 
    3.286816e-11, 3.297785e-11, 3.287913e-11, 3.305014e-11, 3.308738e-11, 
    3.306193e-11, 3.315968e-11, 3.287366e-11, 3.29835e-11, 3.215738e-11, 
    3.216225e-11, 3.218488e-11, 3.208537e-11, 3.207928e-11, 3.198809e-11, 
    3.206923e-11, 3.210379e-11, 3.219151e-11, 3.224339e-11, 3.229271e-11, 
    3.240116e-11, 3.252227e-11, 3.269162e-11, 3.281328e-11, 3.289484e-11, 
    3.284483e-11, 3.288898e-11, 3.283962e-11, 3.281649e-11, 3.307343e-11, 
    3.292915e-11, 3.314562e-11, 3.313364e-11, 3.303568e-11, 3.313499e-11, 
    3.216566e-11, 3.213769e-11, 3.204061e-11, 3.211659e-11, 3.197816e-11, 
    3.205565e-11, 3.21002e-11, 3.227211e-11, 3.230988e-11, 3.23449e-11, 
    3.241407e-11, 3.250284e-11, 3.265856e-11, 3.279405e-11, 3.291773e-11, 
    3.290867e-11, 3.291186e-11, 3.293949e-11, 3.287105e-11, 3.295073e-11, 
    3.29641e-11, 3.292914e-11, 3.313204e-11, 3.307407e-11, 3.313338e-11, 
    3.309564e-11, 3.214678e-11, 3.219383e-11, 3.216841e-11, 3.221622e-11, 
    3.218254e-11, 3.233231e-11, 3.237722e-11, 3.258733e-11, 3.25011e-11, 
    3.263833e-11, 3.251503e-11, 3.253688e-11, 3.264282e-11, 3.25217e-11, 
    3.278658e-11, 3.2607e-11, 3.294056e-11, 3.276125e-11, 3.29518e-11, 
    3.29172e-11, 3.297449e-11, 3.30258e-11, 3.309036e-11, 3.320948e-11, 
    3.318189e-11, 3.328151e-11, 3.226398e-11, 3.232501e-11, 3.231963e-11, 
    3.23835e-11, 3.243073e-11, 3.25331e-11, 3.269729e-11, 3.263555e-11, 
    3.274889e-11, 3.277165e-11, 3.259945e-11, 3.270518e-11, 3.236585e-11, 
    3.242068e-11, 3.238803e-11, 3.22688e-11, 3.264978e-11, 3.245426e-11, 
    3.281529e-11, 3.270938e-11, 3.301849e-11, 3.286477e-11, 3.316671e-11, 
    3.329579e-11, 3.341727e-11, 3.355924e-11, 3.235831e-11, 3.231684e-11, 
    3.239109e-11, 3.249382e-11, 3.258913e-11, 3.271584e-11, 3.27288e-11, 
    3.275254e-11, 3.281402e-11, 3.286572e-11, 3.276005e-11, 3.287868e-11, 
    3.24334e-11, 3.266675e-11, 3.230117e-11, 3.241126e-11, 3.248777e-11, 
    3.24542e-11, 3.262849e-11, 3.266957e-11, 3.283649e-11, 3.27502e-11, 
    3.326394e-11, 3.303665e-11, 3.366733e-11, 3.349109e-11, 3.230236e-11, 
    3.235817e-11, 3.255242e-11, 3.245999e-11, 3.27243e-11, 3.278935e-11, 
    3.284224e-11, 3.290984e-11, 3.291714e-11, 3.29572e-11, 3.289156e-11, 
    3.29546e-11, 3.271611e-11, 3.282269e-11, 3.253021e-11, 3.26014e-11, 
    3.256865e-11, 3.253273e-11, 3.264359e-11, 3.276171e-11, 3.276423e-11, 
    3.28021e-11, 3.290885e-11, 3.272536e-11, 3.329328e-11, 3.294256e-11, 
    3.241903e-11, 3.252654e-11, 3.254189e-11, 3.250024e-11, 3.278283e-11, 
    3.268044e-11, 3.295622e-11, 3.288169e-11, 3.300381e-11, 3.294312e-11, 
    3.29342e-11, 3.285625e-11, 3.280773e-11, 3.268514e-11, 3.258538e-11, 
    3.250628e-11, 3.252467e-11, 3.261157e-11, 3.276894e-11, 3.29178e-11, 
    3.288519e-11, 3.299453e-11, 3.270513e-11, 3.282648e-11, 3.277958e-11, 
    3.290187e-11, 3.263391e-11, 3.286211e-11, 3.257558e-11, 3.26007e-11, 
    3.267841e-11, 3.283472e-11, 3.286929e-11, 3.290622e-11, 3.288343e-11, 
    3.277293e-11, 3.275482e-11, 3.267652e-11, 3.26549e-11, 3.259523e-11, 
    3.254583e-11, 3.259096e-11, 3.263837e-11, 3.277297e-11, 3.289428e-11, 
    3.302654e-11, 3.30589e-11, 3.321344e-11, 3.308764e-11, 3.329523e-11, 
    3.311875e-11, 3.342425e-11, 3.287533e-11, 3.311355e-11, 3.268194e-11, 
    3.272844e-11, 3.281254e-11, 3.300544e-11, 3.29013e-11, 3.302309e-11, 
    3.275412e-11, 3.261457e-11, 3.257846e-11, 3.251109e-11, 3.257999e-11, 
    3.257439e-11, 3.264033e-11, 3.261914e-11, 3.277744e-11, 3.269241e-11, 
    3.293397e-11, 3.302213e-11, 3.327107e-11, 3.342368e-11, 3.357901e-11, 
    3.36476e-11, 3.366847e-11, 3.36772e-11 ;

 SOILC =
  17.34462, 17.3446, 17.34461, 17.3446, 17.3446, 17.34459, 17.34462, 17.3446, 
    17.34461, 17.34462, 17.34457, 17.3446, 17.34455, 17.34457, 17.34453, 
    17.34455, 17.34453, 17.34453, 17.34452, 17.34452, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.3445, 17.34452, 17.34459, 17.34458, 17.34459, 
    17.34459, 17.34459, 17.3446, 17.34461, 17.34462, 17.34462, 17.34461, 
    17.34459, 17.3446, 17.34458, 17.34458, 17.34456, 17.34457, 17.34454, 
    17.34455, 17.34452, 17.34453, 17.34452, 17.34452, 17.34452, 17.34453, 
    17.34453, 17.34454, 17.34457, 17.34456, 17.34459, 17.3446, 17.34462, 
    17.34462, 17.34462, 17.34462, 17.34461, 17.3446, 17.34459, 17.34459, 
    17.34458, 17.34456, 17.34455, 17.34454, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34452, 17.34453, 17.34452, 17.34454, 17.34454, 
    17.34458, 17.34459, 17.3446, 17.34461, 17.34462, 17.34461, 17.34462, 
    17.34461, 17.3446, 17.3446, 17.34459, 17.34459, 17.34455, 17.34457, 
    17.34453, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34451, 17.34451, 17.34451, 17.34453, 17.34452, 17.3446, 17.3446, 
    17.3446, 17.34461, 17.34461, 17.34462, 17.34461, 17.34461, 17.3446, 
    17.34459, 17.34459, 17.34458, 17.34457, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34454, 17.34454, 17.34451, 17.34453, 17.34451, 
    17.34451, 17.34452, 17.34451, 17.3446, 17.3446, 17.34461, 17.34461, 
    17.34462, 17.34461, 17.34461, 17.34459, 17.34459, 17.34459, 17.34458, 
    17.34457, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 17.34453, 
    17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 17.34451, 17.34451, 
    17.34451, 17.3446, 17.3446, 17.3446, 17.3446, 17.3446, 17.34459, 
    17.34458, 17.34456, 17.34457, 17.34456, 17.34457, 17.34457, 17.34455, 
    17.34457, 17.34454, 17.34456, 17.34453, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34451, 17.3445, 17.3445, 17.34449, 17.34459, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34457, 17.34455, 17.34456, 
    17.34455, 17.34454, 17.34456, 17.34455, 17.34458, 17.34458, 17.34458, 
    17.34459, 17.34455, 17.34457, 17.34454, 17.34455, 17.34452, 17.34453, 
    17.34451, 17.34449, 17.34448, 17.34447, 17.34458, 17.34459, 17.34458, 
    17.34457, 17.34456, 17.34455, 17.34455, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34458, 17.34455, 17.34459, 17.34458, 17.34457, 
    17.34457, 17.34456, 17.34455, 17.34454, 17.34455, 17.3445, 17.34452, 
    17.34446, 17.34447, 17.34459, 17.34458, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34455, 17.34454, 17.34457, 17.34456, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34454, 17.34453, 17.34455, 17.34449, 17.34453, 
    17.34458, 17.34457, 17.34457, 17.34457, 17.34454, 17.34455, 17.34452, 
    17.34453, 17.34452, 17.34453, 17.34453, 17.34453, 17.34454, 17.34455, 
    17.34456, 17.34457, 17.34457, 17.34456, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34455, 17.34454, 17.34454, 17.34453, 17.34456, 17.34453, 
    17.34456, 17.34456, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 
    17.34454, 17.34455, 17.34455, 17.34455, 17.34456, 17.34456, 17.34456, 
    17.34456, 17.34454, 17.34453, 17.34452, 17.34451, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.34448, 17.34453, 17.34451, 17.34455, 17.34455, 
    17.34454, 17.34452, 17.34453, 17.34452, 17.34455, 17.34456, 17.34456, 
    17.34457, 17.34456, 17.34456, 17.34456, 17.34456, 17.34454, 17.34455, 
    17.34453, 17.34452, 17.34449, 17.34448, 17.34446, 17.34446, 17.34446, 
    17.34445 ;

 SOILC_HR =
  6.358298e-08, 6.386256e-08, 6.380821e-08, 6.403371e-08, 6.390862e-08, 
    6.405628e-08, 6.363966e-08, 6.387366e-08, 6.372428e-08, 6.360815e-08, 
    6.447134e-08, 6.404377e-08, 6.491543e-08, 6.464276e-08, 6.532771e-08, 
    6.4873e-08, 6.541939e-08, 6.531458e-08, 6.563002e-08, 6.553965e-08, 
    6.594313e-08, 6.567172e-08, 6.615226e-08, 6.58783e-08, 6.592116e-08, 
    6.566277e-08, 6.412981e-08, 6.441811e-08, 6.411273e-08, 6.415384e-08, 
    6.413539e-08, 6.39112e-08, 6.379823e-08, 6.356161e-08, 6.360457e-08, 
    6.377836e-08, 6.417233e-08, 6.403859e-08, 6.437563e-08, 6.436802e-08, 
    6.474324e-08, 6.457406e-08, 6.520471e-08, 6.502547e-08, 6.554342e-08, 
    6.541316e-08, 6.553731e-08, 6.549966e-08, 6.55378e-08, 6.534675e-08, 
    6.542861e-08, 6.52605e-08, 6.460575e-08, 6.479818e-08, 6.422425e-08, 
    6.387916e-08, 6.364992e-08, 6.348726e-08, 6.351026e-08, 6.35541e-08, 
    6.377937e-08, 6.399117e-08, 6.415257e-08, 6.426054e-08, 6.436692e-08, 
    6.468895e-08, 6.485936e-08, 6.524096e-08, 6.517209e-08, 6.528876e-08, 
    6.540021e-08, 6.558732e-08, 6.555653e-08, 6.563896e-08, 6.528568e-08, 
    6.552047e-08, 6.513286e-08, 6.523888e-08, 6.439587e-08, 6.407466e-08, 
    6.393816e-08, 6.381866e-08, 6.352794e-08, 6.372871e-08, 6.364956e-08, 
    6.383784e-08, 6.395748e-08, 6.389831e-08, 6.42635e-08, 6.412152e-08, 
    6.486947e-08, 6.454731e-08, 6.53872e-08, 6.518622e-08, 6.543538e-08, 
    6.530824e-08, 6.552609e-08, 6.533003e-08, 6.566965e-08, 6.57436e-08, 
    6.569307e-08, 6.588719e-08, 6.531916e-08, 6.553731e-08, 6.389665e-08, 
    6.39063e-08, 6.395126e-08, 6.375364e-08, 6.374155e-08, 6.356043e-08, 
    6.372159e-08, 6.379021e-08, 6.396441e-08, 6.406746e-08, 6.416541e-08, 
    6.438078e-08, 6.462131e-08, 6.495763e-08, 6.519925e-08, 6.536121e-08, 
    6.52619e-08, 6.534958e-08, 6.525156e-08, 6.520562e-08, 6.571589e-08, 
    6.542937e-08, 6.585927e-08, 6.583548e-08, 6.564093e-08, 6.583816e-08, 
    6.391308e-08, 6.385754e-08, 6.366474e-08, 6.381563e-08, 6.35407e-08, 
    6.369459e-08, 6.378308e-08, 6.412449e-08, 6.41995e-08, 6.426905e-08, 
    6.440642e-08, 6.458272e-08, 6.489199e-08, 6.516106e-08, 6.540669e-08, 
    6.538869e-08, 6.539503e-08, 6.54499e-08, 6.531398e-08, 6.547221e-08, 
    6.549877e-08, 6.542933e-08, 6.58323e-08, 6.571717e-08, 6.583497e-08, 
    6.576001e-08, 6.38756e-08, 6.396904e-08, 6.391854e-08, 6.40135e-08, 
    6.394661e-08, 6.424406e-08, 6.433323e-08, 6.475051e-08, 6.457925e-08, 
    6.48518e-08, 6.460694e-08, 6.465033e-08, 6.486071e-08, 6.462017e-08, 
    6.514622e-08, 6.478959e-08, 6.545203e-08, 6.50959e-08, 6.547435e-08, 
    6.540562e-08, 6.551941e-08, 6.562132e-08, 6.574952e-08, 6.598609e-08, 
    6.59313e-08, 6.612913e-08, 6.410834e-08, 6.422955e-08, 6.421887e-08, 
    6.434571e-08, 6.443951e-08, 6.464282e-08, 6.496889e-08, 6.484628e-08, 
    6.507138e-08, 6.511657e-08, 6.477458e-08, 6.498456e-08, 6.431066e-08, 
    6.441955e-08, 6.435471e-08, 6.411791e-08, 6.487454e-08, 6.448624e-08, 
    6.520325e-08, 6.49929e-08, 6.560679e-08, 6.53015e-08, 6.590115e-08, 
    6.615751e-08, 6.639875e-08, 6.668071e-08, 6.429569e-08, 6.421333e-08, 
    6.436079e-08, 6.456481e-08, 6.475408e-08, 6.500573e-08, 6.503147e-08, 
    6.507862e-08, 6.520072e-08, 6.53034e-08, 6.509353e-08, 6.532913e-08, 
    6.444481e-08, 6.490824e-08, 6.41822e-08, 6.440084e-08, 6.455278e-08, 
    6.448612e-08, 6.483226e-08, 6.491384e-08, 6.524535e-08, 6.507398e-08, 
    6.609424e-08, 6.564286e-08, 6.689538e-08, 6.654536e-08, 6.418456e-08, 
    6.429541e-08, 6.468117e-08, 6.449763e-08, 6.502253e-08, 6.515172e-08, 
    6.525676e-08, 6.539102e-08, 6.540552e-08, 6.548507e-08, 6.53547e-08, 
    6.547992e-08, 6.500627e-08, 6.521793e-08, 6.463707e-08, 6.477845e-08, 
    6.471341e-08, 6.464207e-08, 6.486225e-08, 6.509683e-08, 6.510184e-08, 
    6.517705e-08, 6.538904e-08, 6.502465e-08, 6.615252e-08, 6.545599e-08, 
    6.441627e-08, 6.462978e-08, 6.466026e-08, 6.457756e-08, 6.513877e-08, 
    6.493543e-08, 6.548313e-08, 6.53351e-08, 6.557763e-08, 6.545712e-08, 
    6.543939e-08, 6.52846e-08, 6.518822e-08, 6.494476e-08, 6.474665e-08, 
    6.458955e-08, 6.462608e-08, 6.479865e-08, 6.511118e-08, 6.540683e-08, 
    6.534207e-08, 6.55592e-08, 6.498447e-08, 6.522547e-08, 6.513232e-08, 
    6.537519e-08, 6.484301e-08, 6.529623e-08, 6.472717e-08, 6.477707e-08, 
    6.493139e-08, 6.524182e-08, 6.531049e-08, 6.538382e-08, 6.533857e-08, 
    6.511911e-08, 6.508316e-08, 6.492764e-08, 6.488471e-08, 6.47662e-08, 
    6.46681e-08, 6.475774e-08, 6.485187e-08, 6.51192e-08, 6.536012e-08, 
    6.562277e-08, 6.568705e-08, 6.599396e-08, 6.574413e-08, 6.61564e-08, 
    6.580591e-08, 6.641262e-08, 6.532247e-08, 6.579559e-08, 6.493841e-08, 
    6.503075e-08, 6.519779e-08, 6.558088e-08, 6.537405e-08, 6.561592e-08, 
    6.508175e-08, 6.480461e-08, 6.473289e-08, 6.459911e-08, 6.473595e-08, 
    6.472482e-08, 6.485576e-08, 6.481368e-08, 6.512808e-08, 6.49592e-08, 
    6.543894e-08, 6.561401e-08, 6.610841e-08, 6.641149e-08, 6.671998e-08, 
    6.685619e-08, 6.689764e-08, 6.691497e-08 ;

 SOILC_LOSS =
  6.358298e-08, 6.386256e-08, 6.380821e-08, 6.403371e-08, 6.390862e-08, 
    6.405628e-08, 6.363966e-08, 6.387366e-08, 6.372428e-08, 6.360815e-08, 
    6.447134e-08, 6.404377e-08, 6.491543e-08, 6.464276e-08, 6.532771e-08, 
    6.4873e-08, 6.541939e-08, 6.531458e-08, 6.563002e-08, 6.553965e-08, 
    6.594313e-08, 6.567172e-08, 6.615226e-08, 6.58783e-08, 6.592116e-08, 
    6.566277e-08, 6.412981e-08, 6.441811e-08, 6.411273e-08, 6.415384e-08, 
    6.413539e-08, 6.39112e-08, 6.379823e-08, 6.356161e-08, 6.360457e-08, 
    6.377836e-08, 6.417233e-08, 6.403859e-08, 6.437563e-08, 6.436802e-08, 
    6.474324e-08, 6.457406e-08, 6.520471e-08, 6.502547e-08, 6.554342e-08, 
    6.541316e-08, 6.553731e-08, 6.549966e-08, 6.55378e-08, 6.534675e-08, 
    6.542861e-08, 6.52605e-08, 6.460575e-08, 6.479818e-08, 6.422425e-08, 
    6.387916e-08, 6.364992e-08, 6.348726e-08, 6.351026e-08, 6.35541e-08, 
    6.377937e-08, 6.399117e-08, 6.415257e-08, 6.426054e-08, 6.436692e-08, 
    6.468895e-08, 6.485936e-08, 6.524096e-08, 6.517209e-08, 6.528876e-08, 
    6.540021e-08, 6.558732e-08, 6.555653e-08, 6.563896e-08, 6.528568e-08, 
    6.552047e-08, 6.513286e-08, 6.523888e-08, 6.439587e-08, 6.407466e-08, 
    6.393816e-08, 6.381866e-08, 6.352794e-08, 6.372871e-08, 6.364956e-08, 
    6.383784e-08, 6.395748e-08, 6.389831e-08, 6.42635e-08, 6.412152e-08, 
    6.486947e-08, 6.454731e-08, 6.53872e-08, 6.518622e-08, 6.543538e-08, 
    6.530824e-08, 6.552609e-08, 6.533003e-08, 6.566965e-08, 6.57436e-08, 
    6.569307e-08, 6.588719e-08, 6.531916e-08, 6.553731e-08, 6.389665e-08, 
    6.39063e-08, 6.395126e-08, 6.375364e-08, 6.374155e-08, 6.356043e-08, 
    6.372159e-08, 6.379021e-08, 6.396441e-08, 6.406746e-08, 6.416541e-08, 
    6.438078e-08, 6.462131e-08, 6.495763e-08, 6.519925e-08, 6.536121e-08, 
    6.52619e-08, 6.534958e-08, 6.525156e-08, 6.520562e-08, 6.571589e-08, 
    6.542937e-08, 6.585927e-08, 6.583548e-08, 6.564093e-08, 6.583816e-08, 
    6.391308e-08, 6.385754e-08, 6.366474e-08, 6.381563e-08, 6.35407e-08, 
    6.369459e-08, 6.378308e-08, 6.412449e-08, 6.41995e-08, 6.426905e-08, 
    6.440642e-08, 6.458272e-08, 6.489199e-08, 6.516106e-08, 6.540669e-08, 
    6.538869e-08, 6.539503e-08, 6.54499e-08, 6.531398e-08, 6.547221e-08, 
    6.549877e-08, 6.542933e-08, 6.58323e-08, 6.571717e-08, 6.583497e-08, 
    6.576001e-08, 6.38756e-08, 6.396904e-08, 6.391854e-08, 6.40135e-08, 
    6.394661e-08, 6.424406e-08, 6.433323e-08, 6.475051e-08, 6.457925e-08, 
    6.48518e-08, 6.460694e-08, 6.465033e-08, 6.486071e-08, 6.462017e-08, 
    6.514622e-08, 6.478959e-08, 6.545203e-08, 6.50959e-08, 6.547435e-08, 
    6.540562e-08, 6.551941e-08, 6.562132e-08, 6.574952e-08, 6.598609e-08, 
    6.59313e-08, 6.612913e-08, 6.410834e-08, 6.422955e-08, 6.421887e-08, 
    6.434571e-08, 6.443951e-08, 6.464282e-08, 6.496889e-08, 6.484628e-08, 
    6.507138e-08, 6.511657e-08, 6.477458e-08, 6.498456e-08, 6.431066e-08, 
    6.441955e-08, 6.435471e-08, 6.411791e-08, 6.487454e-08, 6.448624e-08, 
    6.520325e-08, 6.49929e-08, 6.560679e-08, 6.53015e-08, 6.590115e-08, 
    6.615751e-08, 6.639875e-08, 6.668071e-08, 6.429569e-08, 6.421333e-08, 
    6.436079e-08, 6.456481e-08, 6.475408e-08, 6.500573e-08, 6.503147e-08, 
    6.507862e-08, 6.520072e-08, 6.53034e-08, 6.509353e-08, 6.532913e-08, 
    6.444481e-08, 6.490824e-08, 6.41822e-08, 6.440084e-08, 6.455278e-08, 
    6.448612e-08, 6.483226e-08, 6.491384e-08, 6.524535e-08, 6.507398e-08, 
    6.609424e-08, 6.564286e-08, 6.689538e-08, 6.654536e-08, 6.418456e-08, 
    6.429541e-08, 6.468117e-08, 6.449763e-08, 6.502253e-08, 6.515172e-08, 
    6.525676e-08, 6.539102e-08, 6.540552e-08, 6.548507e-08, 6.53547e-08, 
    6.547992e-08, 6.500627e-08, 6.521793e-08, 6.463707e-08, 6.477845e-08, 
    6.471341e-08, 6.464207e-08, 6.486225e-08, 6.509683e-08, 6.510184e-08, 
    6.517705e-08, 6.538904e-08, 6.502465e-08, 6.615252e-08, 6.545599e-08, 
    6.441627e-08, 6.462978e-08, 6.466026e-08, 6.457756e-08, 6.513877e-08, 
    6.493543e-08, 6.548313e-08, 6.53351e-08, 6.557763e-08, 6.545712e-08, 
    6.543939e-08, 6.52846e-08, 6.518822e-08, 6.494476e-08, 6.474665e-08, 
    6.458955e-08, 6.462608e-08, 6.479865e-08, 6.511118e-08, 6.540683e-08, 
    6.534207e-08, 6.55592e-08, 6.498447e-08, 6.522547e-08, 6.513232e-08, 
    6.537519e-08, 6.484301e-08, 6.529623e-08, 6.472717e-08, 6.477707e-08, 
    6.493139e-08, 6.524182e-08, 6.531049e-08, 6.538382e-08, 6.533857e-08, 
    6.511911e-08, 6.508316e-08, 6.492764e-08, 6.488471e-08, 6.47662e-08, 
    6.46681e-08, 6.475774e-08, 6.485187e-08, 6.51192e-08, 6.536012e-08, 
    6.562277e-08, 6.568705e-08, 6.599396e-08, 6.574413e-08, 6.61564e-08, 
    6.580591e-08, 6.641262e-08, 6.532247e-08, 6.579559e-08, 6.493841e-08, 
    6.503075e-08, 6.519779e-08, 6.558088e-08, 6.537405e-08, 6.561592e-08, 
    6.508175e-08, 6.480461e-08, 6.473289e-08, 6.459911e-08, 6.473595e-08, 
    6.472482e-08, 6.485576e-08, 6.481368e-08, 6.512808e-08, 6.49592e-08, 
    6.543894e-08, 6.561401e-08, 6.610841e-08, 6.641149e-08, 6.671998e-08, 
    6.685619e-08, 6.689764e-08, 6.691497e-08 ;

 SOILICE =
  57.77513, 57.96864, 57.931, 58.08735, 58.0006, 58.10302, 57.81435, 57.9763, 
    57.87289, 57.79257, 58.39167, 58.09434, 58.70219, 58.51152, 58.99155, 
    58.67244, 59.05608, 58.9824, 59.20456, 59.14085, 59.42558, 59.23398, 
    59.57373, 59.37982, 59.41009, 59.22766, 58.15414, 58.35456, 58.14227, 
    58.17081, 58.15802, 58.00236, 57.924, 57.76041, 57.7901, 57.91029, 
    58.18365, 58.09079, 58.32522, 58.31992, 58.58176, 58.46358, 58.90518, 
    58.77941, 59.14351, 59.05176, 59.13918, 59.11267, 59.13953, 59.00502, 
    59.06261, 58.94439, 58.48568, 58.62017, 58.21979, 57.98003, 57.82143, 
    57.70905, 57.72492, 57.75518, 57.91099, 58.05787, 58.16999, 58.24508, 
    58.31916, 58.54366, 58.66293, 58.9306, 58.88229, 58.96421, 59.04264, 
    59.17443, 59.15273, 59.21084, 58.96209, 59.12729, 58.85477, 58.9292, 
    58.33905, 58.11584, 58.02097, 57.93822, 57.73713, 57.87592, 57.82117, 
    57.95155, 58.03449, 57.99347, 58.24714, 58.1484, 58.67001, 58.44486, 
    59.03349, 58.89221, 59.0674, 58.97797, 59.13126, 58.99328, 59.2325, 
    59.28466, 59.249, 59.38615, 58.98563, 59.13916, 57.99231, 57.999, 
    58.03019, 57.89317, 57.88482, 57.75958, 57.87103, 57.91852, 58.03933, 
    58.11083, 58.1789, 58.32878, 58.49651, 58.7318, 58.90136, 59.01522, 
    58.9454, 59.00703, 58.93812, 58.90586, 59.26509, 59.06314, 59.36641, 
    59.34961, 59.21221, 59.3515, 58.0037, 57.96521, 57.83168, 57.93616, 
    57.74596, 57.85233, 57.91354, 58.1504, 58.20261, 58.25098, 58.34666, 
    58.46962, 58.68582, 58.8745, 59.04722, 59.03455, 59.03901, 59.07762, 
    58.98199, 59.09333, 59.11201, 59.06314, 59.34735, 59.26605, 59.34925, 
    59.29631, 57.97773, 58.04252, 58.0075, 58.07335, 58.02693, 58.23352, 
    58.29558, 58.58677, 58.46719, 58.65768, 58.48653, 58.51682, 58.66379, 
    58.49579, 58.86404, 58.61407, 59.07912, 58.82866, 59.09484, 59.04647, 
    59.12659, 59.1984, 59.28889, 59.45606, 59.41732, 59.55738, 58.13924, 
    58.22346, 58.21609, 58.30436, 58.36971, 58.5116, 58.73972, 58.65387, 
    58.81161, 58.84331, 58.60371, 58.75068, 58.27992, 58.35572, 58.31062, 
    58.14585, 58.67358, 58.40223, 58.90415, 58.75656, 59.18815, 58.97314, 
    59.396, 59.57738, 59.74871, 59.94916, 58.26952, 58.21225, 58.31488, 
    58.45705, 58.58935, 58.76554, 58.78362, 58.81667, 58.90241, 58.97456, 
    58.82708, 58.99265, 58.37321, 58.6972, 58.19056, 58.34267, 58.44868, 
    58.40221, 58.64408, 58.70118, 58.9337, 58.81344, 59.53253, 59.21351, 
    60.1023, 59.85284, 58.19223, 58.26935, 58.53835, 58.41024, 58.77735, 
    58.86798, 58.94178, 59.03615, 59.04638, 59.10237, 59.01064, 59.09876, 
    58.76592, 58.91448, 58.50761, 58.6064, 58.56095, 58.51109, 58.66507, 
    58.82938, 58.83298, 58.88574, 59.03448, 58.77884, 59.57366, 59.08165, 
    58.35354, 58.5024, 58.52378, 58.46604, 58.85888, 58.71629, 59.10102, 
    58.99685, 59.16762, 59.08271, 59.07022, 58.96134, 58.89361, 58.7228, 
    58.58414, 58.47442, 58.49993, 58.62051, 58.83947, 59.04728, 59.00169, 
    59.15463, 58.75066, 58.91974, 58.85432, 59.02504, 58.65157, 58.96925, 
    58.57057, 58.60545, 58.71346, 58.93117, 58.97954, 59.03108, 58.99929, 
    58.84505, 58.81985, 58.71085, 58.68074, 58.59786, 58.52928, 58.59192, 
    58.65775, 58.84515, 59.0144, 59.19941, 59.24479, 59.46149, 59.28493, 
    59.5764, 59.32837, 59.75832, 58.98781, 59.32124, 58.7184, 58.78313, 
    58.90026, 59.16979, 59.02424, 59.19453, 58.81886, 58.62463, 58.57456, 
    58.48108, 58.5767, 58.56892, 58.66053, 58.63108, 58.85138, 58.73296, 
    59.06988, 59.1932, 59.54267, 59.75766, 59.97726, 60.07437, 60.10395, 
    60.11632,
  78.08491, 78.38567, 78.32719, 78.56937, 78.43539, 78.59308, 78.1459, 
    78.39755, 78.23689, 78.11207, 79.02924, 78.57996, 79.49915, 79.21082, 
    79.93704, 79.45409, 80.03476, 79.92332, 80.25967, 80.16322, 80.59417, 
    80.30424, 80.81867, 80.52499, 80.57078, 80.29465, 78.67043, 78.97312, 
    78.65247, 78.69559, 78.67629, 78.4381, 78.31622, 78.0621, 78.10822, 
    78.29497, 78.71498, 78.57468, 78.92914, 78.92113, 79.31708, 79.13835, 
    79.80645, 79.61616, 80.16724, 80.02833, 80.16068, 80.12056, 80.16119, 
    79.95756, 80.04474, 79.86581, 79.17175, 79.37514, 78.76965, 78.40327, 
    78.15688, 77.98228, 78.00694, 78.05394, 78.29606, 78.52443, 78.69443, 
    78.80795, 78.91997, 79.25921, 79.43977, 79.84486, 79.77183, 79.89573, 
    80.01453, 80.21403, 80.1812, 80.26913, 79.89261, 80.14262, 79.73021, 
    79.84281, 78.94964, 78.61255, 78.46691, 78.33839, 78.02589, 78.24155, 
    78.15646, 78.35917, 78.48808, 78.42433, 78.81106, 78.66177, 79.45047, 
    79.10997, 80.00066, 79.78683, 80.05202, 79.91665, 80.14864, 79.93983, 
    80.30196, 80.38089, 80.32693, 80.53465, 79.92825, 80.1606, 78.42252, 
    78.43291, 78.48141, 78.26836, 78.25539, 78.0608, 78.23399, 78.30778, 
    78.49562, 78.60497, 78.70786, 78.93448, 79.18807, 79.54401, 79.80067, 
    79.97304, 79.86736, 79.96065, 79.85634, 79.80753, 80.35125, 80.04551, 
    80.50475, 80.47931, 80.2712, 80.48217, 78.44022, 78.38041, 78.17284, 
    78.33524, 78.03964, 78.2049, 78.30001, 78.6647, 78.74374, 78.81683, 
    78.96155, 79.14748, 79.47447, 79.75999, 80.02148, 80.00231, 80.00906, 
    80.06747, 79.92272, 80.09126, 80.1195, 80.04556, 80.47589, 80.35278, 
    80.47877, 80.39861, 78.39986, 78.50056, 78.44613, 78.54829, 78.4763, 
    78.79034, 78.88416, 79.32455, 79.14378, 79.43187, 79.17307, 79.21883, 
    79.44094, 79.18709, 79.74407, 79.36581, 80.06974, 79.69044, 80.09354, 
    80.02035, 80.14165, 80.25031, 80.38735, 80.64045, 80.58182, 80.79398, 
    78.64793, 78.77519, 78.76413, 78.89758, 78.99636, 79.211, 79.55605, 
    79.42621, 79.66489, 79.71282, 79.35035, 79.5726, 78.86057, 78.9751, 
    78.90701, 78.65788, 79.4559, 79.04545, 79.80489, 79.58155, 80.23479, 
    79.90923, 80.54952, 80.82409, 81.08388, 81.38749, 78.84488, 78.75832, 
    78.91351, 79.12836, 79.32857, 79.59513, 79.62253, 79.67252, 79.8023, 
    79.91148, 79.68819, 79.93888, 79.00138, 79.49168, 78.72546, 78.95535, 
    79.11575, 79.04551, 79.41142, 79.4978, 79.84957, 79.66766, 80.75612, 
    80.27308, 81.61976, 81.24155, 78.72805, 78.84466, 79.25137, 79.05766, 
    79.61303, 79.75015, 79.86189, 80.00466, 80.0202, 80.10492, 79.96611, 
    80.09949, 79.5957, 79.82054, 79.20497, 79.35435, 79.28566, 79.21024, 
    79.44316, 79.69165, 79.69721, 79.77699, 80.00171, 79.6153, 80.81818, 
    80.07319, 78.97195, 79.19691, 79.22939, 79.14211, 79.73639, 79.52061, 
    80.10289, 79.94524, 80.20374, 80.07518, 80.05627, 79.89148, 79.78896, 
    79.53045, 79.32068, 79.15479, 79.19336, 79.37568, 79.70693, 80.0215, 
    79.95248, 80.18407, 79.57265, 79.82845, 79.72942, 79.98788, 79.42271, 
    79.90304, 79.30022, 79.35297, 79.51633, 79.84566, 79.91903, 79.99699, 
    79.94893, 79.7154, 79.6773, 79.51242, 79.46682, 79.34151, 79.23776, 
    79.33248, 79.43201, 79.7156, 79.97173, 80.25182, 80.32059, 80.64845, 
    80.38114, 80.8223, 80.44662, 81.09808, 79.93131, 80.43607, 79.52386, 
    79.62179, 79.7989, 80.20686, 79.98666, 80.24435, 79.67583, 79.38186, 
    79.30624, 79.16483, 79.30948, 79.29771, 79.4363, 79.39176, 79.72504, 
    79.54588, 80.05573, 80.24237, 80.77164, 81.0973, 81.43025, 81.57746, 
    81.62233, 81.64108,
  118.461, 119.0176, 118.9093, 119.3593, 119.1095, 119.4044, 118.5737, 
    119.0397, 118.7421, 118.5111, 120.236, 119.3794, 121.1308, 120.5809, 
    121.9608, 121.0451, 122.141, 121.9351, 122.5557, 122.3777, 123.174, 
    122.638, 123.5883, 123.0458, 123.1305, 122.6203, 119.5515, 120.1291, 
    119.5173, 119.5995, 119.5626, 119.1147, 118.8894, 118.4186, 118.504, 
    118.8498, 119.6365, 119.369, 120.044, 120.0287, 120.7834, 120.4427, 
    121.7162, 121.3533, 122.3851, 122.1288, 122.3731, 122.299, 122.374, 
    121.9983, 122.1592, 121.829, 120.5064, 120.8941, 119.7405, 119.0507, 
    118.5941, 118.271, 118.3166, 118.4037, 118.8518, 119.2743, 119.597, 
    119.8132, 120.0266, 120.6739, 121.0176, 121.7897, 121.6501, 121.8844, 
    122.1034, 122.4716, 122.4109, 122.5733, 121.8784, 122.3399, 121.5707, 
    121.7855, 120.0845, 119.4412, 119.1684, 118.9301, 118.3517, 118.7509, 
    118.5934, 118.9684, 119.207, 119.089, 119.8191, 119.5349, 121.038, 
    120.3889, 122.0778, 121.6787, 122.1725, 121.9227, 122.351, 121.9655, 
    122.6339, 122.7797, 122.68, 123.0634, 121.9441, 122.3731, 119.0856, 
    119.1049, 119.1946, 118.8005, 118.7765, 118.4163, 118.7367, 118.8734, 
    119.2209, 119.4268, 119.6227, 120.0543, 120.5377, 121.2161, 121.7052, 
    122.0267, 121.8317, 122.0039, 121.8112, 121.7181, 122.7251, 122.1607, 
    123.0082, 122.9612, 122.5772, 122.9665, 119.1184, 119.0076, 118.6236, 
    118.9241, 118.3771, 118.683, 118.8592, 119.5408, 119.6909, 119.8303, 
    120.1058, 120.4601, 121.0835, 121.6277, 122.1161, 122.0807, 122.0932, 
    122.2011, 121.934, 122.245, 122.2972, 122.1606, 122.9549, 122.7276, 
    122.9602, 122.8122, 119.0436, 119.2301, 119.1293, 119.3189, 119.1853, 
    119.7801, 119.9589, 120.798, 120.4531, 121.0023, 120.5089, 120.5962, 
    121.0202, 120.5355, 121.5977, 120.8768, 122.2053, 121.4957, 122.2492, 
    122.114, 122.3379, 122.5386, 122.7915, 123.259, 123.1507, 123.5425, 
    119.5085, 119.7511, 119.7298, 119.984, 120.1722, 120.5811, 121.2389, 
    120.9912, 121.4462, 121.5377, 120.8466, 121.2705, 119.9137, 120.1321, 
    120.002, 119.5276, 121.0482, 120.2661, 121.7132, 121.2874, 122.5099, 
    121.9094, 123.091, 123.5986, 124.078, 124.6397, 119.8837, 119.7187, 
    120.0143, 120.424, 120.8052, 121.3133, 121.3654, 121.4608, 121.7082, 
    121.9132, 121.491, 121.9637, 120.1828, 121.1163, 119.6563, 120.0946, 
    120.3999, 120.2659, 120.9629, 121.1276, 121.7986, 121.4514, 123.4732, 
    122.581, 125.0687, 124.3698, 119.661, 119.8831, 120.6583, 120.289, 
    121.3473, 121.6088, 121.8216, 122.0853, 122.1138, 122.2702, 122.014, 
    122.2601, 121.3144, 121.743, 120.5695, 120.8544, 120.7233, 120.5796, 
    121.0235, 121.4976, 121.5078, 121.6602, 122.0812, 121.3516, 123.5886, 
    122.2129, 120.1256, 120.5548, 120.6162, 120.4498, 121.5826, 121.1712, 
    122.2664, 121.9754, 122.4525, 122.2153, 122.1804, 121.8763, 121.6828, 
    121.1901, 120.7902, 120.4739, 120.5474, 120.8951, 121.5267, 122.1164, 
    121.9891, 122.4162, 121.2704, 121.7583, 121.5695, 122.0542, 120.9846, 
    121.8989, 120.751, 120.8516, 121.1631, 121.7914, 121.9271, 122.0711, 
    121.9823, 121.5428, 121.47, 121.1555, 121.0688, 120.8297, 120.632, 
    120.8126, 121.0025, 121.543, 122.0246, 122.5414, 122.6682, 123.2745, 
    122.7807, 123.5963, 122.9025, 124.1053, 121.9505, 122.8823, 121.1773, 
    121.364, 121.7022, 122.4588, 122.052, 122.5279, 121.4671, 120.9071, 
    120.7625, 120.4931, 120.7687, 120.7463, 121.0104, 120.9255, 121.5609, 
    121.2193, 122.1795, 122.5241, 123.5013, 124.1032, 124.7182, 124.9903, 
    125.0733, 125.1079,
  187.2937, 188.2959, 188.1007, 188.9114, 188.4613, 188.9927, 187.4965, 
    188.3358, 187.7997, 187.3837, 190.4924, 188.9476, 192.1069, 191.1142, 
    193.6134, 191.9522, 193.9387, 193.5668, 194.6876, 194.366, 195.8053, 
    194.8362, 196.5545, 195.5734, 195.7267, 194.8043, 189.2576, 190.2996, 
    189.1961, 189.3443, 189.2778, 188.4707, 188.065, 187.2172, 187.3709, 
    187.9936, 189.411, 188.9289, 190.1456, 190.1181, 191.4796, 190.8648, 
    193.1642, 192.5085, 194.3794, 193.9165, 194.3577, 194.2238, 194.3594, 
    193.6809, 193.9714, 193.3686, 190.9798, 191.6796, 189.5984, 188.3556, 
    187.5333, 186.9515, 187.0337, 187.1904, 187.9973, 188.7582, 189.3397, 
    189.7295, 190.1141, 191.2822, 191.9025, 193.2971, 193.0447, 193.4723, 
    193.8705, 194.5356, 194.426, 194.7195, 193.4609, 194.2978, 192.9011, 
    193.2894, 190.2191, 189.0589, 188.5676, 188.1382, 187.0969, 187.8156, 
    187.532, 188.2071, 188.637, 188.4243, 189.7402, 189.2278, 191.9393, 
    190.7677, 193.8244, 193.0965, 193.9954, 193.5437, 194.3178, 193.6216, 
    194.8288, 195.0925, 194.9122, 195.6052, 193.583, 194.3577, 188.4183, 
    188.453, 188.6147, 187.905, 187.8616, 187.213, 187.79, 188.0361, 188.662, 
    189.0329, 189.3861, 190.1643, 191.0364, 192.2608, 193.1442, 193.7322, 
    193.3737, 193.6909, 193.3359, 193.1675, 194.9937, 193.9741, 195.5054, 
    195.4204, 194.7265, 195.43, 188.4774, 188.2778, 187.5863, 188.1273, 
    187.1425, 187.6933, 188.0106, 189.2385, 189.5091, 189.7603, 190.2571, 
    190.8962, 192.0213, 193.0044, 193.8935, 193.8297, 193.8521, 194.047, 
    193.5647, 194.1263, 194.2207, 193.974, 195.409, 194.9982, 195.4186, 
    195.151, 188.3427, 188.6786, 188.497, 188.8386, 188.5979, 189.67, 
    189.9923, 191.5061, 190.8836, 191.8749, 190.9841, 191.1418, 191.9074, 
    191.0322, 192.9501, 191.6483, 194.0546, 192.7661, 194.1339, 193.8898, 
    194.294, 194.6566, 195.1136, 195.959, 195.7629, 196.4716, 189.1803, 
    189.6176, 189.579, 190.0374, 190.3769, 191.1144, 192.3019, 191.8547, 
    192.6763, 192.8416, 191.5936, 192.3591, 189.9107, 190.3047, 190.07, 
    189.2148, 191.9578, 190.5463, 193.1588, 192.3896, 194.6049, 193.519, 
    195.6551, 196.5734, 197.4406, 198.4581, 189.8565, 189.559, 190.0919, 
    190.8312, 191.519, 192.4364, 192.5304, 192.7028, 193.1496, 193.5259, 
    192.7573, 193.6184, 190.3962, 192.0806, 189.4467, 190.237, 190.7876, 
    190.5458, 191.8036, 192.101, 193.3131, 192.6858, 196.3465, 194.7334, 
    199.2354, 197.9691, 189.4552, 189.8555, 191.2539, 190.5875, 192.4978, 
    192.9702, 193.3549, 193.838, 193.8894, 194.1719, 193.7091, 194.1536, 
    192.4384, 193.2126, 191.0936, 191.6077, 191.371, 191.1117, 191.9129, 
    192.7694, 192.7877, 193.063, 193.831, 192.5055, 196.5556, 194.0688, 
    190.2928, 191.0671, 191.1778, 190.8775, 192.9228, 192.1798, 194.165, 
    193.6395, 194.5011, 194.0726, 194.0096, 193.457, 193.1038, 192.2138, 
    191.492, 190.921, 191.0536, 191.6813, 192.8219, 193.8941, 193.6643, 
    194.4355, 192.3588, 193.2403, 192.8992, 193.7818, 191.8428, 193.4998, 
    191.4211, 191.6027, 192.1651, 193.3002, 193.5519, 193.8124, 193.6518, 
    192.8509, 192.7194, 192.1514, 191.9948, 191.5631, 191.2063, 191.5323, 
    191.8751, 192.8512, 193.7283, 194.6618, 194.8908, 195.9872, 195.0944, 
    196.5695, 195.315, 197.4906, 193.5948, 195.278, 192.1907, 192.5278, 
    193.1389, 194.5127, 193.7777, 194.6375, 192.7142, 191.703, 191.4419, 
    190.9557, 191.453, 191.4125, 191.8893, 191.736, 192.8837, 192.2665, 
    194.0081, 194.6306, 196.3972, 197.4865, 198.6, 199.0932, 199.2435, 
    199.3064,
  314.8134, 316.5515, 316.2129, 317.6201, 316.8387, 317.7612, 315.165, 
    316.6208, 315.6906, 314.9694, 320.3683, 317.683, 323.18, 321.4505, 
    325.8118, 322.9104, 326.3999, 325.7276, 327.7546, 327.1727, 329.768, 
    328.0236, 331.0811, 329.3589, 329.6303, 327.9658, 318.2215, 320.0328, 
    318.1145, 318.3721, 318.2564, 316.8548, 316.1508, 314.6808, 314.9472, 
    316.0271, 318.488, 317.6505, 319.765, 319.717, 322.0868, 321.0162, 
    325.0244, 323.8803, 327.1969, 326.3598, 327.1576, 326.9155, 327.1607, 
    325.9338, 326.459, 325.3813, 321.2165, 322.4352, 318.8137, 316.6551, 
    315.2287, 314.2204, 314.3628, 314.6343, 316.0334, 317.354, 318.364, 
    319.0414, 319.7102, 321.7431, 322.8237, 325.2563, 324.8158, 325.5622, 
    326.2766, 327.4796, 327.2813, 327.8124, 325.5424, 327.0494, 324.5652, 
    325.2429, 319.8928, 317.8762, 317.0232, 316.278, 314.4723, 315.7182, 
    315.2265, 316.3974, 317.1436, 316.7743, 319.06, 318.1695, 322.8878, 
    320.8473, 326.1932, 324.9062, 326.5024, 325.6869, 327.0854, 325.8265, 
    328.0102, 328.4876, 328.1613, 329.4164, 325.7569, 327.1577, 316.764, 
    316.8242, 317.1048, 315.8733, 315.798, 314.6736, 315.6739, 316.1008, 
    317.1869, 317.8311, 318.4445, 319.7974, 321.3149, 323.4484, 324.9895, 
    326.0265, 325.3902, 325.9519, 325.324, 325.0302, 328.3087, 326.4639, 
    329.2356, 329.0816, 327.825, 329.0989, 316.8665, 316.5201, 315.3207, 
    316.259, 314.5513, 315.5062, 316.0565, 318.1882, 318.6583, 319.0949, 
    319.9589, 321.071, 323.0309, 324.7454, 326.3182, 326.2027, 326.2433, 
    326.5957, 325.7237, 326.739, 326.9098, 326.4636, 329.0609, 328.3169, 
    329.0783, 328.5936, 316.6327, 317.2158, 316.9006, 317.4936, 317.0757, 
    318.938, 319.4984, 322.133, 321.0491, 322.7756, 321.224, 321.4984, 
    322.8323, 321.3076, 324.6508, 322.3808, 326.6094, 324.3297, 326.7528, 
    326.3114, 327.0424, 327.6986, 328.5258, 330.0372, 329.6938, 330.9356, 
    318.087, 318.8469, 318.7798, 319.5767, 320.1673, 321.4509, 323.52, 
    322.7404, 324.1729, 324.4613, 322.2854, 323.6198, 319.3564, 320.0416, 
    319.6334, 318.1469, 322.92, 320.462, 325.015, 323.6728, 327.605, 
    325.6439, 329.5049, 331.1143, 332.6356, 334.423, 319.2623, 318.7451, 
    319.6716, 320.9579, 322.1555, 323.7545, 323.9185, 324.2191, 324.9988, 
    325.6559, 324.3143, 325.8208, 320.201, 323.1342, 318.5499, 319.9239, 
    320.8819, 320.4612, 322.6514, 323.1697, 325.2844, 324.1895, 330.7164, 
    327.8376, 335.7901, 333.5638, 318.5646, 319.2604, 321.6937, 320.5337, 
    323.8615, 324.6858, 325.3572, 326.2177, 326.3107, 326.8217, 325.9847, 
    326.7885, 323.758, 325.1089, 321.4145, 322.31, 321.8977, 321.4461, 
    322.8419, 324.3354, 324.3672, 324.8477, 326.2054, 323.8751, 331.0831, 
    326.6353, 320.0208, 321.3686, 321.5613, 321.0383, 324.6031, 323.3071, 
    326.8092, 325.859, 327.4171, 326.642, 326.5281, 325.5355, 324.919, 
    323.3664, 322.1084, 321.1141, 321.345, 322.4382, 324.427, 326.3192, 
    325.9038, 327.2985, 323.6191, 325.1572, 324.5619, 326.1161, 322.7198, 
    325.6104, 321.9849, 322.3012, 323.2814, 325.2619, 325.7013, 326.1715, 
    325.8813, 324.4776, 324.2481, 323.2575, 322.9846, 322.2323, 321.6108, 
    322.1786, 322.776, 324.4781, 326.0195, 327.708, 328.1224, 330.0868, 
    328.4912, 331.1076, 328.8909, 332.7236, 325.7784, 328.8238, 323.326, 
    323.914, 324.9802, 327.4382, 326.1088, 327.664, 324.2391, 322.476, 
    322.0211, 321.1745, 322.0405, 321.97, 322.8007, 322.5335, 324.5348, 
    323.4583, 326.5253, 327.6516, 330.8053, 332.7162, 334.6725, 335.54, 
    335.8044, 335.9151,
  523.2206, 526.4933, 525.8551, 528.5091, 527.0347, 528.7756, 523.882, 
    526.6239, 524.8715, 523.514, 533.7067, 528.6278, 539.0443, 535.7587, 
    544.0591, 538.5316, 545.1821, 543.8983, 547.7728, 546.6593, 551.6535, 
    548.2877, 554.2643, 550.8471, 551.3801, 548.1771, 529.6448, 533.0712, 
    529.4427, 529.9294, 529.7109, 527.0652, 525.7383, 522.9713, 523.4722, 
    525.5051, 530.1485, 528.5665, 532.564, 532.4733, 536.9666, 534.9349, 
    542.5568, 540.3768, 546.7057, 545.1055, 546.6305, 546.1675, 546.6365, 
    544.2919, 545.295, 543.2374, 535.3147, 537.6284, 530.7641, 526.6887, 
    524.002, 522.1057, 522.3732, 522.8839, 525.517, 528.007, 529.9142, 
    531.1948, 532.4602, 536.314, 538.3668, 542.999, 542.1591, 543.5827, 
    544.9466, 547.2465, 546.8671, 547.8834, 543.5449, 546.4236, 541.6815, 
    542.9734, 532.806, 528.9926, 527.3828, 525.9777, 522.5791, 524.9233, 
    523.9977, 526.2028, 527.6099, 526.9134, 531.2299, 529.5467, 538.4887, 
    534.6146, 544.7873, 542.3314, 545.378, 543.8206, 546.4926, 544.0871, 
    548.2621, 549.1766, 548.5515, 550.9573, 543.9542, 546.6306, 526.8939, 
    527.0074, 527.5366, 525.2153, 525.0737, 522.9576, 524.8398, 525.644, 
    527.6916, 528.9075, 530.0664, 532.6254, 535.5015, 539.5549, 542.4902, 
    544.4689, 543.2544, 544.3264, 543.1282, 542.5677, 548.8339, 545.3044, 
    550.6105, 550.3152, 547.9076, 550.3484, 527.0872, 526.4342, 524.175, 
    525.942, 522.7278, 524.5242, 525.5605, 529.5821, 530.4703, 531.296, 
    532.9311, 535.0386, 538.7606, 542.0249, 545.026, 544.8054, 544.8831, 
    545.5562, 543.8909, 545.8303, 546.1567, 545.3038, 550.2756, 548.8495, 
    550.3089, 549.3797, 526.6463, 527.7462, 527.1515, 528.2704, 527.4819, 
    530.9993, 532.0594, 537.0543, 534.9971, 538.2753, 535.3289, 535.8496, 
    538.3832, 535.4875, 541.8445, 537.525, 545.5824, 541.2326, 545.8564, 
    545.013, 546.4103, 547.6656, 549.2498, 552.1884, 551.5061, 553.9747, 
    529.3908, 530.827, 530.7001, 532.2076, 533.3259, 535.7593, 539.6911, 
    538.2084, 540.9341, 541.4834, 537.3438, 539.881, 531.7906, 533.0879, 
    532.3149, 529.504, 538.5499, 533.8842, 542.5389, 539.9819, 547.4865, 
    543.7385, 551.131, 554.3303, 557.2731, 560.7239, 531.6125, 530.6345, 
    532.3871, 534.8242, 537.097, 540.1375, 540.4496, 541.0221, 542.508, 
    543.7614, 541.2034, 544.0762, 533.3897, 538.9572, 530.2654, 532.8648, 
    534.6801, 533.8826, 538.0392, 539.0247, 543.0526, 540.9656, 553.5388, 
    547.9316, 563.3696, 559.064, 530.2933, 531.6091, 536.2202, 534.0201, 
    540.3411, 541.9112, 543.1916, 544.8341, 545.0117, 545.9882, 544.3892, 
    545.9248, 540.144, 542.7178, 535.6904, 537.3906, 536.6075, 535.7504, 
    538.4012, 541.2437, 541.3042, 542.2197, 544.8107, 540.3669, 554.2684, 
    545.6319, 533.0485, 535.6032, 535.9689, 534.9767, 541.7535, 539.2859, 
    545.9643, 544.1492, 547.127, 545.6448, 545.4272, 543.5316, 542.3558, 
    539.3989, 537.0076, 535.1204, 535.5585, 537.634, 541.418, 545.0279, 
    544.2347, 546.9, 539.8797, 542.8099, 541.6752, 544.6401, 538.1691, 
    543.6746, 536.7731, 537.3738, 539.2371, 543.0096, 543.8481, 544.7458, 
    544.1917, 541.5145, 541.0773, 539.1917, 538.6726, 537.2429, 536.0629, 
    537.141, 538.2761, 541.5154, 544.4556, 547.6836, 548.4771, 552.2869, 
    549.1835, 554.3171, 549.9496, 557.4429, 543.9952, 549.821, 539.322, 
    540.4409, 542.4725, 547.1673, 544.6261, 547.5993, 541.0601, 537.7059, 
    536.8419, 535.235, 536.8787, 536.7448, 538.3229, 537.8151, 541.6234, 
    539.5736, 545.4218, 547.5756, 553.7155, 557.4286, 561.2064, 562.8851, 
    563.3974, 563.6117,
  947.1248, 953.9976, 952.6545, 958.2484, 955.1379, 958.8113, 948.5109, 
    954.2725, 950.5872, 947.7395, 969.1224, 958.4991, 980.1622, 973.3553, 
    990.6236, 979.0976, 992.9783, 990.2868, 998.4278, 996.0826, 1006.636, 
    999.5137, 1012.19, 1004.926, 1006.056, 999.2805, 960.6494, 967.8145, 
    960.2218, 961.2517, 960.7892, 955.2023, 952.4089, 946.6025, 947.6519, 
    951.9185, 961.7155, 958.3695, 966.7713, 966.5849, 975.8534, 971.6542, 
    987.4803, 982.9335, 996.1803, 992.8176, 996.022, 995.0482, 996.0347, 
    991.1115, 993.2153, 988.9034, 972.4383, 977.2244, 963.0198, 954.4091, 
    948.7624, 944.7913, 945.3509, 946.4196, 951.9435, 957.1882, 961.2195, 
    963.933, 966.5581, 974.5031, 978.7556, 988.4049, 986.6498, 989.626, 
    992.4842, 997.3187, 996.5198, 998.6609, 989.5468, 995.5867, 985.6528, 
    988.3514, 967.2691, 959.27, 955.8716, 952.9125, 945.7816, 950.6962, 
    948.7536, 953.3861, 956.3506, 954.8823, 964.0074, 960.4417, 979.0087, 
    970.9935, 992.15, 987.0095, 993.3895, 990.1241, 995.7318, 990.6823, 
    999.4597, 1001.391, 1000.07, 1005.16, 990.4038, 996.0222, 954.8413, 
    955.0805, 956.196, 951.3096, 951.012, 946.5739, 950.5209, 952.2106, 
    956.5228, 959.0901, 961.5416, 966.8977, 972.8239, 981.2234, 987.3412, 
    991.4822, 988.939, 991.1837, 988.6751, 987.5033, 1000.667, 993.235, 
    1004.425, 1003.799, 998.712, 1003.87, 955.2485, 953.8731, 949.1253, 
    952.8373, 946.0928, 949.858, 952.0351, 960.5165, 962.3972, 964.1478, 
    967.5262, 971.8683, 979.5732, 986.3696, 992.6508, 992.188, 992.3509, 
    993.7639, 990.2712, 994.3394, 995.0255, 993.2339, 1003.715, 1000.7, 
    1003.786, 1001.82, 954.3198, 956.6379, 955.384, 957.7443, 956.0806, 
    963.5183, 965.7346, 976.035, 971.7827, 978.5659, 972.4675, 973.5432, 
    978.7897, 972.7952, 985.993, 977.0103, 993.8188, 984.7166, 994.3945, 
    992.6235, 995.5588, 998.2018, 1001.545, 1007.772, 1006.323, 1011.572, 
    960.1119, 963.153, 962.8842, 966.0391, 968.3386, 973.3566, 981.5068, 
    978.427, 984.0943, 985.2396, 976.6346, 981.9017, 965.1827, 967.8488, 
    966.2595, 960.3514, 979.1357, 969.4882, 987.443, 982.1116, 997.8243, 
    989.9521, 1005.528, 1012.33, 1018.811, 1026.49, 964.8172, 962.7449, 
    966.408, 971.426, 976.1237, 982.4354, 983.0851, 984.2776, 987.3785, 
    990.0002, 984.6558, 990.6594, 968.4699, 979.9814, 961.9631, 967.3899, 
    971.1287, 969.4849, 978.076, 980.1216, 988.5169, 984.1601, 1010.644, 
    998.7625, 1032.29, 1022.79, 962.0221, 964.8101, 974.3091, 969.7681, 
    982.8591, 986.1322, 988.8076, 992.2482, 992.6207, 994.6713, 991.3152, 
    994.5381, 982.4489, 987.817, 973.2141, 976.7316, 975.1104, 973.3381, 
    978.8272, 984.7396, 984.8658, 986.7764, 992.1991, 982.9128, 1012.198, 
    993.9227, 967.7677, 973.034, 973.7896, 971.7406, 985.8032, 980.6644, 
    994.6211, 990.8124, 997.0671, 993.9498, 993.4928, 989.5191, 987.0604, 
    980.8991, 975.9384, 972.0372, 972.9417, 977.236, 985.1032, 992.6548, 
    990.9914, 996.5891, 981.899, 988.0095, 985.6396, 991.8413, 978.3456, 
    989.8184, 975.4529, 976.6968, 980.5629, 988.4271, 990.1817, 992.0631, 
    990.9012, 985.3043, 984.3926, 980.4684, 979.3905, 976.4257, 973.984, 
    976.2146, 978.5675, 985.3063, 991.4543, 998.2397, 999.9133, 1007.981, 
    1001.405, 1012.302, 1003.025, 1019.188, 990.4897, 1002.753, 980.7393, 
    983.067, 987.3044, 997.152, 991.812, 998.0621, 984.3569, 977.3852, 
    975.5953, 972.2737, 975.6715, 975.3943, 978.6646, 977.6115, 985.5316, 
    981.2624, 993.4815, 998.0122, 1011.02, 1019.156, 1027.567, 1031.239, 
    1032.35, 1032.816,
  1829.886, 1849.348, 1845.52, 1861.544, 1852.608, 1863.169, 1833.786, 
    1850.133, 1839.651, 1831.614, 1893.766, 1862.268, 1928.089, 1906.809, 
    1960.685, 1924.735, 1968.115, 1959.626, 1985.501, 1977.986, 2012.206, 
    1988.998, 2030.642, 2006.59, 2010.298, 1988.246, 1868.489, 1889.765, 
    1867.249, 1870.237, 1868.894, 1852.792, 1844.821, 1828.42, 1831.368, 
    1843.427, 1871.585, 1861.894, 1886.584, 1886.016, 1914.574, 1901.55, 
    1950.842, 1936.753, 1978.298, 1967.606, 1977.792, 1974.687, 1977.833, 
    1962.22, 1968.865, 1955.288, 1903.971, 1918.857, 1875.385, 1850.523, 
    1834.495, 1823.349, 1824.913, 1827.906, 1843.498, 1858.491, 1870.144, 
    1878.052, 1885.935, 1910.37, 1923.66, 1953.728, 1948.255, 1957.552, 
    1966.552, 1981.941, 1979.383, 1986.251, 1957.303, 1976.403, 1945.158, 
    1953.561, 1888.101, 1864.494, 1854.71, 1846.254, 1826.119, 1839.96, 
    1834.47, 1847.603, 1856.084, 1851.876, 1878.27, 1867.887, 1924.456, 
    1899.514, 1965.496, 1949.375, 1969.418, 1959.115, 1976.866, 1960.869, 
    1988.824, 1995.068, 1990.795, 2007.356, 1959.994, 1977.793, 1851.759, 
    1852.443, 1855.64, 1841.699, 1840.855, 1828.339, 1839.463, 1844.257, 
    1856.578, 1863.974, 1871.08, 1886.969, 1905.163, 1931.442, 1950.408, 
    1963.389, 1955.399, 1962.448, 1954.573, 1950.913, 1992.722, 1968.928, 
    2004.949, 2002.904, 1986.415, 2003.134, 1852.924, 1848.992, 1835.518, 
    1846.04, 1826.99, 1837.588, 1843.758, 1868.104, 1873.57, 1878.68, 
    1888.885, 1902.211, 1926.232, 1947.384, 1967.079, 1965.616, 1966.13, 
    1970.605, 1959.577, 1972.432, 1974.615, 1968.924, 2002.631, 1992.829, 
    2002.861, 1996.46, 1850.268, 1856.909, 1853.312, 1860.092, 1855.309, 
    1876.84, 1883.43, 1915.141, 1901.946, 1923.064, 1904.062, 1907.391, 
    1923.767, 1905.075, 1946.214, 1918.187, 1970.779, 1942.257, 1972.608, 
    1966.992, 1976.314, 1984.775, 1995.569, 2015.952, 2011.177, 2028.578, 
    1866.931, 1875.773, 1874.989, 1884.356, 1891.367, 1906.813, 1932.338, 
    1922.628, 1940.333, 1943.877, 1917.013, 1933.58, 1881.755, 1889.87, 
    1885.026, 1867.625, 1924.855, 1894.888, 1950.725, 1934.225, 1983.562, 
    1958.575, 2008.563, 2031.113, 2053.029, 2079.234, 1880.647, 1874.583, 
    1885.478, 1900.846, 1915.417, 1935.22, 1937.22, 1940.9, 1950.524, 
    1958.726, 1942.069, 1960.797, 1891.769, 1927.519, 1872.306, 1888.469, 
    1899.93, 1894.878, 1921.526, 1927.961, 1954.078, 1940.536, 2025.48, 
    1986.578, 2099.502, 2066.699, 1872.477, 1880.625, 1909.768, 1895.747, 
    1936.524, 1946.646, 1954.988, 1965.806, 1966.983, 1973.488, 1962.862, 
    1973.064, 1935.261, 1951.892, 1906.371, 1917.316, 1912.259, 1906.755, 
    1923.885, 1942.328, 1942.719, 1948.649, 1965.651, 1936.689, 2030.672, 
    1971.109, 1889.623, 1905.814, 1908.155, 1901.817, 1945.625, 1929.674, 
    1973.328, 1961.279, 1981.135, 1971.195, 1969.745, 1957.216, 1949.533, 
    1930.416, 1914.839, 1902.732, 1905.528, 1918.894, 1943.454, 1967.091, 
    1961.842, 1979.605, 1933.571, 1952.493, 1945.117, 1964.521, 1922.372, 
    1958.155, 1913.326, 1917.207, 1929.354, 1953.797, 1959.296, 1965.221, 
    1961.558, 1944.077, 1941.255, 1929.055, 1925.657, 1916.36, 1908.758, 
    1915.701, 1923.069, 1944.083, 1963.301, 1984.896, 1990.287, 2016.644, 
    1995.115, 2031.019, 2000.38, 2054.315, 1960.264, 1999.495, 1929.911, 
    1937.164, 1950.293, 1981.406, 1964.429, 1984.326, 1941.145, 1919.361, 
    1913.769, 1903.462, 1914.007, 1913.143, 1923.374, 1920.069, 1944.782, 
    1931.565, 1969.709, 1984.166, 2026.734, 2054.207, 2082.894, 2095.755, 
    2099.718, 2101.382,
  5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597,
  8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILLIQ =
  4.537545, 4.556073, 4.552467, 4.567442, 4.55913, 4.568943, 4.541296, 
    4.556811, 4.546902, 4.53921, 4.596604, 4.568111, 4.626322, 4.608057, 
    4.654032, 4.623478, 4.660209, 4.653146, 4.674419, 4.668318, 4.695602, 
    4.677237, 4.709784, 4.69121, 4.694114, 4.676632, 4.573833, 4.59305, 
    4.572697, 4.575433, 4.574205, 4.559302, 4.551806, 4.53613, 4.538973, 
    4.550488, 4.576664, 4.567765, 4.590211, 4.589704, 4.614782, 4.603463, 
    4.645752, 4.633706, 4.668572, 4.659788, 4.66816, 4.66562, 4.668193, 
    4.655313, 4.660829, 4.649506, 4.605582, 4.618462, 4.580122, 4.557177, 
    4.541976, 4.531213, 4.532734, 4.535634, 4.550555, 4.564613, 4.575348, 
    4.582538, 4.589631, 4.61115, 4.622563, 4.648191, 4.643558, 4.651408, 
    4.658914, 4.671536, 4.669457, 4.675024, 4.6512, 4.667025, 4.64092, 
    4.64805, 4.591567, 4.570164, 4.561094, 4.55316, 4.533903, 4.547196, 
    4.541953, 4.554432, 4.562375, 4.558445, 4.582735, 4.573281, 4.62324, 
    4.601676, 4.658038, 4.644508, 4.661285, 4.652719, 4.667403, 4.654186, 
    4.677096, 4.682096, 4.678679, 4.691811, 4.653454, 4.66816, 4.558335, 
    4.558976, 4.561962, 4.548849, 4.548047, 4.536052, 4.546723, 4.551273, 
    4.562835, 4.569685, 4.576203, 4.590556, 4.606623, 4.629153, 4.645384, 
    4.656287, 4.649599, 4.655503, 4.648904, 4.645813, 4.680223, 4.660881, 
    4.689921, 4.688311, 4.675157, 4.688492, 4.559426, 4.555739, 4.542957, 
    4.552958, 4.534748, 4.544936, 4.550801, 4.57348, 4.578472, 4.583106, 
    4.592267, 4.604042, 4.624749, 4.642817, 4.659351, 4.658138, 4.658565, 
    4.662264, 4.653105, 4.663769, 4.665561, 4.660878, 4.688095, 4.680308, 
    4.688276, 4.683205, 4.556937, 4.563143, 4.559789, 4.566098, 4.561653, 
    4.581441, 4.587386, 4.61527, 4.60381, 4.622056, 4.605661, 4.608563, 
    4.622654, 4.606545, 4.64182, 4.617887, 4.662408, 4.638439, 4.663913, 
    4.659279, 4.666952, 4.673832, 4.682496, 4.698512, 4.694799, 4.708213, 
    4.572404, 4.580474, 4.579762, 4.588216, 4.594475, 4.60806, 4.629908, 
    4.621684, 4.636788, 4.639825, 4.616879, 4.63096, 4.585879, 4.593144, 
    4.588817, 4.573041, 4.62358, 4.597596, 4.645653, 4.631519, 4.672851, 
    4.652266, 4.692757, 4.710142, 4.726535, 4.745749, 4.584881, 4.579393, 
    4.589221, 4.602846, 4.615508, 4.63238, 4.634109, 4.637275, 4.645483, 
    4.652392, 4.638278, 4.654126, 4.594832, 4.625839, 4.577321, 4.591896, 
    4.602041, 4.597588, 4.620744, 4.626214, 4.648487, 4.636963, 4.705848, 
    4.675288, 4.760407, 4.736519, 4.577477, 4.584862, 4.610628, 4.598356, 
    4.633508, 4.642189, 4.649253, 4.658296, 4.659272, 4.664636, 4.655848, 
    4.664288, 4.632416, 4.646641, 4.607676, 4.61714, 4.612784, 4.60801, 
    4.622755, 4.6385, 4.638835, 4.643892, 4.658167, 4.63365, 4.709806, 
    4.66268, 4.592923, 4.60719, 4.609228, 4.603696, 4.641318, 4.627663, 
    4.664505, 4.654528, 4.670882, 4.66275, 4.661555, 4.651127, 4.644643, 
    4.628288, 4.61501, 4.604498, 4.606941, 4.618493, 4.639464, 4.659361, 
    4.654998, 4.669637, 4.630953, 4.647149, 4.640885, 4.657228, 4.621466, 
    4.651915, 4.613705, 4.617046, 4.627392, 4.64825, 4.65287, 4.65781, 
    4.654761, 4.639997, 4.63758, 4.62714, 4.624261, 4.616319, 4.609752, 
    4.615752, 4.62206, 4.640002, 4.656213, 4.67393, 4.678272, 4.699048, 
    4.682134, 4.71007, 4.686316, 4.727483, 4.65368, 4.685615, 4.627862, 
    4.63406, 4.645288, 4.671103, 4.657152, 4.673469, 4.637486, 4.618893, 
    4.614088, 4.605137, 4.614293, 4.613548, 4.62232, 4.619499, 4.640599, 
    4.629257, 4.661526, 4.673339, 4.706807, 4.727403, 4.748426, 4.757728, 
    4.760561, 4.761745,
  5.631596, 5.65485, 5.650323, 5.669121, 5.658687, 5.671004, 5.636303, 
    5.655776, 5.643338, 5.633685, 5.705736, 5.66996, 5.743062, 5.720119, 
    5.777877, 5.739489, 5.78564, 5.776764, 5.8035, 5.795831, 5.83013, 
    5.807041, 5.847961, 5.824608, 5.828258, 5.806281, 5.677144, 5.701274, 
    5.675717, 5.679153, 5.67761, 5.658903, 5.649494, 5.629819, 5.633387, 
    5.647839, 5.680698, 5.669526, 5.697708, 5.697071, 5.728565, 5.714349, 
    5.767473, 5.752337, 5.796151, 5.78511, 5.795633, 5.79244, 5.795674, 
    5.779488, 5.786419, 5.77219, 5.71701, 5.733188, 5.685039, 5.656235, 
    5.637156, 5.62365, 5.625557, 5.629197, 5.647923, 5.66557, 5.679046, 
    5.688074, 5.696979, 5.724004, 5.73834, 5.770538, 5.764716, 5.77458, 
    5.784013, 5.799877, 5.797263, 5.80426, 5.774318, 5.794206, 5.761401, 
    5.770361, 5.69941, 5.672538, 5.661152, 5.651193, 5.627025, 5.643707, 
    5.637127, 5.65279, 5.66276, 5.657827, 5.688321, 5.676451, 5.739191, 
    5.712104, 5.782912, 5.76591, 5.786992, 5.776227, 5.794682, 5.778071, 
    5.806866, 5.81315, 5.808855, 5.825363, 5.777151, 5.795633, 5.657689, 
    5.658494, 5.662241, 5.645782, 5.644775, 5.629722, 5.643114, 5.648825, 
    5.663338, 5.671937, 5.680119, 5.698141, 5.718318, 5.746618, 5.767011, 
    5.780711, 5.772307, 5.779726, 5.771433, 5.767549, 5.810795, 5.786484, 
    5.822987, 5.820962, 5.804427, 5.82119, 5.659058, 5.65443, 5.638387, 
    5.650939, 5.628085, 5.64087, 5.648232, 5.676701, 5.682968, 5.688787, 
    5.700289, 5.715076, 5.741086, 5.763785, 5.784561, 5.783037, 5.783574, 
    5.788223, 5.776713, 5.790114, 5.792366, 5.78648, 5.820691, 5.810903, 
    5.82092, 5.814544, 5.655934, 5.663724, 5.659514, 5.667433, 5.661854, 
    5.686696, 5.69416, 5.729178, 5.714786, 5.737702, 5.71711, 5.720755, 
    5.738454, 5.718221, 5.762533, 5.732467, 5.788404, 5.758285, 5.790295, 
    5.784472, 5.794115, 5.802762, 5.813653, 5.833788, 5.829121, 5.845986, 
    5.675351, 5.685482, 5.684588, 5.695202, 5.703063, 5.720123, 5.747567, 
    5.737235, 5.756211, 5.760026, 5.731201, 5.748888, 5.692269, 5.701391, 
    5.695957, 5.67615, 5.739617, 5.706982, 5.767349, 5.74959, 5.801529, 
    5.775659, 5.826553, 5.848412, 5.869029, 5.893198, 5.691015, 5.684125, 
    5.696465, 5.713574, 5.729477, 5.750673, 5.752844, 5.756822, 5.767135, 
    5.775817, 5.758082, 5.777995, 5.703511, 5.742455, 5.681523, 5.699823, 
    5.712564, 5.706971, 5.736055, 5.742926, 5.770909, 5.75643, 5.843013, 
    5.804592, 5.911641, 5.881587, 5.681719, 5.690991, 5.723348, 5.707935, 
    5.752089, 5.762996, 5.771872, 5.783236, 5.784462, 5.791203, 5.78016, 
    5.790766, 5.750718, 5.768589, 5.71964, 5.731527, 5.726056, 5.72006, 
    5.73858, 5.758362, 5.758782, 5.765136, 5.783074, 5.752268, 5.84799, 
    5.788745, 5.701114, 5.71903, 5.72159, 5.714643, 5.761902, 5.744746, 
    5.791039, 5.778501, 5.799054, 5.788834, 5.787332, 5.774227, 5.766079, 
    5.745532, 5.728852, 5.71565, 5.718717, 5.733227, 5.759573, 5.784575, 
    5.779091, 5.79749, 5.748879, 5.769228, 5.761358, 5.781895, 5.736961, 
    5.775217, 5.727213, 5.73141, 5.744405, 5.770612, 5.776417, 5.782626, 
    5.778794, 5.760242, 5.757205, 5.744089, 5.740472, 5.730496, 5.722248, 
    5.729784, 5.737708, 5.760249, 5.780619, 5.802886, 5.808343, 5.834462, 
    5.813198, 5.848321, 5.818456, 5.870221, 5.777435, 5.817574, 5.744997, 
    5.752783, 5.76689, 5.799332, 5.781798, 5.802306, 5.757086, 5.733729, 
    5.727694, 5.716452, 5.727952, 5.727015, 5.738034, 5.734491, 5.760998, 
    5.746749, 5.787295, 5.802143, 5.844218, 5.870121, 5.896566, 5.908269, 
    5.911834, 5.913325,
  8.097835, 8.132032, 8.125374, 8.153026, 8.137675, 8.155797, 8.104757, 
    8.133393, 8.115102, 8.100906, 8.20691, 8.154261, 8.261874, 8.228086, 
    8.313172, 8.256612, 8.324615, 8.311533, 8.350945, 8.339639, 8.39022, 
    8.356168, 8.41653, 8.382075, 8.38746, 8.355046, 8.16483, 8.200341, 
    8.162731, 8.167786, 8.165517, 8.137994, 8.124155, 8.095223, 8.10047, 
    8.12172, 8.170059, 8.153622, 8.195093, 8.194155, 8.240523, 8.219591, 
    8.297839, 8.275538, 8.34011, 8.323833, 8.339346, 8.33464, 8.339407, 
    8.315546, 8.325763, 8.30479, 8.223509, 8.247331, 8.176447, 8.134069, 
    8.106012, 8.086152, 8.088958, 8.094308, 8.121844, 8.147801, 8.167628, 
    8.180913, 8.19402, 8.233806, 8.254919, 8.302357, 8.293777, 8.308313, 
    8.322216, 8.345603, 8.341749, 8.352067, 8.307927, 8.337243, 8.288893, 
    8.302095, 8.197598, 8.158053, 8.141302, 8.126654, 8.091115, 8.115644, 
    8.105968, 8.129003, 8.143668, 8.136412, 8.181276, 8.163811, 8.256171, 
    8.216286, 8.320594, 8.295536, 8.326608, 8.31074, 8.337944, 8.313457, 
    8.355908, 8.365176, 8.358842, 8.383189, 8.312102, 8.339347, 8.136209, 
    8.137392, 8.142904, 8.118695, 8.117215, 8.09508, 8.114773, 8.123171, 
    8.144518, 8.157168, 8.169208, 8.195729, 8.225434, 8.267113, 8.297159, 
    8.317348, 8.304963, 8.315898, 8.303676, 8.297952, 8.361703, 8.325859, 
    8.379684, 8.376698, 8.352313, 8.377034, 8.138223, 8.131415, 8.107821, 
    8.126281, 8.092672, 8.111473, 8.122299, 8.164179, 8.1734, 8.181962, 
    8.198892, 8.220661, 8.258964, 8.292404, 8.323025, 8.320778, 8.321568, 
    8.328422, 8.311457, 8.33121, 8.33453, 8.325853, 8.376298, 8.361861, 
    8.376635, 8.367231, 8.133627, 8.145085, 8.138892, 8.150542, 8.142335, 
    8.178886, 8.189871, 8.241426, 8.220233, 8.25398, 8.223655, 8.229022, 
    8.255088, 8.22529, 8.290561, 8.246269, 8.328689, 8.284301, 8.331476, 
    8.322892, 8.337108, 8.349857, 8.365917, 8.395617, 8.388732, 8.413615, 
    8.162191, 8.177099, 8.175783, 8.191405, 8.202974, 8.228092, 8.26851, 
    8.253292, 8.281245, 8.286867, 8.244404, 8.270457, 8.187087, 8.200513, 
    8.192515, 8.163367, 8.2568, 8.208744, 8.297657, 8.271491, 8.348039, 
    8.309902, 8.384944, 8.417194, 8.447623, 8.483309, 8.185243, 8.175102, 
    8.193264, 8.21845, 8.241867, 8.273086, 8.276284, 8.282146, 8.297341, 
    8.310137, 8.284002, 8.313346, 8.203634, 8.260981, 8.171273, 8.198206, 
    8.216962, 8.208728, 8.251554, 8.261674, 8.302903, 8.281569, 8.409227, 
    8.352556, 8.51055, 8.466164, 8.171562, 8.185206, 8.23284, 8.210148, 
    8.275172, 8.291242, 8.304322, 8.321071, 8.322879, 8.332816, 8.316537, 
    8.332171, 8.273152, 8.299485, 8.227381, 8.244885, 8.236828, 8.228, 
    8.255273, 8.284414, 8.285033, 8.294396, 8.320832, 8.275436, 8.416572, 
    8.329192, 8.200106, 8.226482, 8.230251, 8.220022, 8.28963, 8.264355, 
    8.332573, 8.314091, 8.34439, 8.329323, 8.327108, 8.307793, 8.295786, 
    8.265512, 8.240946, 8.221504, 8.226022, 8.247389, 8.286198, 8.323044, 
    8.314962, 8.342084, 8.270444, 8.300426, 8.288829, 8.319094, 8.252889, 
    8.309252, 8.238533, 8.244713, 8.263853, 8.302465, 8.311021, 8.320171, 
    8.314524, 8.287185, 8.282711, 8.263387, 8.25806, 8.243366, 8.231219, 
    8.242318, 8.253987, 8.287194, 8.317213, 8.350039, 8.358088, 8.396612, 
    8.365246, 8.417061, 8.373001, 8.449383, 8.312521, 8.371699, 8.264724, 
    8.276195, 8.296979, 8.344799, 8.318952, 8.349184, 8.282535, 8.248129, 
    8.239241, 8.222687, 8.239619, 8.238241, 8.254468, 8.24925, 8.288299, 
    8.267305, 8.327054, 8.348945, 8.411006, 8.449235, 8.488283, 8.505569, 
    8.510836, 8.513039,
  12.66455, 12.72001, 12.70921, 12.75408, 12.72917, 12.75858, 12.67577, 
    12.72222, 12.69255, 12.66953, 12.84158, 12.75608, 12.93093, 12.87599, 
    13.01441, 12.92237, 13.03304, 13.01174, 13.07593, 13.05751, 13.13994, 
    13.08444, 13.18286, 13.12667, 13.13544, 13.08261, 12.77324, 12.83091, 
    12.76983, 12.77804, 12.77435, 12.72968, 12.70723, 12.66031, 12.66882, 
    12.70328, 12.78173, 12.75505, 12.82238, 12.82086, 12.89621, 12.86218, 
    12.98945, 12.95316, 13.05828, 13.03177, 13.05703, 13.04936, 13.05713, 
    13.01827, 13.03491, 13.00076, 12.86855, 12.90728, 12.7921, 12.72332, 
    12.67781, 12.64561, 12.65016, 12.65883, 12.70348, 12.7456, 12.77778, 
    12.79935, 12.82064, 12.88529, 12.91962, 12.9968, 12.98283, 13.0065, 
    13.02913, 13.06722, 13.06095, 13.07775, 13.00587, 13.0536, 12.97488, 
    12.99637, 12.82645, 12.76224, 12.73505, 12.71129, 12.65365, 12.69343, 
    12.67774, 12.7151, 12.73889, 12.72712, 12.79994, 12.77158, 12.92165, 
    12.85681, 13.02649, 12.9857, 13.03628, 13.01045, 13.05475, 13.01487, 
    13.08401, 13.09912, 13.08879, 13.12848, 13.01266, 13.05703, 12.72679, 
    12.72871, 12.73765, 12.69838, 12.69598, 12.66008, 12.69201, 12.70564, 
    12.74027, 12.7608, 12.78035, 12.82342, 12.87168, 12.93945, 12.98834, 
    13.02121, 13.00104, 13.01884, 12.99895, 12.98963, 13.09346, 13.03506, 
    13.12277, 13.1179, 13.07816, 13.11845, 12.73005, 12.71901, 12.68074, 
    12.71068, 12.65618, 12.68666, 12.70422, 12.77218, 12.78715, 12.80106, 
    12.82855, 12.86392, 12.92619, 12.9806, 13.03045, 13.02679, 13.02808, 
    13.03924, 13.01161, 13.04378, 13.04919, 13.03505, 13.11725, 13.09372, 
    13.11779, 13.10247, 12.7226, 12.74119, 12.73114, 12.75005, 12.73673, 
    12.79606, 12.8139, 12.89768, 12.86323, 12.91809, 12.86879, 12.87751, 
    12.91989, 12.87145, 12.9776, 12.90555, 13.03967, 12.96741, 13.04421, 
    13.03023, 13.05338, 13.07415, 13.10032, 13.14875, 13.13752, 13.1781, 
    12.76896, 12.79316, 12.79102, 12.81639, 12.83519, 12.876, 12.94172, 
    12.91697, 12.96244, 12.97159, 12.90252, 12.94489, 12.80938, 12.83119, 
    12.8182, 12.77086, 12.92268, 12.84456, 12.98915, 12.94657, 13.07119, 
    13.00908, 13.13134, 13.18394, 13.2336, 13.29188, 12.80638, 12.78992, 
    12.81941, 12.86033, 12.89839, 12.94917, 12.95437, 12.96391, 12.98864, 
    13.00946, 12.96693, 13.01469, 12.83626, 12.92948, 12.7837, 12.82744, 
    12.85791, 12.84453, 12.91414, 12.9306, 12.99769, 12.96297, 13.17094, 
    13.07855, 13.3364, 13.26388, 12.78417, 12.80632, 12.88372, 12.84684, 
    12.95256, 12.97871, 13, 13.02727, 13.03021, 13.04639, 13.01988, 13.04534, 
    12.94927, 12.99212, 12.87485, 12.9033, 12.8902, 12.87585, 12.92019, 
    12.9676, 12.96861, 12.98384, 13.02688, 12.95299, 13.18293, 13.04049, 
    12.83053, 12.87339, 12.87951, 12.86289, 12.97608, 12.93496, 13.046, 
    13.0159, 13.06525, 13.0407, 13.0371, 13.00565, 12.9861, 12.93685, 
    12.8969, 12.8653, 12.87264, 12.90737, 12.9705, 13.03048, 13.01732, 
    13.06149, 12.94487, 12.99366, 12.97478, 13.02405, 12.91632, 13.00802, 
    12.89297, 12.90302, 12.93415, 12.99697, 13.0109, 13.0258, 13.01661, 
    12.97211, 12.96483, 12.93339, 12.92472, 12.90083, 12.88109, 12.89913, 
    12.9181, 12.97212, 13.02098, 13.07445, 13.08756, 13.15037, 13.09923, 
    13.18372, 13.11187, 13.23648, 13.01334, 13.10975, 12.93556, 12.95422, 
    12.98805, 13.06591, 13.02382, 13.07306, 12.96454, 12.90858, 12.89412, 
    12.86722, 12.89474, 12.8925, 12.91888, 12.9104, 12.97392, 12.93976, 
    13.03701, 13.07267, 13.17385, 13.23623, 13.30001, 13.32826, 13.33687, 
    13.34047,
  20.59553, 20.69158, 20.67287, 20.75063, 20.70745, 20.75843, 20.61496, 
    20.69541, 20.64401, 20.60415, 20.90251, 20.75411, 21.05789, 20.96231, 
    21.20334, 21.04299, 21.23583, 21.19868, 21.3107, 21.27854, 21.42258, 
    21.32556, 21.49767, 21.39936, 21.41471, 21.32237, 20.78387, 20.88397, 
    20.77796, 20.79219, 20.7858, 20.70834, 20.66944, 20.5882, 20.60292, 
    20.6626, 20.7986, 20.75231, 20.86917, 20.86652, 20.99748, 20.93832, 
    21.15982, 21.09659, 21.27988, 21.23362, 21.27771, 21.26432, 21.27788, 
    21.21008, 21.2391, 21.17954, 20.94938, 21.01673, 20.8166, 20.69731, 
    20.61848, 20.56276, 20.57063, 20.58563, 20.66295, 20.73593, 20.79175, 
    20.82918, 20.86614, 20.97848, 21.0382, 21.17263, 21.14829, 21.18954, 
    21.22902, 21.2955, 21.28454, 21.31389, 21.18845, 21.27173, 21.13444, 
    21.17189, 20.87623, 20.76479, 20.71765, 20.67646, 20.57668, 20.64553, 
    20.61836, 20.68306, 20.7243, 20.70389, 20.83021, 20.781, 21.04175, 
    20.92898, 21.22441, 21.15329, 21.2415, 21.19643, 21.27372, 21.20415, 
    21.32483, 21.35121, 21.33318, 21.40253, 21.2003, 21.27771, 20.70332, 
    20.70665, 20.72215, 20.6541, 20.64994, 20.5878, 20.64308, 20.66668, 
    20.72669, 20.76229, 20.7962, 20.87096, 20.95482, 21.07273, 21.15789, 
    21.2152, 21.18003, 21.21107, 21.17638, 21.16014, 21.34132, 21.23937, 
    21.39254, 21.38403, 21.31459, 21.38499, 20.70899, 20.68985, 20.62356, 
    20.67542, 20.58105, 20.63381, 20.66423, 20.78203, 20.80801, 20.83214, 
    20.87988, 20.94134, 21.04965, 21.1444, 21.23132, 21.22494, 21.22718, 
    21.24665, 21.19846, 21.25458, 21.26401, 21.23935, 21.38289, 21.34177, 
    21.38385, 21.35707, 20.69607, 20.72829, 20.71087, 20.74364, 20.72055, 
    20.82347, 20.85443, 21.00003, 20.94013, 21.03554, 20.9498, 20.96496, 
    21.03868, 20.95442, 21.13917, 21.01373, 21.24741, 21.12143, 21.25533, 
    21.23094, 21.27134, 21.30761, 21.35332, 21.43797, 21.41833, 21.48934, 
    20.77644, 20.81843, 20.81472, 20.85876, 20.8914, 20.96234, 21.07668, 
    21.0336, 21.11276, 21.1287, 21.00845, 21.0822, 20.84659, 20.88446, 
    20.86189, 20.77975, 21.04353, 20.90769, 21.1593, 21.08513, 21.30243, 
    21.19405, 21.40754, 21.49956, 21.58656, 21.68877, 20.84138, 20.81281, 
    20.864, 20.93509, 21.00128, 21.08964, 21.09871, 21.11532, 21.15841, 
    21.19472, 21.12058, 21.20383, 20.89326, 21.05536, 20.80202, 20.87795, 
    20.93089, 20.90764, 21.02868, 21.05732, 21.17419, 21.11368, 21.47681, 
    21.31528, 21.76694, 21.63964, 20.80283, 20.84128, 20.97575, 20.91165, 
    21.09555, 21.14111, 21.17821, 21.22577, 21.2309, 21.25914, 21.21289, 
    21.25731, 21.08983, 21.16449, 20.96033, 21.00982, 20.98703, 20.96207, 
    21.03921, 21.12175, 21.1235, 21.15005, 21.22509, 21.0963, 21.49779, 
    21.24884, 20.88331, 20.95779, 20.96844, 20.93954, 21.13653, 21.06491, 
    21.25845, 21.20594, 21.29205, 21.24921, 21.24292, 21.18806, 21.15399, 
    21.06819, 20.99867, 20.94372, 20.95648, 21.0169, 21.1268, 21.23137, 
    21.20842, 21.28549, 21.08216, 21.16716, 21.13426, 21.22015, 21.03246, 
    21.1922, 20.99185, 21.00933, 21.06349, 21.17294, 21.19723, 21.22321, 
    21.20717, 21.1296, 21.11692, 21.06217, 21.04709, 21.00552, 20.97117, 
    21.00255, 21.03557, 21.12963, 21.21481, 21.30812, 21.33103, 21.44081, 
    21.35141, 21.49918, 21.3735, 21.59159, 21.20149, 21.36979, 21.06596, 
    21.09845, 21.15738, 21.29321, 21.21975, 21.30569, 21.11642, 21.01899, 
    20.99385, 20.94706, 20.99492, 20.99102, 21.03693, 21.02216, 21.13276, 
    21.07327, 21.24277, 21.30501, 21.48189, 21.59117, 21.70304, 21.75264, 
    21.76776, 21.77409,
  34.63897, 34.81973, 34.78447, 34.93106, 34.84963, 34.94577, 34.6755, 
    34.82694, 34.73015, 34.65517, 35.21813, 34.93762, 35.51293, 35.33146, 
    35.78991, 35.48461, 35.85193, 35.78102, 35.99502, 35.93352, 36.20935, 
    36.02346, 36.35355, 36.16482, 36.19426, 36.01735, 34.99379, 35.18303, 
    34.98262, 35.00951, 34.99744, 34.85131, 34.77802, 34.6252, 34.65287, 
    34.76514, 35.0216, 34.93423, 35.15501, 35.15001, 35.39817, 35.28596, 
    35.70693, 35.58653, 35.93608, 35.8477, 35.93193, 35.90635, 35.93226, 
    35.80277, 35.85817, 35.74452, 35.30694, 35.43473, 35.05561, 34.83052, 
    34.68213, 34.57739, 34.59217, 34.62037, 34.7658, 34.90333, 35.00867, 
    35.0794, 35.14928, 35.36213, 35.47551, 35.73136, 35.68497, 35.7636, 
    35.83892, 35.96595, 35.945, 36.00113, 35.76151, 35.9205, 35.65859, 
    35.72994, 35.16838, 34.95776, 34.86885, 34.79125, 34.60354, 34.73301, 
    34.68189, 34.80368, 34.8814, 34.84293, 35.08133, 34.98837, 35.48225, 
    35.26827, 35.83013, 35.69448, 35.86275, 35.77674, 35.92431, 35.79145, 
    36.02205, 36.07256, 36.03803, 36.17091, 35.78411, 35.93193, 34.84185, 
    34.84812, 34.87735, 34.74914, 34.74132, 34.62444, 34.7284, 34.77282, 
    34.88591, 34.95306, 35.01707, 35.15841, 35.31726, 35.54113, 35.70325, 
    35.81254, 35.74546, 35.80467, 35.73849, 35.70753, 36.05362, 35.85868, 
    36.15175, 36.13544, 36.00246, 36.13728, 34.85253, 34.81646, 34.69168, 
    34.78928, 34.61175, 34.71097, 34.76821, 34.99032, 35.03938, 35.08498, 
    35.17529, 35.29169, 35.49726, 35.67756, 35.84331, 35.83113, 35.83541, 
    35.8726, 35.78061, 35.88773, 35.90576, 35.85865, 36.13326, 36.05449, 
    36.13509, 36.08377, 34.82817, 34.88892, 34.85608, 34.91788, 34.87433, 
    35.0686, 35.12715, 35.40302, 35.2894, 35.47046, 35.30773, 35.33649, 
    35.47642, 35.31649, 35.66759, 35.42902, 35.87404, 35.6338, 35.88918, 
    35.84259, 35.91977, 35.9891, 36.0766, 36.2389, 36.20121, 36.33756, 
    34.97976, 35.05908, 35.05207, 35.13533, 35.1971, 35.3315, 35.54866, 
    35.46676, 35.61731, 35.64765, 35.41901, 35.55915, 35.1123, 35.18395, 
    35.14126, 34.98601, 35.48563, 35.22794, 35.70594, 35.56472, 35.97921, 
    35.7722, 36.1805, 36.3572, 36.52462, 36.72183, 35.10247, 35.04845, 
    35.14525, 35.27985, 35.40538, 35.57331, 35.59055, 35.62217, 35.70424, 
    35.77346, 35.63218, 35.79085, 35.20062, 35.50812, 35.02806, 35.17163, 
    35.27189, 35.22785, 35.45742, 35.51185, 35.73432, 35.61905, 36.31348, 
    36.00379, 36.87302, 36.62696, 35.0296, 35.10228, 35.35695, 35.23544, 
    35.58456, 35.67128, 35.74199, 35.83271, 35.84252, 35.89645, 35.80814, 
    35.89295, 35.57367, 35.71583, 35.32769, 35.42159, 35.37835, 35.33101, 
    35.47742, 35.63441, 35.63775, 35.68832, 35.83142, 35.58598, 36.35378, 
    35.87677, 35.18178, 35.32288, 35.34307, 35.28827, 35.66257, 35.52628, 
    35.89513, 35.79488, 35.95935, 35.87749, 35.86547, 35.76077, 35.69583, 
    35.53252, 35.40044, 35.29621, 35.32041, 35.43504, 35.64404, 35.84341, 
    35.7996, 35.94681, 35.55907, 35.72091, 35.65824, 35.82199, 35.4646, 
    35.76867, 35.38749, 35.42067, 35.52358, 35.73195, 35.77826, 35.82784, 
    35.79723, 35.64936, 35.62521, 35.52107, 35.4924, 35.41344, 35.34827, 
    35.40781, 35.4705, 35.64942, 35.8118, 35.99009, 36.03392, 36.24434, 
    36.07294, 36.35647, 36.11525, 36.53432, 35.78638, 36.10815, 35.52827, 
    35.59007, 35.70228, 35.96158, 35.82122, 35.98544, 35.62427, 35.43901, 
    35.39129, 35.30254, 35.39332, 35.38593, 35.47309, 35.44504, 35.65538, 
    35.54217, 35.86517, 35.98413, 36.32324, 36.53351, 36.7494, 36.84533, 
    36.87461, 36.88686,
  60.67812, 61.07083, 60.99409, 61.31372, 61.13599, 61.34588, 60.75732, 
    61.08654, 60.87596, 60.71325, 61.9436, 61.32805, 62.59597, 62.19373, 
    63.21417, 62.53306, 63.35332, 63.19427, 63.67535, 63.53676, 64.1604, 
    63.73951, 64.48857, 64.05934, 64.12612, 63.72573, 61.45091, 61.86631, 
    61.42648, 61.48533, 61.4589, 61.13966, 60.98005, 60.64828, 60.70824, 
    60.95203, 61.51183, 61.32064, 61.80466, 61.79365, 62.34135, 62.09321, 
    63.02843, 62.75974, 63.54253, 63.34382, 63.53318, 63.47563, 63.53393, 
    63.243, 63.36732, 63.11252, 62.13954, 62.42237, 61.58636, 61.09434, 
    60.77169, 60.54478, 60.57676, 60.63782, 60.95346, 61.25314, 61.48349, 
    61.63854, 61.79206, 62.26156, 62.51286, 63.08306, 62.97934, 63.15522, 
    63.32412, 63.60981, 63.5626, 63.68912, 63.15054, 63.50746, 62.92043, 
    63.0799, 61.83408, 61.3721, 61.17791, 61.00883, 60.60137, 60.88219, 
    60.77119, 61.03589, 61.20528, 61.12138, 61.64279, 61.43905, 62.52781, 
    62.05416, 63.30437, 63.0006, 63.37762, 63.18466, 63.51603, 63.21764, 
    63.73632, 63.85044, 63.77242, 64.07315, 63.20118, 63.53319, 61.11904, 
    61.13271, 61.19645, 60.91724, 60.90023, 60.64664, 60.87217, 60.96872, 
    61.21512, 61.36181, 61.5019, 61.81213, 62.16233, 62.65868, 63.0202, 
    63.26491, 63.11462, 63.24727, 63.09903, 63.02978, 63.80764, 63.36849, 
    64.02972, 63.99275, 63.69214, 63.99691, 61.14231, 61.06372, 60.79243, 
    61.00453, 60.61915, 60.8343, 60.95869, 61.44332, 61.55079, 61.65081, 
    61.84927, 62.10587, 62.56117, 62.96279, 63.33397, 63.30662, 63.31624, 
    63.39974, 63.19334, 63.43375, 63.4743, 63.36842, 63.98781, 63.80959, 
    63.99197, 63.8758, 61.08924, 61.22169, 61.15005, 61.28492, 61.18985, 
    61.61485, 61.7434, 62.35209, 62.1008, 62.50164, 62.14127, 62.20483, 
    62.51487, 62.16063, 62.94054, 62.40971, 63.40299, 62.8651, 63.43701, 
    63.33235, 63.50581, 63.66199, 63.85958, 64.22751, 64.14191, 64.4521, 
    61.4202, 61.59397, 61.57861, 61.76139, 61.89728, 62.19381, 62.67543, 
    62.49343, 62.82833, 62.89601, 62.38752, 62.69877, 61.71079, 61.86833, 
    61.77442, 61.43389, 62.53532, 61.96521, 63.02622, 62.71117, 63.63968, 
    63.17449, 64.0949, 64.49689, 64.87986, 65.33361, 61.68919, 61.57065, 
    61.7832, 62.07972, 62.35733, 62.7303, 62.7687, 62.83917, 63.02241, 
    63.17733, 62.86151, 63.21629, 61.90504, 62.58529, 61.52598, 61.84122, 
    62.06215, 61.96502, 62.4727, 62.59358, 63.08968, 62.83222, 64.39722, 
    63.69513, 65.68346, 65.11497, 61.52935, 61.68877, 62.2501, 61.98175, 
    62.75534, 62.94876, 63.10686, 63.31018, 63.33218, 63.45336, 63.25504, 
    63.44549, 62.7311, 63.04832, 62.18539, 62.39325, 62.29744, 62.19271, 
    62.51709, 62.86647, 62.87393, 62.98683, 63.30727, 62.75852, 64.48909, 
    63.40913, 61.86354, 62.17475, 62.2194, 62.09831, 62.92932, 62.62565, 
    63.45039, 63.22533, 63.59494, 63.41073, 63.38372, 63.14891, 63.00361, 
    62.63952, 62.34637, 62.11584, 62.16929, 62.42305, 62.88795, 63.3342, 
    63.23591, 63.56669, 62.6986, 63.0597, 62.91965, 63.28613, 62.48862, 
    63.16659, 62.31769, 62.39119, 62.61966, 63.08437, 63.18806, 63.29924, 
    63.23058, 62.89984, 62.84597, 62.61407, 62.55037, 62.37517, 62.23088, 
    62.3627, 62.50174, 62.89996, 63.26326, 63.66423, 63.76313, 64.23988, 
    63.8513, 64.49522, 63.94703, 64.90211, 63.20626, 63.93095, 62.63008, 
    62.76763, 63.01803, 63.59995, 63.2844, 63.65373, 62.84385, 62.43187, 
    62.3261, 62.12981, 62.3306, 62.31422, 62.50748, 62.44524, 62.91327, 
    62.66099, 63.38305, 63.65079, 64.41946, 64.90024, 65.39728, 65.61927, 
    65.68715, 65.71558,
  116.3177, 117.5456, 117.3041, 118.3151, 117.7513, 118.4176, 116.5637, 
    117.5951, 116.9338, 116.4267, 120.3481, 118.3608, 122.5137, 121.171, 
    124.6257, 122.3021, 125.1096, 124.5568, 126.2417, 125.7524, 127.9808, 
    126.4694, 129.1813, 127.615, 127.8565, 126.4205, 118.7533, 120.0957, 
    118.6751, 118.8636, 118.7789, 117.7629, 117.26, 116.2252, 116.4112, 
    117.1721, 118.9486, 118.3372, 119.895, 119.8591, 121.6609, 120.8392, 
    123.9848, 123.0673, 125.7727, 125.0765, 125.7398, 125.5376, 125.7424, 
    124.7257, 125.1585, 124.2743, 120.992, 121.9312, 119.1884, 117.6198, 
    116.6085, 115.9052, 116.004, 116.1928, 117.1766, 118.1225, 118.8577, 
    119.3567, 119.854, 121.3957, 122.2342, 124.1727, 123.8163, 124.4217, 
    125.0078, 126.0099, 125.8434, 126.2906, 124.4055, 125.6493, 123.6146, 
    124.1618, 119.9907, 118.5013, 117.8839, 117.3504, 116.08, 116.9533, 
    116.6069, 117.4356, 117.9706, 117.7051, 119.3704, 118.7153, 122.2844, 
    120.7108, 124.939, 123.8892, 125.1944, 124.5235, 125.6795, 124.6378, 
    126.4581, 126.8647, 126.5865, 127.6649, 124.5807, 125.7398, 117.6977, 
    117.7409, 117.9426, 117.063, 117.0098, 116.2201, 116.922, 117.2244, 
    118.0018, 118.4685, 118.9168, 119.9193, 121.0672, 122.7252, 123.9565, 
    124.8018, 124.2815, 124.7405, 124.2277, 123.9894, 126.712, 125.1625, 
    127.5082, 127.375, 126.3013, 127.39, 117.7713, 117.5232, 116.6731, 
    117.3369, 116.135, 116.8037, 117.193, 118.729, 119.0739, 119.3963, 
    120.0402, 120.8809, 122.3965, 123.7596, 125.0421, 124.9468, 124.9804, 
    125.2717, 124.5536, 125.3907, 125.5329, 125.1623, 127.3572, 126.7189, 
    127.3722, 126.9554, 117.6037, 118.0227, 117.7958, 118.2235, 117.9217, 
    119.2802, 119.696, 121.6967, 120.8642, 122.1966, 120.9977, 121.2077, 
    122.241, 121.0616, 123.6834, 121.8889, 125.2831, 123.4257, 125.4021, 
    125.0365, 125.6435, 126.1945, 126.8974, 128.2247, 127.9137, 129.0469, 
    118.655, 119.2129, 119.1634, 119.7544, 120.1967, 121.1713, 122.7818, 
    122.1691, 123.3005, 123.5312, 121.8148, 122.8607, 119.5903, 120.1023, 
    119.7967, 118.6988, 122.3096, 120.4189, 123.9772, 122.9027, 126.1155, 
    124.4883, 127.7435, 129.212, 130.6391, 132.3671, 119.5204, 119.1378, 
    119.8252, 120.7948, 121.7141, 122.9675, 123.0977, 123.3373, 123.9641, 
    124.4982, 123.4135, 124.6331, 120.2221, 122.4777, 118.9941, 120.0139, 
    120.737, 120.4182, 122.0996, 122.5056, 124.1955, 123.3137, 128.8451, 
    126.3119, 133.7281, 131.5293, 119.0049, 119.519, 121.3577, 120.4731, 
    123.0524, 123.7116, 124.2547, 124.9592, 125.0359, 125.4594, 124.7675, 
    125.4319, 122.9702, 124.0532, 121.1434, 121.8339, 121.5149, 121.1676, 
    122.2484, 123.4304, 123.4558, 123.842, 124.9491, 123.0632, 129.1832, 
    125.3046, 120.0867, 121.1082, 121.256, 120.856, 123.645, 122.6137, 
    125.4491, 124.6644, 125.9574, 125.3102, 125.2157, 124.3999, 123.8996, 
    122.6605, 121.6777, 120.9138, 121.0902, 121.9335, 123.5037, 125.0429, 
    124.7011, 125.8578, 122.8601, 124.0923, 123.612, 124.8756, 122.153, 
    124.461, 121.5822, 121.8271, 122.5935, 124.1772, 124.5353, 124.9212, 
    124.6826, 123.5443, 123.3605, 122.5746, 122.3602, 121.7736, 121.294, 
    121.7321, 122.1969, 123.5447, 124.7961, 126.2024, 126.5534, 128.2697, 
    126.8678, 129.2058, 127.2107, 130.7228, 124.5983, 127.153, 122.6286, 
    123.0941, 123.9491, 125.9751, 124.8695, 126.1652, 123.3533, 121.963, 
    121.6102, 120.9599, 121.6252, 121.5707, 122.2162, 122.0077, 123.5901, 
    122.733, 125.2134, 126.1548, 128.9268, 130.7158, 132.6128, 133.4764, 
    133.7426, 133.8543,
  366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466,
  603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILPSI =
  -0.02027925, -0.01994774, -0.02001173, -0.01974766, -0.01989369, 
    -0.01972144, -0.02021158, -0.01993468, -0.02011098, -0.02024919, 
    -0.01924578, -0.01973597, -0.01875059, -0.01905304, -0.0183031, 
    -0.01879729, -0.01820517, -0.01831719, -0.01798235, -0.01807759, 
    -0.01765646, -0.01793857, -0.0174424, -0.01772341, -0.01767912, 
    -0.01794796, -0.01963629, -0.01930608, -0.01965603, -0.01960853, 
    -0.01962983, -0.01989065, -0.02002348, -0.02030485, -0.02025346, 
    -0.02004696, -0.01958721, -0.01974201, -0.01935442, -0.01936308, 
    -0.01894098, -0.01913005, -0.0184354, -0.01863003, -0.01807361, 
    -0.01821183, -0.01808007, -0.01811992, -0.01807955, -0.01828273, 
    -0.01819538, -0.01837528, -0.01909448, -0.01888, -0.01952747, 
    -0.01992821, -0.02019934, -0.02039412, -0.02036646, -0.02031384, 
    -0.02004576, -0.01979721, -0.01961, -0.01948584, -0.01936433, 
    -0.01900139, -0.01881234, -0.0183963, -0.01847067, -0.01834489, 
    -0.01822564, -0.01802727, -0.01805976, -0.01797293, -0.01834822, 
    -0.01809786, -0.01851317, -0.01839856, -0.01933132, -0.01970012, 
    -0.01985907, -0.01999941, -0.02034522, -0.02010573, -0.02019977, 
    -0.01997682, -0.01983652, -0.01990579, -0.01948246, -0.01964587, 
    -0.0188012, -0.01916013, -0.01823951, -0.01845538, -0.01818817, 
    -0.018324, -0.01809193, -0.01830065, -0.01794074, -0.01786338, 
    -0.0179162, -0.01771424, -0.01831229, -0.01808006, -0.01990772, 
    -0.01989641, -0.01984379, -0.0200762, -0.02009051, -0.02030626, 
    -0.02011418, -0.02003297, -0.01982843, -0.01970848, -0.01959519, 
    -0.01934855, -0.01907703, -0.01870425, -0.0184413, -0.01826727, 
    -0.01837378, -0.01827971, -0.0183849, -0.01843443, -0.01789232, 
    -0.01819456, -0.01774313, -0.0177678, -0.01797087, -0.01776502, 
    -0.01988847, -0.01995365, -0.02018171, -0.020003, -0.02032991, 
    -0.0201462, -0.02004137, -0.01964241, -0.01955594, -0.01947608, 
    -0.01931941, -0.01912033, -0.0187764, -0.01848259, -0.01821873, 
    -0.01823793, -0.01823117, -0.01817273, -0.01831784, -0.01814902, 
    -0.01812084, -0.0181946, -0.0177711, -0.017891, -0.01776832, -0.01784628, 
    -0.01993244, -0.01982302, -0.01988207, -0.01977119, -0.01984922, 
    -0.01950472, -0.01940269, -0.01893288, -0.01912422, -0.0188207, 
    -0.01909316, -0.01904457, -0.01881084, -0.01907833, -0.01849864, 
    -0.0188895, -0.01817046, -0.01855325, -0.01814676, -0.01821987, 
    -0.018099, -0.01799148, -0.01785721, -0.01761227, -0.01766867, 
    -0.01746595, -0.01966111, -0.01952138, -0.01953366, -0.0193885, 
    -0.01928188, -0.01905297, -0.01869191, -0.01882682, -0.01857997, 
    -0.01853083, -0.01890619, -0.01867474, -0.01942848, -0.01930449, 
    -0.01937823, -0.01965004, -0.01879561, -0.01922898, -0.01843699, 
    -0.01866563, -0.01800677, -0.01833121, -0.0176998, -0.01743704, 
    -0.0171937, -0.01691387, -0.0194456, -0.01954002, -0.01937131, 
    -0.01914044, -0.01892892, -0.0186516, -0.01862348, -0.01857209, 
    -0.01843972, -0.0183292, -0.01855586, -0.01830161, -0.01927582, 
    -0.0187585, -0.01957583, -0.01932573, -0.01915397, -0.01922913, 
    -0.01884231, -0.01875236, -0.01839157, -0.01857715, -0.01750148, 
    -0.01796883, -0.0167042, -0.01704757, -0.01957313, -0.01944593, 
    -0.0190101, -0.01921614, -0.01863325, -0.01849271, -0.01837932, 
    -0.01823543, -0.01821998, -0.01813538, -0.01827423, -0.01814085, 
    -0.01865101, -0.01842114, -0.0190594, -0.01890188, -0.01897418, 
    -0.01905381, -0.01880919, -0.01855226, -0.01854684, -0.01846528, 
    -0.01823747, -0.01863093, -0.01744207, -0.01816618, -0.01930824, 
    -0.01906754, -0.01903346, -0.01912613, -0.01850674, -0.01872863, 
    -0.01813745, -0.01829521, -0.01803749, -0.01816506, -0.01818391, 
    -0.01834938, -0.01845321, -0.01871839, -0.01893719, -0.01911267, 
    -0.01907171, -0.01887949, -0.01853667, -0.01821857, -0.01828774, 
    -0.01805694, -0.01867487, -0.018413, -0.01851373, -0.01825233, 
    -0.01883041, -0.01833682, -0.01895886, -0.01890342, -0.01873306, 
    -0.01839536, -0.01832159, -0.01824312, -0.0182915, -0.01852806, 
    -0.01856715, -0.01873719, -0.01878442, -0.01891548, -0.01902471, 
    -0.01892488, -0.01882063, -0.01852798, -0.01826844, -0.01798995, 
    -0.01792251, -0.01760415, -0.0178628, -0.01743812, -0.0177984, 
    -0.01717976, -0.0183087, -0.01780918, -0.01872536, -0.01862426, 
    -0.01844286, -0.01803404, -0.01825355, -0.01799714, -0.01856869, 
    -0.01887288, -0.01895249, -0.01910194, -0.01894909, -0.01896148, 
    -0.01881635, -0.01886285, -0.01851835, -0.01870255, -0.01818438, 
    -0.01799916, -0.01748706, -0.01718093, -0.01687533, -0.01674228, 
    -0.01670201, -0.01668521,
  -0.05400472, -0.05296151, -0.05316266, -0.05233337, -0.05279174, 
    -0.05225114, -0.05379153, -0.05292049, -0.05347484, -0.05390999, 
    -0.05076257, -0.05229671, -0.04921966, -0.05016121, -0.04783148, 
    -0.04936488, -0.04752846, -0.0478751, -0.04684005, -0.04713414, 
    -0.0458359, -0.04670498, -0.04517806, -0.04604194, -0.0459056, 
    -0.04673393, -0.05198419, -0.05095092, -0.05204607, -0.05189721, 
    -0.05196397, -0.05278219, -0.05319959, -0.05408542, -0.05392347, 
    -0.05327345, -0.05183041, -0.05231566, -0.05110202, -0.0511291, 
    -0.04981206, -0.05040139, -0.0482413, -0.04884512, -0.04712183, 
    -0.04754905, -0.04714178, -0.0472649, -0.04714018, -0.04776842, 
    -0.04749817, -0.048055, -0.05029044, -0.04962223, -0.05164335, 
    -0.05290014, -0.053753, -0.05436689, -0.05427966, -0.05411374, 
    -0.05326967, -0.05248883, -0.05190184, -0.05151305, -0.051133, 
    -0.05000024, -0.0494117, -0.04812012, -0.04835062, -0.04796088, 
    -0.04759178, -0.04697872, -0.04707906, -0.046811, -0.04797119, 
    -0.04719674, -0.04848243, -0.04812713, -0.05102981, -0.05218429, 
    -0.05268299, -0.05312392, -0.05421267, -0.0534583, -0.05375434, 
    -0.05305294, -0.05261222, -0.05282972, -0.05150247, -0.05201422, 
    -0.04937704, -0.05049522, -0.04763468, -0.04830323, -0.0474759, 
    -0.0478962, -0.04717841, -0.04782389, -0.04671167, -0.0464731, 
    -0.04663599, -0.04601369, -0.04785994, -0.04714175, -0.05283581, 
    -0.05280027, -0.05263505, -0.05336539, -0.05341044, -0.05408985, 
    -0.05348491, -0.05322943, -0.05258682, -0.0522105, -0.05185543, 
    -0.05108368, -0.05023602, -0.04907565, -0.04825959, -0.0477206, 
    -0.04805036, -0.0477591, -0.04808481, -0.04823829, -0.04656232, 
    -0.04749564, -0.04610265, -0.0461786, -0.04680463, -0.04617004, 
    -0.05277533, -0.05298011, -0.05369748, -0.05313521, -0.05416439, 
    -0.05358569, -0.05325587, -0.05200339, -0.05173249, -0.0514825, 
    -0.0509926, -0.05037104, -0.04929992, -0.0483876, -0.04757041, 
    -0.0476298, -0.04760888, -0.04742814, -0.04787713, -0.04735485, 
    -0.04726776, -0.04749579, -0.04618878, -0.04655825, -0.04618022, 
    -0.04642039, -0.05291346, -0.05256985, -0.05275523, -0.05240719, 
    -0.0526521, -0.05157214, -0.05125293, -0.04978683, -0.05038318, 
    -0.0494377, -0.0502863, -0.0501348, -0.04940702, -0.05024008, 
    -0.04843737, -0.04965179, -0.04742113, -0.04860676, -0.04734785, 
    -0.04757392, -0.04720028, -0.04686824, -0.0464541, -0.04569999, 
    -0.04587347, -0.04525035, -0.052062, -0.05162429, -0.05166275, 
    -0.05120854, -0.05087532, -0.05016102, -0.04903733, -0.04945675, 
    -0.04868972, -0.04853724, -0.04970374, -0.04898399, -0.05133358, 
    -0.05094598, -0.05117644, -0.05202729, -0.04935967, -0.05071013, 
    -0.0482462, -0.04895568, -0.04691542, -0.04791851, -0.04596925, 
    -0.0451616, -0.04441552, -0.04355986, -0.05138713, -0.05168267, 
    -0.05115483, -0.05043377, -0.04977453, -0.04891208, -0.04882477, 
    -0.04866525, -0.04825468, -0.04791228, -0.04861486, -0.04782686, 
    -0.05085639, -0.04924429, -0.0517948, -0.05101232, -0.050476, -0.0507106, 
    -0.04950494, -0.0492252, -0.04810547, -0.04868094, -0.04535947, 
    -0.04679833, -0.0429203, -0.04396839, -0.05178633, -0.05138818, 
    -0.05002738, -0.05067005, -0.04885511, -0.04841897, -0.04806751, 
    -0.04762205, -0.04757427, -0.0473127, -0.04774213, -0.04732961, 
    -0.04891026, -0.04819711, -0.05018106, -0.04969032, -0.04991547, 
    -0.05016363, -0.0494019, -0.04860369, -0.0485869, -0.04833392, 
    -0.04762835, -0.0488479, -0.04517701, -0.04740787, -0.05095769, 
    -0.05020641, -0.0501002, -0.05038915, -0.0484625, -0.04915142, 
    -0.04731907, -0.04780707, -0.04701029, -0.04740444, -0.04746272, 
    -0.04797479, -0.04829651, -0.04911959, -0.04980025, -0.05034715, 
    -0.05021943, -0.04962062, -0.04855534, -0.0475699, -0.04778393, 
    -0.04707034, -0.04898436, -0.04817187, -0.04848416, -0.04767436, 
    -0.04946792, -0.04793586, -0.04986774, -0.04969514, -0.0491652, 
    -0.04811721, -0.04788873, -0.04764584, -0.04779558, -0.04852863, 
    -0.04864991, -0.04917804, -0.04932487, -0.04973267, -0.05007294, 
    -0.04976192, -0.04943748, -0.04852837, -0.04772419, -0.04686351, 
    -0.04665545, -0.045675, -0.04647131, -0.04516489, -0.04627284, 
    -0.04437285, -0.0478488, -0.04630607, -0.04914127, -0.0488272, 
    -0.04826441, -0.04699963, -0.04767814, -0.0468857, -0.04865468, 
    -0.04960005, -0.04984793, -0.0503137, -0.04983734, -0.04987591, 
    -0.04942417, -0.04956887, -0.04849849, -0.04907038, -0.04746415, 
    -0.04689192, -0.04531519, -0.04437644, -0.04344219, -0.04303636, 
    -0.04291365, -0.04286246,
  -0.07871422, -0.07706323, -0.07738139, -0.07607025, -0.07679477, 
    -0.07594033, -0.07837664, -0.07699836, -0.07787535, -0.07856421, 
    -0.07359091, -0.07601232, -0.071161, -0.07264318, -0.06897949, 
    -0.07138947, -0.06850391, -0.06904797, -0.06742429, -0.06788536, 
    -0.06585159, -0.0672126, -0.06482265, -0.06617408, -0.06596068, 
    -0.06725796, -0.07551863, -0.07388791, -0.07561637, -0.07538126, 
    -0.0754867, -0.07677967, -0.07743981, -0.07884203, -0.07858555, 
    -0.07755666, -0.07527579, -0.07604226, -0.07412623, -0.07416894, 
    -0.07209331, -0.0730216, -0.06962305, -0.07057196, -0.06786605, 
    -0.06853621, -0.06789735, -0.06809043, -0.06789484, -0.06888051, 
    -0.06845637, -0.06933043, -0.07284677, -0.07179447, -0.07498045, 
    -0.07696617, -0.07831563, -0.07928794, -0.07914972, -0.0788869, 
    -0.07755069, -0.07631592, -0.07538859, -0.07477478, -0.07417509, 
    -0.07238965, -0.07146313, -0.06943271, -0.06979479, -0.06918265, 
    -0.06860327, -0.06764167, -0.06779899, -0.06737875, -0.06919883, 
    -0.06798354, -0.07000188, -0.06944371, -0.07401233, -0.07583472, 
    -0.07662284, -0.07732011, -0.07904361, -0.07784916, -0.07831776, 
    -0.07720783, -0.07651095, -0.07685482, -0.07475808, -0.07556607, 
    -0.0714086, -0.07316948, -0.06867059, -0.06972032, -0.06842145, 
    -0.06908108, -0.06795479, -0.06896758, -0.06722309, -0.06684929, 
    -0.06710448, -0.06612986, -0.06902417, -0.0678973, -0.07686445, 
    -0.07680825, -0.07654704, -0.07770214, -0.07777342, -0.07884905, 
    -0.07789126, -0.07748702, -0.07647081, -0.07587612, -0.0753153, 
    -0.07409729, -0.07276104, -0.07093447, -0.06965177, -0.06880543, 
    -0.06932315, -0.06886587, -0.06937724, -0.06961831, -0.06698906, 
    -0.0684524, -0.06626914, -0.06638805, -0.06736878, -0.06637464, 
    -0.07676882, -0.07709263, -0.07822774, -0.07733796, -0.07896712, 
    -0.07805078, -0.07752884, -0.07554896, -0.07512117, -0.07472657, 
    -0.07395365, -0.07297378, -0.07128726, -0.06985288, -0.06856973, 
    -0.06866293, -0.0686301, -0.0683465, -0.06905115, -0.06823154, 
    -0.06809492, -0.06845264, -0.06640399, -0.06698269, -0.06639057, 
    -0.06676671, -0.07698724, -0.07644399, -0.07673703, -0.0761869, 
    -0.076574, -0.07486805, -0.0743643, -0.07205359, -0.07299291, 
    -0.07150405, -0.07284026, -0.07260158, -0.07145578, -0.07276743, 
    -0.06993107, -0.071841, -0.0683355, -0.07019726, -0.06822055, 
    -0.06857523, -0.06798908, -0.06746848, -0.06681952, -0.06563892, 
    -0.06591038, -0.06493566, -0.07564154, -0.07495037, -0.07501107, 
    -0.07429426, -0.07376869, -0.07264287, -0.0708742, -0.07153402, 
    -0.07032766, -0.070088, -0.07192276, -0.07079032, -0.07449156, 
    -0.07388011, -0.07424362, -0.07558671, -0.07138126, -0.07350823, 
    -0.06963075, -0.0707458, -0.06754243, -0.06911613, -0.0660603, 
    -0.06479692, -0.06363132, -0.06229629, -0.07457605, -0.07504252, 
    -0.07420953, -0.07307262, -0.07203422, -0.07067724, -0.07053997, 
    -0.07028919, -0.06964406, -0.06910634, -0.07020999, -0.06897224, 
    -0.07373884, -0.07119974, -0.07521956, -0.07398475, -0.07313918, 
    -0.07350898, -0.07160987, -0.0711697, -0.06940971, -0.07031386, 
    -0.06510629, -0.0673589, -0.0612997, -0.06293346, -0.07520619, 
    -0.0745777, -0.07243238, -0.07344504, -0.07058766, -0.06990215, 
    -0.06935008, -0.06865078, -0.0685758, -0.06816541, -0.06883924, 
    -0.06819194, -0.07067438, -0.06955363, -0.07267445, -0.07190165, 
    -0.07225614, -0.07264699, -0.07144771, -0.07019246, -0.07016606, 
    -0.06976855, -0.06866066, -0.07057633, -0.06482102, -0.06831471, 
    -0.07389858, -0.07271439, -0.07254707, -0.07300232, -0.06997056, 
    -0.07105365, -0.06817541, -0.06894117, -0.06769116, -0.06830932, 
    -0.06840076, -0.06920448, -0.06970978, -0.07100358, -0.07207472, 
    -0.07293613, -0.07273489, -0.07179195, -0.07011646, -0.06856894, 
    -0.06890484, -0.06778533, -0.07079091, -0.06951399, -0.0700046, 
    -0.06873287, -0.07155161, -0.06914337, -0.07218099, -0.07190923, 
    -0.07107533, -0.06942814, -0.06906936, -0.0686881, -0.06892314, 
    -0.07007449, -0.07026509, -0.07109552, -0.07132651, -0.07196832, 
    -0.07250413, -0.07201438, -0.0715037, -0.07007407, -0.06881107, 
    -0.06746107, -0.06713498, -0.06559983, -0.06684648, -0.06480206, 
    -0.06653563, -0.0635647, -0.06900668, -0.06658766, -0.07103768, 
    -0.0705438, -0.06965935, -0.06767445, -0.0687388, -0.06749584, 
    -0.07027258, -0.07175955, -0.07214979, -0.07288342, -0.07213311, 
    -0.07219384, -0.07148276, -0.07171047, -0.07002712, -0.07092618, 
    -0.06840301, -0.06750561, -0.06503705, -0.0635703, -0.06211286, 
    -0.06148047, -0.06128934, -0.06120962,
  -0.08618436, -0.08427431, -0.08464228, -0.08312619, -0.08396385, 
    -0.08297601, -0.08579369, -0.08419929, -0.08521368, -0.08601075, 
    -0.08026178, -0.08305923, -0.07745771, -0.07916772, -0.07494314, 
    -0.07772122, -0.07439532, -0.07502203, -0.07315222, -0.07368302, 
    -0.07134265, -0.07290855, -0.07015957, -0.07171358, -0.07146812, 
    -0.07296077, -0.08248862, -0.08060474, -0.08260158, -0.08232987, 
    -0.08245172, -0.08394639, -0.08470985, -0.08633227, -0.08603545, 
    -0.08484502, -0.08220799, -0.08309384, -0.08087995, -0.08092929, 
    -0.07853318, -0.0796045, -0.07568466, -0.07677846, -0.07366079, 
    -0.07443253, -0.07369683, -0.07391915, -0.07369393, -0.07482911, 
    -0.07434057, -0.07534748, -0.0794027, -0.0781884, -0.08186672, 
    -0.08416208, -0.08572309, -0.08684841, -0.08668841, -0.0863842, 
    -0.08483811, -0.0834102, -0.08233833, -0.0816291, -0.08093638, 
    -0.07887513, -0.07780617, -0.07546532, -0.07588258, -0.0751772, 
    -0.07450975, -0.07340246, -0.07358358, -0.0730998, -0.07519584, 
    -0.07379606, -0.07612127, -0.07547799, -0.08074843, -0.08285394, 
    -0.08376505, -0.0845714, -0.08656559, -0.08518338, -0.08572555, 
    -0.08444153, -0.08363569, -0.0840333, -0.0816098, -0.08254344, 
    -0.07774328, -0.07977521, -0.07458729, -0.07579676, -0.07430034, 
    -0.07506018, -0.07376297, -0.07492942, -0.07292063, -0.07249044, 
    -0.07278412, -0.07166272, -0.07499461, -0.07369677, -0.08404443, 
    -0.08397944, -0.08367741, -0.08501331, -0.08509577, -0.08634039, 
    -0.08523209, -0.08476447, -0.08358926, -0.08290179, -0.08225363, 
    -0.08084653, -0.07930375, -0.07719647, -0.07571775, -0.07474263, 
    -0.07533909, -0.07481224, -0.07540141, -0.0756792, -0.07265128, 
    -0.074336, -0.07182293, -0.07195973, -0.07308831, -0.0719443, 
    -0.08393385, -0.08430831, -0.08562139, -0.08459204, -0.08647705, 
    -0.08541664, -0.08481284, -0.08252367, -0.08202932, -0.0815734, 
    -0.08068064, -0.07954931, -0.07760333, -0.07594954, -0.07447114, 
    -0.07457847, -0.07454067, -0.07421403, -0.0750257, -0.07408164, 
    -0.07392433, -0.07433628, -0.07197806, -0.07264394, -0.07196264, 
    -0.07239541, -0.08418642, -0.08355825, -0.08389708, -0.08326104, 
    -0.08370858, -0.08173687, -0.08115494, -0.07848736, -0.07957138, 
    -0.07785338, -0.07939518, -0.0791197, -0.0777977, -0.07931112, 
    -0.07603967, -0.07824208, -0.07420137, -0.0763465, -0.07406899, 
    -0.07447747, -0.07380244, -0.07320308, -0.07245617, -0.07109807, 
    -0.07141027, -0.07028947, -0.08263066, -0.08183198, -0.0819021, 
    -0.08107403, -0.08046705, -0.07916736, -0.07712696, -0.07788795, 
    -0.07649681, -0.07622054, -0.07833641, -0.07703023, -0.08130193, 
    -0.08059572, -0.08101553, -0.08256729, -0.07771175, -0.0801663, 
    -0.07569353, -0.07697891, -0.07328822, -0.07510056, -0.07158269, 
    -0.07012999, -0.06879062, -0.06725767, -0.08139953, -0.08193844, 
    -0.08097615, -0.0796634, -0.07846501, -0.07689986, -0.07674158, 
    -0.07645247, -0.07570887, -0.07508928, -0.07636117, -0.07493478, 
    -0.08043259, -0.07750238, -0.08214301, -0.08071657, -0.07974024, 
    -0.08016717, -0.07797544, -0.07746773, -0.07543882, -0.0764809, 
    -0.07048563, -0.07307696, -0.0661141, -0.06798916, -0.08212756, 
    -0.08140144, -0.07892445, -0.08009335, -0.07679657, -0.07600633, 
    -0.07537011, -0.07456449, -0.07447812, -0.07400549, -0.07478157, 
    -0.07403603, -0.07689656, -0.07560466, -0.07920381, -0.07831205, 
    -0.07872106, -0.07917211, -0.07778838, -0.07634095, -0.07631052, 
    -0.07585235, -0.07457589, -0.0767835, -0.07015771, -0.07417744, 
    -0.08061705, -0.0792499, -0.0790568, -0.07958224, -0.07608518, 
    -0.0773339, -0.074017, -0.07489899, -0.07345943, -0.07417122, 
    -0.07427651, -0.07520235, -0.07578461, -0.07727616, -0.07851173, 
    -0.07950584, -0.07927357, -0.07818548, -0.07625335, -0.07447021, 
    -0.07485714, -0.07356784, -0.07703091, -0.07555899, -0.07612441, 
    -0.07465903, -0.07790823, -0.07513196, -0.07863434, -0.07832079, 
    -0.0773589, -0.07546006, -0.07504667, -0.07460748, -0.07487822, 
    -0.07620497, -0.07642468, -0.07738218, -0.07764859, -0.07838897, 
    -0.07900725, -0.0784421, -0.07785297, -0.07620449, -0.07474913, 
    -0.07319456, -0.07281922, -0.07105312, -0.07248721, -0.07013591, 
    -0.07212954, -0.0687141, -0.07497447, -0.07218941, -0.07731548, 
    -0.07674599, -0.0757265, -0.07344021, -0.07466587, -0.07323458, 
    -0.07643332, -0.07814811, -0.07859835, -0.079445, -0.0785791, 
    -0.07864918, -0.0778288, -0.07809149, -0.07615037, -0.0771869, 
    -0.07427911, -0.07324582, -0.07040603, -0.06872053, -0.06704713, 
    -0.06632148, -0.06610221, -0.06601077,
  -0.06732005, -0.06577259, -0.06607072, -0.0648424, -0.06552106, 
    -0.06472072, -0.06700355, -0.06571181, -0.06653364, -0.06717939, 
    -0.06252159, -0.06478814, -0.06024957, -0.06163512, -0.05821211, 
    -0.06046309, -0.05776824, -0.05827603, -0.056761, -0.05719108, 
    -0.05529481, -0.05656356, -0.05433624, -0.05559535, -0.05539647, 
    -0.05660588, -0.06432582, -0.06279946, -0.06441735, -0.06419721, 
    -0.06429593, -0.06550692, -0.06612546, -0.06743988, -0.0671994, 
    -0.06623497, -0.06409846, -0.06481618, -0.06302244, -0.06306241, 
    -0.06112098, -0.06198902, -0.05881293, -0.0596992, -0.05717307, 
    -0.05779838, -0.05720227, -0.05738241, -0.05719993, -0.05811971, 
    -0.05772388, -0.05853973, -0.06182551, -0.06084162, -0.06382196, 
    -0.06568167, -0.06694635, -0.06785802, -0.0677284, -0.06748194, 
    -0.06622937, -0.06507249, -0.06420406, -0.06362943, -0.06306817, 
    -0.06139806, -0.06053193, -0.05863521, -0.0589733, -0.05840176, 
    -0.05786096, -0.05696376, -0.05711051, -0.05671853, -0.05841686, 
    -0.05728268, -0.0591667, -0.05864548, -0.06291588, -0.06462181, -0.06536, 
    -0.06601329, -0.0676289, -0.0665091, -0.06694835, -0.06590807, 
    -0.06525518, -0.06557732, -0.06361379, -0.06437024, -0.06048096, 
    -0.06212734, -0.05792378, -0.05890377, -0.05769127, -0.05830694, 
    -0.05725586, -0.05820099, -0.05657335, -0.05622479, -0.05646275, 
    -0.05555413, -0.05825381, -0.05720222, -0.06558634, -0.06553369, 
    -0.06528898, -0.06637131, -0.06643812, -0.06744646, -0.06654856, 
    -0.0661697, -0.06521757, -0.06466059, -0.06413543, -0.06299537, 
    -0.06174534, -0.0600379, -0.05883975, -0.05804964, -0.05853293, 
    -0.05810605, -0.05858343, -0.05880851, -0.05635512, -0.05772017, 
    -0.05568394, -0.05579478, -0.05670922, -0.05578228, -0.06549675, 
    -0.06580014, -0.06686395, -0.06603001, -0.06755716, -0.06669808, 
    -0.0662089, -0.06435423, -0.0639537, -0.0635843, -0.06286095, -0.0619443, 
    -0.06036756, -0.05902756, -0.05782966, -0.05791663, -0.057886, 
    -0.05762134, -0.058279, -0.05751407, -0.0573866, -0.05772039, 
    -0.05580964, -0.05634917, -0.05579714, -0.05614779, -0.06570138, 
    -0.06519245, -0.06546697, -0.06495164, -0.06531424, -0.06371675, 
    -0.06324524, -0.06108386, -0.06196219, -0.06057017, -0.06181942, 
    -0.06159622, -0.06052506, -0.06175131, -0.05910059, -0.06088512, 
    -0.05761108, -0.05934921, -0.05750381, -0.05783479, -0.05728785, 
    -0.05680221, -0.05619702, -0.05509663, -0.05534959, -0.05444149, 
    -0.06444091, -0.0637938, -0.06385062, -0.06317969, -0.0626879, 
    -0.06163483, -0.05998158, -0.06059818, -0.05947099, -0.05924714, 
    -0.06096155, -0.05990321, -0.06336434, -0.06279216, -0.0631323, 
    -0.06438956, -0.06045542, -0.06244422, -0.05882013, -0.05986162, 
    -0.05687119, -0.05833966, -0.05548929, -0.05431228, -0.05322711, 
    -0.05198516, -0.06344342, -0.06388006, -0.06310039, -0.06203675, 
    -0.06106574, -0.05979756, -0.05966932, -0.05943506, -0.05883255, 
    -0.05833052, -0.05936109, -0.05820533, -0.06265998, -0.06028577, 
    -0.06404581, -0.06289007, -0.062099, -0.06244492, -0.06066907, 
    -0.0602577, -0.05861374, -0.0594581, -0.05460043, -0.05670002, 
    -0.05105871, -0.05257778, -0.06403328, -0.06344496, -0.06143801, 
    -0.06238511, -0.05971387, -0.05907357, -0.05855807, -0.0579053, 
    -0.05783532, -0.05745237, -0.05808119, -0.05747712, -0.05979489, 
    -0.05874812, -0.06166436, -0.06094181, -0.06127321, -0.06163868, 
    -0.0605175, -0.05934471, -0.05932004, -0.05894881, -0.05791454, 
    -0.05970329, -0.05433474, -0.0575917, -0.06280943, -0.06170171, 
    -0.06154525, -0.06197098, -0.05913746, -0.06014926, -0.05746169, 
    -0.05817633, -0.05700992, -0.05758665, -0.05767197, -0.05842214, 
    -0.05889392, -0.06010247, -0.0611036, -0.06190908, -0.06172088, 
    -0.06083926, -0.05927372, -0.05782892, -0.05814243, -0.05709776, 
    -0.05990376, -0.05871111, -0.05916926, -0.05798191, -0.06061461, 
    -0.05836511, -0.06120295, -0.06094889, -0.06016951, -0.05863095, 
    -0.058296, -0.05794013, -0.0581595, -0.05923453, -0.05941255, 
    -0.06018838, -0.06040423, -0.06100413, -0.06150509, -0.06104719, 
    -0.06056984, -0.05923413, -0.05805491, -0.0567953, -0.05649118, 
    -0.05506022, -0.05622217, -0.05431708, -0.05593238, -0.05316512, 
    -0.0582375, -0.05598088, -0.06013433, -0.05967289, -0.05884684, 
    -0.05699435, -0.05798744, -0.05682774, -0.05941955, -0.06080898, 
    -0.06117379, -0.06185979, -0.06115819, -0.06121497, -0.06055026, 
    -0.0607631, -0.05919028, -0.06003015, -0.05767407, -0.05683684, 
    -0.05453593, -0.05317033, -0.05181458, -0.05122671, -0.05104908, 
    -0.05097499,
  -0.06391456, -0.06222175, -0.06254764, -0.06120573, -0.0619469, -0.0610729, 
    -0.06356808, -0.06215534, -0.06305389, -0.06376056, -0.05867596, 
    -0.0611465, -0.05620686, -0.05771168, -0.05399928, -0.05643857, 
    -0.05351921, -0.05406844, -0.05243101, -0.05289546, -0.05084996, 
    -0.05221789, -0.04981826, -0.05117374, -0.05095946, -0.05226356, 
    -0.06064199, -0.05897845, -0.06074184, -0.06050169, -0.06060938, 
    -0.06193145, -0.0626075, -0.06404578, -0.06378247, -0.06272724, 
    -0.06039399, -0.0611771, -0.05922126, -0.0592648, -0.05715295, 
    -0.05809651, -0.0546496, -0.0556099, -0.052876, -0.0535518, -0.05290755, 
    -0.05310217, -0.05290501, -0.05389932, -0.05347124, -0.05435381, 
    -0.05791869, -0.05684952, -0.06009248, -0.06212239, -0.06350548, 
    -0.06450379, -0.06436179, -0.06409185, -0.0627211, -0.06145694, 
    -0.06050916, -0.0598826, -0.05927106, -0.05745402, -0.05651328, 
    -0.05445718, -0.05482328, -0.05420449, -0.05361946, -0.05264993, 
    -0.05280843, -0.05238516, -0.05422083, -0.05299442, -0.05503277, 
    -0.0544683, -0.05910522, -0.06096495, -0.06177095, -0.06248485, 
    -0.06425279, -0.06302705, -0.06350766, -0.06236983, -0.06165646, 
    -0.06200837, -0.05986556, -0.06069045, -0.05645797, -0.05824696, 
    -0.0536874, -0.05474796, -0.053436, -0.05410188, -0.05296544, 
    -0.05398725, -0.05222845, -0.05185237, -0.0521091, -0.05112933, 
    -0.0540444, -0.0529075, -0.06201823, -0.0619607, -0.06169338, 
    -0.06287634, -0.0629494, -0.06405298, -0.06307022, -0.06265587, 
    -0.06161538, -0.06100727, -0.06043432, -0.05919177, -0.05783151, 
    -0.05597721, -0.05467864, -0.05382352, -0.05434645, -0.05388454, 
    -0.05440112, -0.05464481, -0.05199297, -0.05346724, -0.05126922, 
    -0.05138869, -0.05237511, -0.05137522, -0.06192034, -0.06225186, 
    -0.0634153, -0.06250314, -0.06417423, -0.06323379, -0.06269873, 
    -0.06067298, -0.06023612, -0.05983341, -0.0590454, -0.05804787, 
    -0.05633489, -0.05488204, -0.05358563, -0.05367967, -0.05364654, 
    -0.0533604, -0.05407165, -0.05324445, -0.0531067, -0.05346747, 
    -0.05140471, -0.05198655, -0.05139123, -0.05176932, -0.06214393, 
    -0.06158794, -0.0618878, -0.061325, -0.06172096, -0.05997778, 
    -0.05946396, -0.05711262, -0.05806733, -0.0565548, -0.05791207, 
    -0.0576694, -0.05650584, -0.057838, -0.05496115, -0.05689676, 
    -0.05334931, -0.05523052, -0.05323337, -0.05359117, -0.053, -0.0524755, 
    -0.05182242, -0.05063653, -0.05090896, -0.04993146, -0.06076755, 
    -0.06006179, -0.06012373, -0.05939254, -0.05885698, -0.05771137, 
    -0.05591612, -0.0565852, -0.05536251, -0.05511993, -0.05697977, 
    -0.05583112, -0.05959372, -0.05897049, -0.05934092, -0.06071154, 
    -0.05643024, -0.05859175, -0.05465739, -0.05578602, -0.05254998, 
    -0.05413729, -0.05105947, -0.04979249, -0.04862653, -0.04729471, 
    -0.05967988, -0.06015583, -0.05930616, -0.05814842, -0.05709295, 
    -0.05571656, -0.0555775, -0.05532357, -0.05467084, -0.0541274, 
    -0.0552434, -0.05399195, -0.05882659, -0.05624613, -0.06033657, 
    -0.0590771, -0.05821614, -0.05859251, -0.05666216, -0.05621567, 
    -0.05443393, -0.05534854, -0.05010244, -0.05236518, -0.04630309, 
    -0.04792986, -0.06032291, -0.05968157, -0.05749743, -0.05852742, 
    -0.05562581, -0.05493188, -0.05437366, -0.05366741, -0.05359174, 
    -0.05317777, -0.05385765, -0.05320452, -0.05571366, -0.05457941, 
    -0.05774348, -0.05695833, -0.05731835, -0.05771555, -0.05649763, 
    -0.05522564, -0.05519892, -0.05479674, -0.05367741, -0.05561433, 
    -0.04981665, -0.05332836, -0.0589893, -0.05778408, -0.05761399, 
    -0.05807689, -0.05500109, -0.05609801, -0.05318785, -0.05396057, 
    -0.05269978, -0.0533229, -0.05341513, -0.05422654, -0.0547373, 
    -0.05604725, -0.05713408, -0.05800956, -0.05780492, -0.05684696, 
    -0.05514873, -0.05358482, -0.05392389, -0.05279465, -0.05583171, 
    -0.05453935, -0.05503554, -0.05375027, -0.05660304, -0.05416483, 
    -0.057242, -0.05696603, -0.05611999, -0.05445257, -0.05409005, 
    -0.05370509, -0.05394236, -0.05510625, -0.05529917, -0.05614045, 
    -0.05637469, -0.05702602, -0.05757035, -0.05707279, -0.05655444, 
    -0.05510583, -0.05382922, -0.05246804, -0.05213978, -0.05059732, 
    -0.05184955, -0.04979766, -0.05153703, -0.04855999, -0.05402675, 
    -0.05158933, -0.05608182, -0.05558137, -0.05468632, -0.05268296, 
    -0.05375625, -0.05250306, -0.05530675, -0.05681408, -0.05721032, 
    -0.05795596, -0.05719337, -0.05725506, -0.05653318, -0.05676426, 
    -0.05505832, -0.0559688, -0.05341741, -0.05251289, -0.05003305, 
    -0.04856558, -0.04711202, -0.04648279, -0.0462928, -0.04621357,
  -0.04035198, -0.0390736, -0.03931955, -0.03830725, -0.03886621, 
    -0.03820712, -0.04009017, -0.03902348, -0.03970178, -0.04023561, 
    -0.03640242, -0.0382626, -0.03454812, -0.03567765, -0.03289467, 
    -0.03472192, -0.03253571, -0.03294641, -0.03172284, -0.03206963, 
    -0.03054396, -0.03156378, -0.02977613, -0.03078517, -0.03062552, 
    -0.03159786, -0.03788237, -0.03662993, -0.0379576, -0.03777666, 
    -0.03785779, -0.03885456, -0.03936474, -0.04045115, -0.04025216, 
    -0.03945513, -0.03769552, -0.03828567, -0.03681261, -0.03684536, 
    -0.03525804, -0.03596681, -0.03338129, -0.03410058, -0.0320551, 
    -0.03256007, -0.03207866, -0.03222405, -0.03207677, -0.03281992, 
    -0.03249985, -0.03315992, -0.03583318, -0.03503028, -0.03746842, 
    -0.03899862, -0.04004287, -0.0407974, -0.04069004, -0.04048598, 
    -0.0394505, -0.03849667, -0.03778229, -0.03731038, -0.03685008, 
    -0.03548411, -0.03477797, -0.03323727, -0.03351132, -0.03304819, 
    -0.03261065, -0.03188627, -0.03200463, -0.03168861, -0.03306042, 
    -0.03214355, -0.0336682, -0.03324559, -0.0367253, -0.03812575, 
    -0.03873349, -0.03927216, -0.04060763, -0.03968151, -0.04004452, 
    -0.03918535, -0.03864713, -0.03891259, -0.03729755, -0.03791888, 
    -0.03473647, -0.03607989, -0.03266145, -0.03345493, -0.03247351, 
    -0.03297143, -0.0321219, -0.03288567, -0.03157166, -0.03129109, 
    -0.0314826, -0.03075208, -0.03292842, -0.03207862, -0.03892003, 
    -0.03887663, -0.03867498, -0.03956771, -0.03962288, -0.0404566, 
    -0.03971411, -0.03940125, -0.03861615, -0.03815765, -0.0377259, 
    -0.03679042, -0.03576768, -0.03437592, -0.03340304, -0.03276323, 
    -0.03315441, -0.03280886, -0.03319532, -0.03337771, -0.03139596, 
    -0.03249686, -0.03085632, -0.03094536, -0.03168111, -0.03093532, 
    -0.03884618, -0.03909632, -0.03997475, -0.03928596, -0.04054825, 
    -0.03983765, -0.03943361, -0.03790571, -0.0375766, -0.03727335, 
    -0.0366803, -0.03593025, -0.03464415, -0.03355532, -0.03258536, 
    -0.03265567, -0.0326309, -0.03241701, -0.03294881, -0.03233036, 
    -0.03222743, -0.03249704, -0.0309573, -0.03139117, -0.03094725, 
    -0.03122915, -0.03901488, -0.03859545, -0.03882163, -0.03839717, 
    -0.03869578, -0.03738205, -0.03699524, -0.03522776, -0.03594487, 
    -0.03480912, -0.0358282, -0.03564588, -0.03477238, -0.03577255, 
    -0.03361456, -0.03506573, -0.03240872, -0.03381632, -0.03232208, 
    -0.0325895, -0.03214772, -0.03175605, -0.03126875, -0.03038502, 
    -0.0305879, -0.02986032, -0.03797698, -0.03744531, -0.03749195, 
    -0.03694149, -0.03653856, -0.03567742, -0.03433011, -0.03483193, 
    -0.0339152, -0.03373348, -0.03512803, -0.03426639, -0.03709291, 
    -0.03662394, -0.03690264, -0.03793477, -0.03471567, -0.0363391, 
    -0.03338712, -0.03423258, -0.03181165, -0.03299792, -0.03070002, 
    -0.02975697, -0.0288907, -0.02790317, -0.03715777, -0.03751613, 
    -0.03687649, -0.03600582, -0.035213, -0.03418051, -0.0340763, 
    -0.03388602, -0.0333972, -0.03299051, -0.03382597, -0.03288919, 
    -0.03651571, -0.03457757, -0.03765227, -0.03670414, -0.03605672, 
    -0.03633967, -0.03488967, -0.03455473, -0.03321987, -0.03390473, 
    -0.02998751, -0.0316737, -0.02716935, -0.02837386, -0.03764197, 
    -0.03715903, -0.03551672, -0.03629073, -0.0341125, -0.03359265, 
    -0.03317477, -0.0326465, -0.03258993, -0.03228053, -0.03278875, 
    -0.03230052, -0.03417834, -0.03332876, -0.03570154, -0.03511194, 
    -0.03538223, -0.03568056, -0.03476623, -0.03381266, -0.03379264, 
    -0.03349146, -0.03265398, -0.0341039, -0.02977493, -0.03239306, 
    -0.03663809, -0.03573205, -0.03560426, -0.03595206, -0.03364448, 
    -0.03446649, -0.03228806, -0.03286573, -0.0319235, -0.03238898, 
    -0.03245791, -0.03306469, -0.03344695, -0.03442843, -0.03524387, 
    -0.03590146, -0.0357477, -0.03502835, -0.03375505, -0.03258475, 
    -0.03283829, -0.03199435, -0.03426683, -0.03329877, -0.03367027, 
    -0.03270845, -0.03484531, -0.03301852, -0.0353249, -0.03511772, 
    -0.03448297, -0.03323382, -0.03296257, -0.03267467, -0.03285211, 
    -0.03372324, -0.03386774, -0.03449832, -0.034674, -0.03516275, 
    -0.03557148, -0.03519786, -0.03480885, -0.03372291, -0.03276749, 
    -0.03175048, -0.0315055, -0.03035583, -0.03128899, -0.02976081, 
    -0.03105594, -0.02884131, -0.03291522, -0.03109493, -0.03445435, 
    -0.0340792, -0.03340878, -0.03191094, -0.03271293, -0.03177662, 
    -0.03387342, -0.03500368, -0.03530111, -0.03586118, -0.03528839, 
    -0.03533471, -0.0347929, -0.03496629, -0.03368733, -0.03436961, 
    -0.03245961, -0.03178396, -0.02993589, -0.02884545, -0.02776788, 
    -0.02730224, -0.02716173, -0.02710316,
  -0.01970498, -0.01870054, -0.01889315, -0.01810236, -0.01853836, 
    -0.01802443, -0.01949861, -0.01866132, -0.0191931, -0.01961321, 
    -0.01662923, -0.0180676, -0.01521544, -0.01607415, -0.01397336, 
    -0.01534705, -0.01370618, -0.01401194, -0.01310463, -0.01336067, 
    -0.01224115, -0.0129875, -0.01168477, -0.01241693, -0.01230054, 
    -0.01301258, -0.01777204, -0.01680411, -0.01783047, -0.01769001, 
    -0.01775297, -0.01852925, -0.01892857, -0.01978323, -0.01962626, 
    -0.01899946, -0.01762709, -0.01808556, -0.01694474, -0.01696998, 
    -0.01575423, -0.01629523, -0.01433699, -0.01487744, -0.01334993, 
    -0.01372429, -0.01336735, -0.01347497, -0.01336595, -0.01391764, 
    -0.01367955, -0.01417136, -0.016193, -0.01558102, -0.01745117, 
    -0.01864188, -0.01946137, -0.02005681, -0.01997192, -0.01981072, 
    -0.01899583, -0.01824993, -0.01769438, -0.01732891, -0.01697361, 
    -0.01592645, -0.01538954, -0.0142292, -0.01443443, -0.0140879, 
    -0.01376189, -0.01322518, -0.01331261, -0.01307941, -0.01409703, 
    -0.01341536, -0.01455215, -0.01423542, -0.01687751, -0.01796114, 
    -0.01843468, -0.01885602, -0.0199068, -0.01917717, -0.01946267, 
    -0.01878802, -0.01836728, -0.01857461, -0.01731899, -0.01780039, 
    -0.01535808, -0.01638183, -0.01379967, -0.01439216, -0.01365998, 
    -0.0140306, -0.01339934, -0.01396665, -0.0129933, -0.01278713, 
    -0.01292779, -0.01239279, -0.01399853, -0.01336732, -0.01858043, 
    -0.0185465, -0.01838901, -0.0190878, -0.01913112, -0.01978753, 
    -0.01920278, -0.01895721, -0.01834311, -0.01798595, -0.01765065, 
    -0.01692765, -0.01614293, -0.01508524, -0.01435328, -0.01387542, 
    -0.01416725, -0.0139094, -0.01419783, -0.01433431, -0.01286412, 
    -0.01367732, -0.01246887, -0.01253393, -0.01307388, -0.01252659, 
    -0.01852271, -0.01871832, -0.01940775, -0.01886683, -0.01985989, 
    -0.01929989, -0.01898258, -0.01779017, -0.01753494, -0.01730028, 
    -0.01684286, -0.01626726, -0.01528814, -0.01446743, -0.01374308, 
    -0.01379537, -0.01377694, -0.01361804, -0.01401373, -0.01355376, 
    -0.01347748, -0.01367746, -0.01254266, -0.0128606, -0.01253532, 
    -0.0127417, -0.01865459, -0.01832696, -0.01850353, -0.01817239, 
    -0.01840525, -0.01738434, -0.01708553, -0.01573118, -0.01627845, 
    -0.01541315, -0.0161892, -0.01604989, -0.0153853, -0.01614666, 
    -0.01451188, -0.01560796, -0.01361189, -0.01466344, -0.01354762, 
    -0.01374616, -0.01341845, -0.01312911, -0.01277075, -0.01212558, 
    -0.01227314, -0.01174553, -0.01784551, -0.01743328, -0.01746939, 
    -0.01704408, -0.01673384, -0.01607397, -0.01505064, -0.01543046, 
    -0.01473782, -0.01460118, -0.01565532, -0.01500252, -0.0171609, 
    -0.01679951, -0.01701413, -0.01781273, -0.01534232, -0.01658061, 
    -0.01434136, -0.014977, -0.01317011, -0.01405037, -0.01235483, 
    -0.01167095, -0.01104943, -0.01034922, -0.01721098, -0.0174881, 
    -0.01699397, -0.0163251, -0.01571995, -0.01493772, -0.01485914, 
    -0.01471587, -0.0143489, -0.01404485, -0.0146707, -0.01396927, 
    -0.01671627, -0.01523773, -0.01759356, -0.01686122, -0.01636408, 
    -0.01658105, -0.01547426, -0.01522044, -0.01421619, -0.01472995, 
    -0.01183745, -0.01306842, -0.009834968, -0.01068182, -0.01758559, 
    -0.01721196, -0.01595132, -0.01654349, -0.01488643, -0.01449544, 
    -0.01418246, -0.01378855, -0.01374648, -0.01351682, -0.01389443, 
    -0.01353163, -0.01493608, -0.01429766, -0.0160924, -0.01564309, 
    -0.0158488, -0.01607637, -0.01538063, -0.0146607, -0.01464565, 
    -0.01441954, -0.01379411, -0.01487995, -0.0116839, -0.01360027, 
    -0.01681039, -0.0161157, -0.01601812, -0.01628395, -0.01453434, 
    -0.0151537, -0.0135224, -0.01395178, -0.01325267, -0.01359724, 
    -0.0136484, -0.01410022, -0.01438618, -0.01512493, -0.01574344, 
    -0.01624523, -0.01612766, -0.01557956, -0.01461739, -0.01374263, 
    -0.01393133, -0.01330501, -0.01500286, -0.01427521, -0.01455371, 
    -0.01383464, -0.01544061, -0.01406575, -0.01580513, -0.01564748, 
    -0.01516616, -0.01422662, -0.014024, -0.0138095, -0.01394163, 
    -0.01459349, -0.01470212, -0.01517777, -0.01531075, -0.01568172, 
    -0.0159931, -0.01570843, -0.01541295, -0.01459324, -0.01387859, 
    -0.01312501, -0.01294462, -0.01210438, -0.01278559, -0.01167372, 
    -0.01261482, -0.01101419, -0.01398868, -0.01264336, -0.01514452, 
    -0.01486133, -0.01435758, -0.0132434, -0.01383797, -0.01314428, 
    -0.01470639, -0.01556082, -0.01578701, -0.01621442, -0.01577733, 
    -0.0158126, -0.01540086, -0.01553242, -0.01456652, -0.01508047, 
    -0.01364966, -0.01314969, -0.01180012, -0.01101715, -0.01025401, 
    -0.009927696, -0.009829662, -0.009788851,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15 ;

 SOILWATER_10CM =
  297.7622, 299.0222, 298.777, 299.7947, 299.2303, 299.8961, 298.0175, 
    299.0722, 298.3986, 297.8757, 301.7654, 299.8399, 303.777, 302.5413, 
    305.6483, 303.5843, 306.0594, 305.5899, 307.0056, 306.5996, 308.4153, 
    307.1932, 309.3603, 308.1233, 308.3164, 307.1529, 300.2269, 301.525, 
    300.1501, 300.3349, 300.252, 299.2419, 298.7317, 297.6663, 297.8595, 
    298.6422, 300.4181, 299.8169, 301.3345, 301.3001, 302.9964, 302.2307, 
    305.093, 304.2775, 306.6165, 306.0319, 306.589, 306.42, 306.5912, 
    305.7341, 306.101, 305.347, 302.3739, 303.2453, 300.6519, 299.0967, 
    298.0636, 297.332, 297.4353, 297.6324, 298.6468, 299.6033, 300.3295, 
    300.8156, 301.2952, 302.7498, 303.5226, 305.258, 304.9445, 305.4737, 
    305.9738, 306.8137, 306.6753, 307.0457, 305.4601, 306.5132, 304.766, 
    305.2488, 301.4246, 299.979, 299.3633, 298.8241, 297.5148, 298.4184, 
    298.0619, 298.9108, 299.451, 299.1838, 300.8289, 300.1897, 303.5685, 
    302.1095, 305.9154, 305.0089, 306.1315, 305.5616, 306.5385, 305.6592, 
    307.1838, 307.5164, 307.2891, 308.1635, 305.6105, 306.5889, 299.1763, 
    299.2198, 299.423, 298.5308, 298.4763, 297.6609, 298.3865, 298.6958, 
    299.4825, 299.9466, 300.3871, 301.3576, 302.4441, 303.9689, 305.0682, 
    305.799, 305.3533, 305.7469, 305.3067, 305.0974, 307.3917, 306.1044, 
    308.0377, 307.9305, 307.0545, 307.9425, 299.2505, 298.9998, 298.1303, 
    298.8106, 297.5723, 298.2648, 298.6635, 300.2028, 300.5406, 300.8538, 
    301.4734, 302.2698, 303.6709, 304.8942, 306.0029, 305.9222, 305.9506, 
    306.1966, 305.5873, 306.2968, 306.4159, 306.1044, 307.9161, 307.3977, 
    307.9282, 307.5906, 299.0813, 299.5033, 299.2752, 299.704, 299.4019, 
    300.7409, 301.1428, 303.029, 302.2541, 303.4885, 302.3794, 302.5756, 
    303.5283, 302.4393, 304.8264, 303.206, 306.2062, 304.5971, 306.3064, 
    305.9981, 306.5087, 306.9665, 307.5433, 308.6095, 308.3624, 309.2559, 
    300.1305, 300.6758, 300.6279, 301.1995, 301.6227, 302.5417, 304.0202, 
    303.4637, 304.4862, 304.6918, 303.1386, 304.0913, 301.0413, 301.5322, 
    301.24, 300.1733, 303.5916, 301.8334, 305.0864, 304.1293, 306.9011, 
    305.5309, 308.2264, 309.3837, 310.477, 311.7573, 300.9739, 300.603, 
    301.2675, 302.1885, 303.0456, 304.1876, 304.3047, 304.5191, 305.075, 
    305.5398, 304.5867, 305.6552, 301.6457, 303.7446, 300.4627, 301.4477, 
    302.1342, 301.8332, 303.4001, 303.7703, 305.2781, 304.4981, 309.0976, 
    307.0629, 312.7355, 311.142, 300.4734, 300.9727, 302.7151, 301.8852, 
    304.2641, 304.8518, 305.3302, 305.9324, 305.9976, 306.3544, 305.7698, 
    306.3314, 304.19, 305.1533, 302.5158, 303.156, 302.8615, 302.5385, 
    303.5362, 304.6017, 304.6248, 304.967, 305.9222, 304.2737, 309.3603, 
    306.2228, 301.5179, 302.4823, 302.6207, 302.2466, 304.7928, 303.8683, 
    306.3457, 305.682, 306.7702, 306.229, 306.1494, 305.4553, 305.018, 
    303.9105, 303.0118, 302.3008, 302.4661, 303.2475, 304.667, 306.0033, 
    305.7129, 306.6874, 304.0911, 305.1875, 304.7633, 305.8616, 303.4488, 
    305.5063, 302.9238, 303.1499, 303.8499, 305.2618, 305.5717, 305.9001, 
    305.6975, 304.7032, 304.5397, 303.833, 303.6379, 303.1006, 302.6563, 
    303.0622, 303.4889, 304.7037, 305.7939, 306.9729, 307.2621, 308.6444, 
    307.5183, 309.3778, 307.7956, 310.5388, 305.6246, 307.7499, 303.8819, 
    304.3015, 305.0612, 306.7842, 305.8565, 306.9419, 304.5333, 303.2743, 
    302.9497, 302.344, 302.9635, 302.9131, 303.5068, 303.3159, 304.7441, 
    303.9763, 306.1474, 306.9334, 309.1621, 310.5343, 311.9366, 312.557, 
    312.746, 312.8251 ;

 SOMC_FIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOMHR =
  6.358298e-08, 6.386256e-08, 6.380821e-08, 6.403371e-08, 6.390862e-08, 
    6.405628e-08, 6.363966e-08, 6.387366e-08, 6.372428e-08, 6.360815e-08, 
    6.447134e-08, 6.404377e-08, 6.491543e-08, 6.464276e-08, 6.532771e-08, 
    6.4873e-08, 6.541939e-08, 6.531458e-08, 6.563002e-08, 6.553965e-08, 
    6.594313e-08, 6.567172e-08, 6.615226e-08, 6.58783e-08, 6.592116e-08, 
    6.566277e-08, 6.412981e-08, 6.441811e-08, 6.411273e-08, 6.415384e-08, 
    6.413539e-08, 6.39112e-08, 6.379823e-08, 6.356161e-08, 6.360457e-08, 
    6.377836e-08, 6.417233e-08, 6.403859e-08, 6.437563e-08, 6.436802e-08, 
    6.474324e-08, 6.457406e-08, 6.520471e-08, 6.502547e-08, 6.554342e-08, 
    6.541316e-08, 6.553731e-08, 6.549966e-08, 6.55378e-08, 6.534675e-08, 
    6.542861e-08, 6.52605e-08, 6.460575e-08, 6.479818e-08, 6.422425e-08, 
    6.387916e-08, 6.364992e-08, 6.348726e-08, 6.351026e-08, 6.35541e-08, 
    6.377937e-08, 6.399117e-08, 6.415257e-08, 6.426054e-08, 6.436692e-08, 
    6.468895e-08, 6.485936e-08, 6.524096e-08, 6.517209e-08, 6.528876e-08, 
    6.540021e-08, 6.558732e-08, 6.555653e-08, 6.563896e-08, 6.528568e-08, 
    6.552047e-08, 6.513286e-08, 6.523888e-08, 6.439587e-08, 6.407466e-08, 
    6.393816e-08, 6.381866e-08, 6.352794e-08, 6.372871e-08, 6.364956e-08, 
    6.383784e-08, 6.395748e-08, 6.389831e-08, 6.42635e-08, 6.412152e-08, 
    6.486947e-08, 6.454731e-08, 6.53872e-08, 6.518622e-08, 6.543538e-08, 
    6.530824e-08, 6.552609e-08, 6.533003e-08, 6.566965e-08, 6.57436e-08, 
    6.569307e-08, 6.588719e-08, 6.531916e-08, 6.553731e-08, 6.389665e-08, 
    6.39063e-08, 6.395126e-08, 6.375364e-08, 6.374155e-08, 6.356043e-08, 
    6.372159e-08, 6.379021e-08, 6.396441e-08, 6.406746e-08, 6.416541e-08, 
    6.438078e-08, 6.462131e-08, 6.495763e-08, 6.519925e-08, 6.536121e-08, 
    6.52619e-08, 6.534958e-08, 6.525156e-08, 6.520562e-08, 6.571589e-08, 
    6.542937e-08, 6.585927e-08, 6.583548e-08, 6.564093e-08, 6.583816e-08, 
    6.391308e-08, 6.385754e-08, 6.366474e-08, 6.381563e-08, 6.35407e-08, 
    6.369459e-08, 6.378308e-08, 6.412449e-08, 6.41995e-08, 6.426905e-08, 
    6.440642e-08, 6.458272e-08, 6.489199e-08, 6.516106e-08, 6.540669e-08, 
    6.538869e-08, 6.539503e-08, 6.54499e-08, 6.531398e-08, 6.547221e-08, 
    6.549877e-08, 6.542933e-08, 6.58323e-08, 6.571717e-08, 6.583497e-08, 
    6.576001e-08, 6.38756e-08, 6.396904e-08, 6.391854e-08, 6.40135e-08, 
    6.394661e-08, 6.424406e-08, 6.433323e-08, 6.475051e-08, 6.457925e-08, 
    6.48518e-08, 6.460694e-08, 6.465033e-08, 6.486071e-08, 6.462017e-08, 
    6.514622e-08, 6.478959e-08, 6.545203e-08, 6.50959e-08, 6.547435e-08, 
    6.540562e-08, 6.551941e-08, 6.562132e-08, 6.574952e-08, 6.598609e-08, 
    6.59313e-08, 6.612913e-08, 6.410834e-08, 6.422955e-08, 6.421887e-08, 
    6.434571e-08, 6.443951e-08, 6.464282e-08, 6.496889e-08, 6.484628e-08, 
    6.507138e-08, 6.511657e-08, 6.477458e-08, 6.498456e-08, 6.431066e-08, 
    6.441955e-08, 6.435471e-08, 6.411791e-08, 6.487454e-08, 6.448624e-08, 
    6.520325e-08, 6.49929e-08, 6.560679e-08, 6.53015e-08, 6.590115e-08, 
    6.615751e-08, 6.639875e-08, 6.668071e-08, 6.429569e-08, 6.421333e-08, 
    6.436079e-08, 6.456481e-08, 6.475408e-08, 6.500573e-08, 6.503147e-08, 
    6.507862e-08, 6.520072e-08, 6.53034e-08, 6.509353e-08, 6.532913e-08, 
    6.444481e-08, 6.490824e-08, 6.41822e-08, 6.440084e-08, 6.455278e-08, 
    6.448612e-08, 6.483226e-08, 6.491384e-08, 6.524535e-08, 6.507398e-08, 
    6.609424e-08, 6.564286e-08, 6.689538e-08, 6.654536e-08, 6.418456e-08, 
    6.429541e-08, 6.468117e-08, 6.449763e-08, 6.502253e-08, 6.515172e-08, 
    6.525676e-08, 6.539102e-08, 6.540552e-08, 6.548507e-08, 6.53547e-08, 
    6.547992e-08, 6.500627e-08, 6.521793e-08, 6.463707e-08, 6.477845e-08, 
    6.471341e-08, 6.464207e-08, 6.486225e-08, 6.509683e-08, 6.510184e-08, 
    6.517705e-08, 6.538904e-08, 6.502465e-08, 6.615252e-08, 6.545599e-08, 
    6.441627e-08, 6.462978e-08, 6.466026e-08, 6.457756e-08, 6.513877e-08, 
    6.493543e-08, 6.548313e-08, 6.53351e-08, 6.557763e-08, 6.545712e-08, 
    6.543939e-08, 6.52846e-08, 6.518822e-08, 6.494476e-08, 6.474665e-08, 
    6.458955e-08, 6.462608e-08, 6.479865e-08, 6.511118e-08, 6.540683e-08, 
    6.534207e-08, 6.55592e-08, 6.498447e-08, 6.522547e-08, 6.513232e-08, 
    6.537519e-08, 6.484301e-08, 6.529623e-08, 6.472717e-08, 6.477707e-08, 
    6.493139e-08, 6.524182e-08, 6.531049e-08, 6.538382e-08, 6.533857e-08, 
    6.511911e-08, 6.508316e-08, 6.492764e-08, 6.488471e-08, 6.47662e-08, 
    6.46681e-08, 6.475774e-08, 6.485187e-08, 6.51192e-08, 6.536012e-08, 
    6.562277e-08, 6.568705e-08, 6.599396e-08, 6.574413e-08, 6.61564e-08, 
    6.580591e-08, 6.641262e-08, 6.532247e-08, 6.579559e-08, 6.493841e-08, 
    6.503075e-08, 6.519779e-08, 6.558088e-08, 6.537405e-08, 6.561592e-08, 
    6.508175e-08, 6.480461e-08, 6.473289e-08, 6.459911e-08, 6.473595e-08, 
    6.472482e-08, 6.485576e-08, 6.481368e-08, 6.512808e-08, 6.49592e-08, 
    6.543894e-08, 6.561401e-08, 6.610841e-08, 6.641149e-08, 6.671998e-08, 
    6.685619e-08, 6.689764e-08, 6.691497e-08 ;

 SOM_C_LEACHED =
  -2.223797e-20, -5.202761e-20, -6.1968e-21, -4.252685e-21, 1.225423e-20, 
    2.675787e-20, -2.124882e-20, -2.153454e-20, 5.112679e-20, 5.38149e-20, 
    -7.521117e-20, 3.421186e-20, -2.459155e-20, 1.447693e-20, 6.011282e-20, 
    3.372518e-21, -7.137694e-20, 4.708659e-20, -2.273515e-20, -1.666837e-20, 
    -5.638862e-20, 1.421885e-20, -6.742819e-20, -7.228885e-20, 7.827053e-20, 
    1.126088e-20, -4.267727e-20, 6.610116e-20, -1.063266e-20, -3.057475e-20, 
    3.413492e-20, -1.644827e-20, 1.076703e-20, 2.081516e-20, 8.05783e-20, 
    -2.728366e-20, 1.427799e-20, -6.257526e-20, 8.741224e-21, 2.188234e-20, 
    2.389386e-20, -1.526928e-20, 2.176049e-20, 4.550534e-20, -1.571619e-20, 
    2.937337e-20, -5.659279e-20, 9.753454e-21, -1.104938e-20, 3.400927e-20, 
    1.686119e-20, -1.762136e-21, -3.821576e-20, -9.77524e-20, -4.832142e-20, 
    2.039208e-21, -5.739467e-20, -9.791103e-21, 2.672248e-20, -4.64421e-21, 
    -3.109905e-21, -4.195872e-20, 2.213919e-21, -1.093254e-20, 3.690402e-20, 
    -4.402832e-20, -2.306055e-20, 1.228793e-20, 4.071221e-20, 6.482651e-20, 
    2.153361e-20, 4.604599e-21, 1.282182e-20, -2.648278e-20, 6.958326e-21, 
    -6.577641e-20, 1.540388e-20, 3.5756e-21, -4.947176e-20, 6.818034e-20, 
    3.20635e-20, -3.309649e-20, 4.880414e-20, 3.784079e-20, 1.412069e-20, 
    1.558751e-20, -2.533604e-20, -3.716054e-20, -1.22903e-21, -8.631225e-20, 
    3.332803e-20, 1.043664e-20, 3.306648e-20, -1.816995e-20, 3.427514e-20, 
    -5.868562e-21, -1.130259e-20, 2.870768e-21, 1.106104e-20, -7.193995e-21, 
    -3.9398e-20, 1.885334e-20, -4.648365e-20, -1.141754e-20, -1.198276e-20, 
    -3.202359e-20, 5.094408e-20, 8.061835e-20, -3.341136e-20, 1.939364e-20, 
    -1.854e-20, 8.559573e-21, -2.995358e-20, -3.460148e-20, -3.87773e-20, 
    2.11958e-20, -2.993575e-20, 9.214168e-20, 8.443755e-21, 3.676055e-20, 
    5.123637e-21, 8.777982e-21, 5.80989e-20, -4.003784e-20, -2.271953e-20, 
    4.634401e-20, 6.085826e-21, 5.066711e-20, -1.079063e-20, 6.75566e-20, 
    1.490086e-20, 3.887903e-20, 1.355153e-20, -3.226133e-20, -2.12791e-20, 
    -5.537252e-20, 6.461627e-20, -4.958244e-20, 3.031862e-20, -4.766319e-20, 
    1.077816e-20, 3.66924e-20, 6.837876e-21, 4.786225e-21, -1.332016e-20, 
    7.671508e-20, 1.354065e-20, -3.229185e-20, 4.824912e-20, 4.345599e-20, 
    3.434971e-20, 1.892053e-20, 1.27041e-20, -5.760588e-20, -1.325098e-20, 
    3.449634e-20, 1.076742e-20, -6.54829e-21, -3.273555e-21, 5.171955e-20, 
    -3.80579e-20, 4.001184e-21, -4.159458e-20, 1.743163e-20, 2.348224e-20, 
    3.792314e-20, -7.207389e-20, 4.408261e-22, -1.587462e-20, -7.919484e-21, 
    -2.06827e-21, -3.310806e-21, -1.583431e-21, 1.929723e-20, -2.737654e-21, 
    -1.452459e-20, -9.401354e-21, -7.935338e-20, 4.23973e-20, 3.071554e-20, 
    3.952595e-20, 2.097118e-20, -2.435287e-20, -2.426268e-21, -2.14688e-20, 
    -3.166871e-20, -7.626869e-21, 5.688116e-20, -1.770157e-20, 6.75487e-20, 
    -6.501684e-20, -3.647561e-20, -5.243606e-20, -5.4787e-20, 8.701713e-20, 
    1.60387e-20, -5.002666e-20, 1.881594e-20, -1.005869e-20, -1.253205e-20, 
    -6.73924e-20, -5.205705e-20, 3.278813e-20, 4.391977e-20, 3.032959e-20, 
    1.973726e-20, 6.834211e-20, 5.651418e-20, 2.27319e-21, 1.659029e-20, 
    6.110557e-20, -1.24881e-21, -8.00206e-21, -1.854993e-20, -2.52828e-20, 
    3.24319e-20, -5.161256e-20, 5.337239e-20, 4.177545e-20, 2.29369e-20, 
    3.830731e-20, 1.82251e-20, -4.911847e-21, 3.968935e-21, -4.221221e-21, 
    -6.921879e-20, 5.166927e-20, 8.154457e-22, -1.717649e-20, -2.663136e-21, 
    2.603328e-20, -1.502519e-20, -3.946289e-20, 8.468988e-20, 1.601859e-21, 
    3.505915e-20, 2.75448e-20, 1.084218e-22, -3.793549e-20, -3.572481e-20, 
    -9.602171e-22, -5.101267e-20, 2.309779e-20, -5.098517e-20, 2.272713e-20, 
    -4.852941e-20, 2.668059e-20, 2.212031e-20, 5.005751e-20, -2.454467e-21, 
    -2.786692e-20, -1.342589e-20, -2.368768e-20, -3.534884e-20, 
    -5.589144e-21, 4.723392e-20, -4.755218e-20, 3.298229e-20, -3.844398e-20, 
    1.636814e-20, -3.945383e-20, -3.377157e-20, 1.671995e-20, -4.181757e-20, 
    7.316284e-20, 1.124621e-20, -5.555521e-20, 4.008826e-20, -1.948983e-20, 
    -6.103573e-21, -2.041127e-21, 5.594649e-20, -8.746828e-21, 1.19673e-20, 
    2.013692e-20, -5.883433e-20, -3.0347e-20, -3.497904e-20, -2.229049e-20, 
    -2.002508e-20, 6.358039e-21, 2.252112e-20, -7.398351e-20, 6.178532e-21, 
    -3.823069e-20, 1.465145e-20, 3.376874e-20, -2.457565e-20, 3.302312e-20, 
    3.925869e-20, -5.272225e-20, 1.443428e-20, 3.001516e-20, 4.502797e-20, 
    -1.197266e-20, 7.473942e-20, -1.473354e-20, 1.841806e-20, -8.592446e-22, 
    -2.89722e-20, -3.219509e-20, -2.320575e-20, 4.188482e-21, 6.736523e-21, 
    -2.230177e-20, 9.776845e-20, -4.835648e-20, 2.395332e-20, 7.176027e-22, 
    2.325508e-20, 2.349993e-20, -2.25638e-20, 3.041519e-21, -2.253057e-20, 
    -2.618901e-22, 2.451379e-20, -3.986113e-20, 3.733807e-21, 3.430637e-20, 
    3.906661e-20, 2.069844e-20, 4.498759e-22, 4.893834e-21, -1.566504e-20, 
    5.655004e-20, -5.676762e-21, 4.867069e-21, -5.429501e-20, 4.356163e-20, 
    7.219913e-22, 2.435606e-20, -6.065307e-20, -3.183123e-20, -2.545161e-20, 
    1.936009e-20, 6.699051e-20, -2.037428e-20, -7.384228e-21 ;

 SR =
  6.358388e-08, 6.386347e-08, 6.380911e-08, 6.403462e-08, 6.390952e-08, 
    6.405718e-08, 6.364056e-08, 6.387457e-08, 6.372518e-08, 6.360905e-08, 
    6.447225e-08, 6.404468e-08, 6.491634e-08, 6.464366e-08, 6.532863e-08, 
    6.487392e-08, 6.542031e-08, 6.53155e-08, 6.563094e-08, 6.554057e-08, 
    6.594404e-08, 6.567264e-08, 6.615318e-08, 6.587923e-08, 6.592209e-08, 
    6.566369e-08, 6.413072e-08, 6.441902e-08, 6.411364e-08, 6.415475e-08, 
    6.41363e-08, 6.391211e-08, 6.379913e-08, 6.356251e-08, 6.360547e-08, 
    6.377926e-08, 6.417324e-08, 6.403949e-08, 6.437654e-08, 6.436893e-08, 
    6.474416e-08, 6.457498e-08, 6.520563e-08, 6.502638e-08, 6.554434e-08, 
    6.541408e-08, 6.553822e-08, 6.550058e-08, 6.553871e-08, 6.534768e-08, 
    6.542952e-08, 6.526142e-08, 6.460666e-08, 6.47991e-08, 6.422516e-08, 
    6.388007e-08, 6.365083e-08, 6.348817e-08, 6.351116e-08, 6.3555e-08, 
    6.378028e-08, 6.399208e-08, 6.415348e-08, 6.426145e-08, 6.436783e-08, 
    6.468986e-08, 6.486028e-08, 6.524188e-08, 6.5173e-08, 6.528968e-08, 
    6.540112e-08, 6.558825e-08, 6.555744e-08, 6.563989e-08, 6.528659e-08, 
    6.55214e-08, 6.513378e-08, 6.52398e-08, 6.439678e-08, 6.407557e-08, 
    6.393907e-08, 6.381956e-08, 6.352884e-08, 6.372961e-08, 6.365047e-08, 
    6.383875e-08, 6.395839e-08, 6.389921e-08, 6.426441e-08, 6.412242e-08, 
    6.487038e-08, 6.454822e-08, 6.538812e-08, 6.518714e-08, 6.54363e-08, 
    6.530916e-08, 6.5527e-08, 6.533094e-08, 6.567057e-08, 6.574452e-08, 
    6.569399e-08, 6.588811e-08, 6.532007e-08, 6.553822e-08, 6.389756e-08, 
    6.390721e-08, 6.395216e-08, 6.375454e-08, 6.374245e-08, 6.356133e-08, 
    6.372249e-08, 6.379111e-08, 6.396532e-08, 6.406837e-08, 6.416632e-08, 
    6.438169e-08, 6.462222e-08, 6.495855e-08, 6.520017e-08, 6.536213e-08, 
    6.526282e-08, 6.53505e-08, 6.525248e-08, 6.520654e-08, 6.571682e-08, 
    6.543029e-08, 6.586019e-08, 6.58364e-08, 6.564185e-08, 6.583908e-08, 
    6.391399e-08, 6.385844e-08, 6.366564e-08, 6.381653e-08, 6.354161e-08, 
    6.36955e-08, 6.378399e-08, 6.41254e-08, 6.420041e-08, 6.426996e-08, 
    6.440733e-08, 6.458363e-08, 6.489289e-08, 6.516198e-08, 6.54076e-08, 
    6.538961e-08, 6.539594e-08, 6.545082e-08, 6.531489e-08, 6.547314e-08, 
    6.54997e-08, 6.543026e-08, 6.583321e-08, 6.571809e-08, 6.58359e-08, 
    6.576094e-08, 6.38765e-08, 6.396994e-08, 6.391945e-08, 6.40144e-08, 
    6.394751e-08, 6.424496e-08, 6.433414e-08, 6.475143e-08, 6.458016e-08, 
    6.485271e-08, 6.460785e-08, 6.465124e-08, 6.486162e-08, 6.462108e-08, 
    6.514714e-08, 6.47905e-08, 6.545295e-08, 6.509682e-08, 6.547527e-08, 
    6.540655e-08, 6.552033e-08, 6.562224e-08, 6.575045e-08, 6.598701e-08, 
    6.593223e-08, 6.613006e-08, 6.410925e-08, 6.423046e-08, 6.421978e-08, 
    6.434662e-08, 6.444042e-08, 6.464373e-08, 6.496981e-08, 6.484719e-08, 
    6.507229e-08, 6.511748e-08, 6.477549e-08, 6.498548e-08, 6.431157e-08, 
    6.442045e-08, 6.435562e-08, 6.411882e-08, 6.487545e-08, 6.448715e-08, 
    6.520416e-08, 6.499381e-08, 6.560771e-08, 6.530242e-08, 6.590207e-08, 
    6.615844e-08, 6.639969e-08, 6.668164e-08, 6.42966e-08, 6.421424e-08, 
    6.43617e-08, 6.456572e-08, 6.4755e-08, 6.500665e-08, 6.503239e-08, 
    6.507953e-08, 6.520164e-08, 6.530431e-08, 6.509445e-08, 6.533005e-08, 
    6.444572e-08, 6.490915e-08, 6.418311e-08, 6.440175e-08, 6.455369e-08, 
    6.448703e-08, 6.483317e-08, 6.491475e-08, 6.524627e-08, 6.507489e-08, 
    6.609517e-08, 6.564377e-08, 6.689631e-08, 6.654629e-08, 6.418547e-08, 
    6.429631e-08, 6.468208e-08, 6.449854e-08, 6.502344e-08, 6.515264e-08, 
    6.525767e-08, 6.539194e-08, 6.540643e-08, 6.548598e-08, 6.535562e-08, 
    6.548083e-08, 6.500718e-08, 6.521884e-08, 6.463799e-08, 6.477936e-08, 
    6.471433e-08, 6.464298e-08, 6.486317e-08, 6.509775e-08, 6.510275e-08, 
    6.517797e-08, 6.538995e-08, 6.502557e-08, 6.615345e-08, 6.545692e-08, 
    6.441718e-08, 6.463069e-08, 6.466117e-08, 6.457847e-08, 6.513969e-08, 
    6.493634e-08, 6.548404e-08, 6.533602e-08, 6.557855e-08, 6.545803e-08, 
    6.54403e-08, 6.528551e-08, 6.518914e-08, 6.494567e-08, 6.474756e-08, 
    6.459047e-08, 6.4627e-08, 6.479956e-08, 6.51121e-08, 6.540775e-08, 
    6.534299e-08, 6.556012e-08, 6.498538e-08, 6.522639e-08, 6.513324e-08, 
    6.537611e-08, 6.484393e-08, 6.529714e-08, 6.472809e-08, 6.477798e-08, 
    6.493231e-08, 6.524274e-08, 6.53114e-08, 6.538474e-08, 6.533948e-08, 
    6.512003e-08, 6.508407e-08, 6.492856e-08, 6.488562e-08, 6.476711e-08, 
    6.466901e-08, 6.475865e-08, 6.485278e-08, 6.512012e-08, 6.536104e-08, 
    6.562369e-08, 6.568797e-08, 6.599488e-08, 6.574506e-08, 6.615733e-08, 
    6.580684e-08, 6.641355e-08, 6.532339e-08, 6.579651e-08, 6.493933e-08, 
    6.503167e-08, 6.519871e-08, 6.558179e-08, 6.537497e-08, 6.561685e-08, 
    6.508266e-08, 6.480552e-08, 6.47338e-08, 6.460002e-08, 6.473686e-08, 
    6.472573e-08, 6.485668e-08, 6.48146e-08, 6.512899e-08, 6.496011e-08, 
    6.543986e-08, 6.561493e-08, 6.610933e-08, 6.641241e-08, 6.672092e-08, 
    6.685712e-08, 6.689857e-08, 6.69159e-08 ;

 STORVEGC =
  0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 0.7217537, 
    0.7217537, 0.7217537 ;

 STORVEGN =
  0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 0.0288706, 
    0.0288706, 0.0288706 ;

 SUPPLEMENT_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SoilAlpha =
  0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999944, 0.9999943, 
    0.9999943, 0.9999943, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999943, 0.9999942, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999942, 0.9999943, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999943, 0.9999942, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999943, 0.9999942, 0.9999943, 0.9999942, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999944, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999942, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999942, 0.9999942, 0.9999942, 0.9999942, 
    0.9999943, 0.9999942, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999944, 0.9999944, 0.9999944, 0.9999942, 0.9999942, 
    0.9999942, 0.9999942, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999942, 0.9999943, 
    0.9999942, 0.9999942, 0.9999942, 0.9999942, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999944, 0.9999943, 0.9999945, 0.9999944, 
    0.9999942, 0.9999942, 0.9999943, 0.9999942, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999944, 0.9999943, 0.9999942, 0.9999943, 0.9999943, 0.9999942, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999942, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999944, 0.9999943, 0.9999944, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999942, 
    0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 0.9999943, 
    0.9999943, 0.9999943, 0.9999944, 0.9999944, 0.9999944, 0.9999945, 
    0.9999945, 0.9999945 ;

 SoilAlpha_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TAUX =
  -0.1478002, -0.1478152, -0.1478124, -0.1478243, -0.1478178, -0.1478255, 
    -0.1478034, -0.1478157, -0.1478079, -0.1478017, -0.1478458, -0.1478249, 
    -0.1478621, -0.1478534, -0.1478862, -0.1478606, -0.147889, -0.1478859, 
    -0.1478956, -0.1478929, -0.1479049, -0.1478969, -0.1479115, -0.1479031, 
    -0.1479044, -0.1478966, -0.1478294, -0.1478432, -0.1478286, -0.1478305, 
    -0.1478297, -0.1478178, -0.1478115, -0.1477992, -0.1478015, -0.1478107, 
    -0.1478314, -0.1478248, -0.1478418, -0.1478415, -0.1478567, -0.1478509, 
    -0.1478826, -0.1478657, -0.147893, -0.147889, -0.1478928, -0.1478917, 
    -0.1478928, -0.1478869, -0.1478894, -0.1478843, -0.147852, -0.1478584, 
    -0.1478341, -0.1478157, -0.1478038, -0.1477952, -0.1477964, -0.1477987, 
    -0.1478107, -0.1478222, -0.1478307, -0.147836, -0.1478414, -0.1478546, 
    -0.1478603, -0.1478836, -0.1478816, -0.1478851, -0.1478886, -0.1478943, 
    -0.1478934, -0.1478959, -0.1478851, -0.1478922, -0.1478804, -0.1478837, 
    -0.147842, -0.1478267, -0.147819, -0.1478129, -0.1477973, -0.147808, 
    -0.1478038, -0.147814, -0.1478204, -0.1478173, -0.1478362, -0.1478291, 
    -0.1478606, -0.1478499, -0.1478882, -0.147882, -0.1478897, -0.1478858, 
    -0.1478924, -0.1478865, -0.1478968, -0.147899, -0.1478975, -0.1479035, 
    -0.1478861, -0.1478927, -0.1478172, -0.1478177, -0.1478201, -0.1478093, 
    -0.1478087, -0.1477991, -0.1478077, -0.1478114, -0.1478208, -0.1478263, 
    -0.1478312, -0.147842, -0.1478525, -0.1478635, -0.1478824, -0.1478874, 
    -0.1478844, -0.1478871, -0.1478841, -0.1478827, -0.1478982, -0.1478894, 
    -0.1479026, -0.1479019, -0.1478959, -0.147902, -0.147818, -0.1478151, 
    -0.1478047, -0.1478128, -0.1477981, -0.1478062, -0.1478108, -0.147829, 
    -0.147833, -0.1478364, -0.1478433, -0.1478512, -0.1478614, -0.1478812, 
    -0.1478888, -0.1478883, -0.1478885, -0.1478901, -0.147886, -0.1478908, 
    -0.1478916, -0.1478895, -0.1479018, -0.1478983, -0.1479019, -0.1478996, 
    -0.1478161, -0.147821, -0.1478183, -0.1478234, -0.1478198, -0.147835, 
    -0.1478394, -0.1478567, -0.1478511, -0.1478601, -0.1478521, -0.1478536, 
    -0.1478601, -0.1478527, -0.1478806, -0.1478579, -0.1478902, -0.1478675, 
    -0.1478909, -0.1478888, -0.1478923, -0.1478953, -0.1478993, -0.1479064, 
    -0.1479048, -0.1479108, -0.1478284, -0.1478343, -0.147834, -0.1478403, 
    -0.1478449, -0.1478535, -0.147864, -0.1478601, -0.1478671, -0.1478799, 
    -0.1478578, -0.1478644, -0.1478384, -0.1478437, -0.1478407, -0.1478288, 
    -0.1478608, -0.1478471, -0.1478825, -0.1478647, -0.1478949, -0.1478854, 
    -0.1479039, -0.1479115, -0.1479191, -0.1479275, -0.1478378, -0.1478337, 
    -0.1478411, -0.1478504, -0.147857, -0.1478651, -0.1478659, -0.1478673, 
    -0.1478825, -0.1478857, -0.1478676, -0.1478865, -0.1478446, -0.1478619, 
    -0.147832, -0.1478427, -0.1478501, -0.1478473, -0.1478596, -0.1478623, 
    -0.1478838, -0.1478672, -0.1479095, -0.1478958, -0.1479342, -0.1479234, 
    -0.1478322, -0.1478378, -0.1478546, -0.1478478, -0.1478656, -0.147881, 
    -0.1478842, -0.1478883, -0.1478888, -0.1478912, -0.1478872, -0.147891, 
    -0.1478651, -0.147883, -0.1478533, -0.1478578, -0.1478558, -0.1478535, 
    -0.1478606, -0.1478677, -0.147868, -0.1478817, -0.1478876, -0.1478657, 
    -0.1479109, -0.1478898, -0.1478438, -0.1478528, -0.147854, -0.1478511, 
    -0.1478806, -0.1478629, -0.1478911, -0.1478866, -0.1478941, -0.1478903, 
    -0.1478898, -0.1478851, -0.1478821, -0.1478632, -0.1478568, -0.1478516, 
    -0.1478529, -0.1478584, -0.1478682, -0.1478887, -0.1478867, -0.1478935, 
    -0.1478645, -0.1478832, -0.1478803, -0.1478878, -0.1478599, -0.1478849, 
    -0.1478562, -0.1478578, -0.1478628, -0.1478835, -0.1478859, -0.147888, 
    -0.1478867, -0.1478799, -0.1478674, -0.1478627, -0.1478612, -0.1478575, 
    -0.1478543, -0.1478572, -0.1478601, -0.14788, -0.1478873, -0.1478954, 
    -0.1478974, -0.1479064, -0.1478988, -0.147911, -0.1479003, -0.147919, 
    -0.1478859, -0.1479003, -0.147863, -0.1478659, -0.1478822, -0.1478939, 
    -0.1478878, -0.147895, -0.1478674, -0.1478585, -0.1478564, -0.1478519, 
    -0.1478565, -0.1478561, -0.1478604, -0.147859, -0.1478802, -0.1478637, 
    -0.1478897, -0.147895, -0.1479101, -0.1479193, -0.1479289, -0.1479331, 
    -0.1479343, -0.1479349 ;

 TAUY =
  -0.1478002, -0.1478152, -0.1478124, -0.1478243, -0.1478178, -0.1478255, 
    -0.1478034, -0.1478157, -0.1478079, -0.1478017, -0.1478458, -0.1478249, 
    -0.1478621, -0.1478534, -0.1478862, -0.1478606, -0.147889, -0.1478859, 
    -0.1478956, -0.1478929, -0.1479049, -0.1478969, -0.1479115, -0.1479031, 
    -0.1479044, -0.1478966, -0.1478294, -0.1478432, -0.1478286, -0.1478305, 
    -0.1478297, -0.1478178, -0.1478115, -0.1477992, -0.1478015, -0.1478107, 
    -0.1478314, -0.1478248, -0.1478418, -0.1478415, -0.1478567, -0.1478509, 
    -0.1478826, -0.1478657, -0.147893, -0.147889, -0.1478928, -0.1478917, 
    -0.1478928, -0.1478869, -0.1478894, -0.1478843, -0.147852, -0.1478584, 
    -0.1478341, -0.1478157, -0.1478038, -0.1477952, -0.1477964, -0.1477987, 
    -0.1478107, -0.1478222, -0.1478307, -0.147836, -0.1478414, -0.1478546, 
    -0.1478603, -0.1478836, -0.1478816, -0.1478851, -0.1478886, -0.1478943, 
    -0.1478934, -0.1478959, -0.1478851, -0.1478922, -0.1478804, -0.1478837, 
    -0.147842, -0.1478267, -0.147819, -0.1478129, -0.1477973, -0.147808, 
    -0.1478038, -0.147814, -0.1478204, -0.1478173, -0.1478362, -0.1478291, 
    -0.1478606, -0.1478499, -0.1478882, -0.147882, -0.1478897, -0.1478858, 
    -0.1478924, -0.1478865, -0.1478968, -0.147899, -0.1478975, -0.1479035, 
    -0.1478861, -0.1478927, -0.1478172, -0.1478177, -0.1478201, -0.1478093, 
    -0.1478087, -0.1477991, -0.1478077, -0.1478114, -0.1478208, -0.1478263, 
    -0.1478312, -0.147842, -0.1478525, -0.1478635, -0.1478824, -0.1478874, 
    -0.1478844, -0.1478871, -0.1478841, -0.1478827, -0.1478982, -0.1478894, 
    -0.1479026, -0.1479019, -0.1478959, -0.147902, -0.147818, -0.1478151, 
    -0.1478047, -0.1478128, -0.1477981, -0.1478062, -0.1478108, -0.147829, 
    -0.147833, -0.1478364, -0.1478433, -0.1478512, -0.1478614, -0.1478812, 
    -0.1478888, -0.1478883, -0.1478885, -0.1478901, -0.147886, -0.1478908, 
    -0.1478916, -0.1478895, -0.1479018, -0.1478983, -0.1479019, -0.1478996, 
    -0.1478161, -0.147821, -0.1478183, -0.1478234, -0.1478198, -0.147835, 
    -0.1478394, -0.1478567, -0.1478511, -0.1478601, -0.1478521, -0.1478536, 
    -0.1478601, -0.1478527, -0.1478806, -0.1478579, -0.1478902, -0.1478675, 
    -0.1478909, -0.1478888, -0.1478923, -0.1478953, -0.1478993, -0.1479064, 
    -0.1479048, -0.1479108, -0.1478284, -0.1478343, -0.147834, -0.1478403, 
    -0.1478449, -0.1478535, -0.147864, -0.1478601, -0.1478671, -0.1478799, 
    -0.1478578, -0.1478644, -0.1478384, -0.1478437, -0.1478407, -0.1478288, 
    -0.1478608, -0.1478471, -0.1478825, -0.1478647, -0.1478949, -0.1478854, 
    -0.1479039, -0.1479115, -0.1479191, -0.1479275, -0.1478378, -0.1478337, 
    -0.1478411, -0.1478504, -0.147857, -0.1478651, -0.1478659, -0.1478673, 
    -0.1478825, -0.1478857, -0.1478676, -0.1478865, -0.1478446, -0.1478619, 
    -0.147832, -0.1478427, -0.1478501, -0.1478473, -0.1478596, -0.1478623, 
    -0.1478838, -0.1478672, -0.1479095, -0.1478958, -0.1479342, -0.1479234, 
    -0.1478322, -0.1478378, -0.1478546, -0.1478478, -0.1478656, -0.147881, 
    -0.1478842, -0.1478883, -0.1478888, -0.1478912, -0.1478872, -0.147891, 
    -0.1478651, -0.147883, -0.1478533, -0.1478578, -0.1478558, -0.1478535, 
    -0.1478606, -0.1478677, -0.147868, -0.1478817, -0.1478876, -0.1478657, 
    -0.1479109, -0.1478898, -0.1478438, -0.1478528, -0.147854, -0.1478511, 
    -0.1478806, -0.1478629, -0.1478911, -0.1478866, -0.1478941, -0.1478903, 
    -0.1478898, -0.1478851, -0.1478821, -0.1478632, -0.1478568, -0.1478516, 
    -0.1478529, -0.1478584, -0.1478682, -0.1478887, -0.1478867, -0.1478935, 
    -0.1478645, -0.1478832, -0.1478803, -0.1478878, -0.1478599, -0.1478849, 
    -0.1478562, -0.1478578, -0.1478628, -0.1478835, -0.1478859, -0.147888, 
    -0.1478867, -0.1478799, -0.1478674, -0.1478627, -0.1478612, -0.1478575, 
    -0.1478543, -0.1478572, -0.1478601, -0.14788, -0.1478873, -0.1478954, 
    -0.1478974, -0.1479064, -0.1478988, -0.147911, -0.1479003, -0.147919, 
    -0.1478859, -0.1479003, -0.147863, -0.1478659, -0.1478822, -0.1478939, 
    -0.1478878, -0.147895, -0.1478674, -0.1478585, -0.1478564, -0.1478519, 
    -0.1478565, -0.1478561, -0.1478604, -0.147859, -0.1478802, -0.1478637, 
    -0.1478897, -0.147895, -0.1479101, -0.1479193, -0.1479289, -0.1479331, 
    -0.1479343, -0.1479349 ;

 TBOT =
  256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044 ;

 TBUILD =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TG =
  261.6477, 261.6642, 261.661, 261.6743, 261.6669, 261.6756, 261.651, 
    261.6648, 261.656, 261.6492, 261.7, 261.6749, 261.7263, 261.7102, 
    261.7506, 261.7238, 261.7561, 261.7499, 261.7686, 261.7632, 261.787, 
    261.7711, 261.7994, 261.7832, 261.7858, 261.7705, 261.68, 261.6968, 
    261.679, 261.6814, 261.6803, 261.6671, 261.6603, 261.6464, 261.649, 
    261.6592, 261.6824, 261.6746, 261.6945, 261.694, 261.7162, 261.7062, 
    261.7434, 261.7329, 261.7635, 261.7557, 261.7631, 261.7609, 261.7631, 
    261.7518, 261.7567, 261.7467, 261.7081, 261.7195, 261.6855, 261.6651, 
    261.6516, 261.6421, 261.6434, 261.646, 261.6593, 261.6718, 261.6813, 
    261.6877, 261.694, 261.7129, 261.723, 261.7455, 261.7415, 261.7484, 
    261.755, 261.7661, 261.7642, 261.7691, 261.7482, 261.7621, 261.7392, 
    261.7454, 261.6955, 261.6767, 261.6686, 261.6616, 261.6444, 261.6563, 
    261.6516, 261.6628, 261.6698, 261.6663, 261.6879, 261.6795, 261.7236, 
    261.7046, 261.7542, 261.7423, 261.757, 261.7495, 261.7624, 261.7508, 
    261.7709, 261.7753, 261.7723, 261.7838, 261.7502, 261.7631, 261.6662, 
    261.6668, 261.6694, 261.6577, 261.657, 261.6464, 261.6559, 261.6599, 
    261.6702, 261.6763, 261.6821, 261.6948, 261.709, 261.7289, 261.7431, 
    261.7527, 261.7468, 261.752, 261.7462, 261.7435, 261.7736, 261.7567, 
    261.7821, 261.7807, 261.7692, 261.7809, 261.6672, 261.6639, 261.6525, 
    261.6614, 261.6452, 261.6543, 261.6595, 261.6796, 261.6841, 261.6882, 
    261.6963, 261.7067, 261.725, 261.7408, 261.7554, 261.7543, 261.7547, 
    261.7579, 261.7499, 261.7592, 261.7608, 261.7567, 261.7805, 261.7737, 
    261.7807, 261.7763, 261.665, 261.6705, 261.6675, 261.6731, 261.6691, 
    261.6867, 261.6919, 261.7166, 261.7065, 261.7226, 261.7081, 261.7107, 
    261.7231, 261.7089, 261.7399, 261.7189, 261.7581, 261.737, 261.7594, 
    261.7553, 261.7621, 261.7681, 261.7757, 261.7896, 261.7864, 261.7981, 
    261.6787, 261.6858, 261.6852, 261.6927, 261.6982, 261.7103, 261.7296, 
    261.7223, 261.7357, 261.7382, 261.7181, 261.7305, 261.6906, 261.697, 
    261.6932, 261.6792, 261.7239, 261.701, 261.7433, 261.731, 261.7672, 
    261.7491, 261.7846, 261.7997, 261.8141, 261.8306, 261.6898, 261.6849, 
    261.6936, 261.7056, 261.7169, 261.7318, 261.7333, 261.7361, 261.7432, 
    261.7493, 261.7369, 261.7508, 261.6985, 261.726, 261.683, 261.6959, 
    261.7049, 261.701, 261.7215, 261.7263, 261.7458, 261.7358, 261.796, 
    261.7693, 261.8434, 261.8227, 261.6832, 261.6898, 261.7125, 261.7017, 
    261.7328, 261.7403, 261.7465, 261.7544, 261.7553, 261.76, 261.7523, 
    261.7597, 261.7318, 261.7442, 261.7099, 261.7183, 261.7144, 261.7102, 
    261.7233, 261.7371, 261.7375, 261.7418, 261.7542, 261.7329, 261.7993, 
    261.7581, 261.6969, 261.7094, 261.7113, 261.7064, 261.7395, 261.7276, 
    261.7599, 261.7511, 261.7655, 261.7584, 261.7573, 261.7481, 261.7424, 
    261.7281, 261.7164, 261.7071, 261.7093, 261.7195, 261.738, 261.7553, 
    261.7515, 261.7644, 261.7305, 261.7446, 261.7391, 261.7535, 261.7221, 
    261.7487, 261.7153, 261.7182, 261.7274, 261.7455, 261.7497, 261.754, 
    261.7513, 261.7383, 261.7363, 261.7271, 261.7246, 261.7176, 261.7118, 
    261.7171, 261.7226, 261.7383, 261.7526, 261.7681, 261.772, 261.79, 
    261.7752, 261.7995, 261.7788, 261.8147, 261.7503, 261.7783, 261.7278, 
    261.7332, 261.743, 261.7656, 261.7534, 261.7677, 261.7362, 261.7198, 
    261.7156, 261.7077, 261.7158, 261.7151, 261.7229, 261.7204, 261.7389, 
    261.729, 261.7573, 261.7676, 261.7968, 261.8148, 261.833, 261.8411, 
    261.8435, 261.8445 ;

 TG_R =
  261.6477, 261.6642, 261.661, 261.6743, 261.6669, 261.6756, 261.651, 
    261.6648, 261.656, 261.6492, 261.7, 261.6749, 261.7263, 261.7102, 
    261.7506, 261.7238, 261.7561, 261.7499, 261.7686, 261.7632, 261.787, 
    261.7711, 261.7994, 261.7832, 261.7858, 261.7705, 261.68, 261.6968, 
    261.679, 261.6814, 261.6803, 261.6671, 261.6603, 261.6464, 261.649, 
    261.6592, 261.6824, 261.6746, 261.6945, 261.694, 261.7162, 261.7062, 
    261.7434, 261.7329, 261.7635, 261.7557, 261.7631, 261.7609, 261.7631, 
    261.7518, 261.7567, 261.7467, 261.7081, 261.7195, 261.6855, 261.6651, 
    261.6516, 261.6421, 261.6434, 261.646, 261.6593, 261.6718, 261.6813, 
    261.6877, 261.694, 261.7129, 261.723, 261.7455, 261.7415, 261.7484, 
    261.755, 261.7661, 261.7642, 261.7691, 261.7482, 261.7621, 261.7392, 
    261.7454, 261.6955, 261.6767, 261.6686, 261.6616, 261.6444, 261.6563, 
    261.6516, 261.6628, 261.6698, 261.6663, 261.6879, 261.6795, 261.7236, 
    261.7046, 261.7542, 261.7423, 261.757, 261.7495, 261.7624, 261.7508, 
    261.7709, 261.7753, 261.7723, 261.7838, 261.7502, 261.7631, 261.6662, 
    261.6668, 261.6694, 261.6577, 261.657, 261.6464, 261.6559, 261.6599, 
    261.6702, 261.6763, 261.6821, 261.6948, 261.709, 261.7289, 261.7431, 
    261.7527, 261.7468, 261.752, 261.7462, 261.7435, 261.7736, 261.7567, 
    261.7821, 261.7807, 261.7692, 261.7809, 261.6672, 261.6639, 261.6525, 
    261.6614, 261.6452, 261.6543, 261.6595, 261.6796, 261.6841, 261.6882, 
    261.6963, 261.7067, 261.725, 261.7408, 261.7554, 261.7543, 261.7547, 
    261.7579, 261.7499, 261.7592, 261.7608, 261.7567, 261.7805, 261.7737, 
    261.7807, 261.7763, 261.665, 261.6705, 261.6675, 261.6731, 261.6691, 
    261.6867, 261.6919, 261.7166, 261.7065, 261.7226, 261.7081, 261.7107, 
    261.7231, 261.7089, 261.7399, 261.7189, 261.7581, 261.737, 261.7594, 
    261.7553, 261.7621, 261.7681, 261.7757, 261.7896, 261.7864, 261.7981, 
    261.6787, 261.6858, 261.6852, 261.6927, 261.6982, 261.7103, 261.7296, 
    261.7223, 261.7357, 261.7382, 261.7181, 261.7305, 261.6906, 261.697, 
    261.6932, 261.6792, 261.7239, 261.701, 261.7433, 261.731, 261.7672, 
    261.7491, 261.7846, 261.7997, 261.8141, 261.8306, 261.6898, 261.6849, 
    261.6936, 261.7056, 261.7169, 261.7318, 261.7333, 261.7361, 261.7432, 
    261.7493, 261.7369, 261.7508, 261.6985, 261.726, 261.683, 261.6959, 
    261.7049, 261.701, 261.7215, 261.7263, 261.7458, 261.7358, 261.796, 
    261.7693, 261.8434, 261.8227, 261.6832, 261.6898, 261.7125, 261.7017, 
    261.7328, 261.7403, 261.7465, 261.7544, 261.7553, 261.76, 261.7523, 
    261.7597, 261.7318, 261.7442, 261.7099, 261.7183, 261.7144, 261.7102, 
    261.7233, 261.7371, 261.7375, 261.7418, 261.7542, 261.7329, 261.7993, 
    261.7581, 261.6969, 261.7094, 261.7113, 261.7064, 261.7395, 261.7276, 
    261.7599, 261.7511, 261.7655, 261.7584, 261.7573, 261.7481, 261.7424, 
    261.7281, 261.7164, 261.7071, 261.7093, 261.7195, 261.738, 261.7553, 
    261.7515, 261.7644, 261.7305, 261.7446, 261.7391, 261.7535, 261.7221, 
    261.7487, 261.7153, 261.7182, 261.7274, 261.7455, 261.7497, 261.754, 
    261.7513, 261.7383, 261.7363, 261.7271, 261.7246, 261.7176, 261.7118, 
    261.7171, 261.7226, 261.7383, 261.7526, 261.7681, 261.772, 261.79, 
    261.7752, 261.7995, 261.7788, 261.8147, 261.7503, 261.7783, 261.7278, 
    261.7332, 261.743, 261.7656, 261.7534, 261.7677, 261.7362, 261.7198, 
    261.7156, 261.7077, 261.7158, 261.7151, 261.7229, 261.7204, 261.7389, 
    261.729, 261.7573, 261.7676, 261.7968, 261.8148, 261.833, 261.8411, 
    261.8435, 261.8445 ;

 TG_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TH2OSFC =
  254.0223, 254.0242, 254.0238, 254.0253, 254.0245, 254.0254, 254.0227, 
    254.0242, 254.0233, 254.0225, 254.028, 254.0253, 254.031, 254.0293, 
    254.0337, 254.0307, 254.0343, 254.0336, 254.0357, 254.0351, 254.0377, 
    254.0359, 254.039, 254.0373, 254.0375, 254.0359, 254.0259, 254.0277, 
    254.0258, 254.0261, 254.026, 254.0245, 254.0237, 254.0222, 254.0225, 
    254.0236, 254.0262, 254.0253, 254.0275, 254.0275, 254.0299, 254.0288, 
    254.0329, 254.0318, 254.0351, 254.0343, 254.0351, 254.0348, 254.0351, 
    254.0338, 254.0343, 254.0333, 254.029, 254.0302, 254.0265, 254.0242, 
    254.0228, 254.0217, 254.0219, 254.0222, 254.0236, 254.025, 254.0261, 
    254.0268, 254.0275, 254.0295, 254.0306, 254.0331, 254.0327, 254.0334, 
    254.0342, 254.0354, 254.0352, 254.0357, 254.0334, 254.0349, 254.0324, 
    254.0331, 254.0275, 254.0256, 254.0246, 254.0239, 254.022, 254.0233, 
    254.0228, 254.024, 254.0248, 254.0244, 254.0268, 254.0259, 254.0307, 
    254.0286, 254.0341, 254.0328, 254.0344, 254.0336, 254.035, 254.0337, 
    254.0359, 254.0364, 254.0361, 254.0374, 254.0336, 254.035, 254.0244, 
    254.0245, 254.0248, 254.0235, 254.0234, 254.0222, 254.0233, 254.0237, 
    254.0248, 254.0255, 254.0262, 254.0275, 254.0291, 254.0313, 254.0329, 
    254.0339, 254.0333, 254.0338, 254.0332, 254.0329, 254.0362, 254.0343, 
    254.0372, 254.037, 254.0357, 254.037, 254.0245, 254.0242, 254.0229, 
    254.0239, 254.0221, 254.0231, 254.0236, 254.0259, 254.0264, 254.0268, 
    254.0277, 254.0289, 254.0309, 254.0326, 254.0342, 254.0341, 254.0341, 
    254.0345, 254.0336, 254.0346, 254.0348, 254.0344, 254.037, 254.0362, 
    254.037, 254.0365, 254.0243, 254.0249, 254.0245, 254.0251, 254.0247, 
    254.0266, 254.0272, 254.0299, 254.0288, 254.0306, 254.029, 254.0293, 
    254.0306, 254.0291, 254.0325, 254.0302, 254.0345, 254.0321, 254.0347, 
    254.0342, 254.035, 254.0356, 254.0365, 254.038, 254.0376, 254.0389, 
    254.0258, 254.0266, 254.0265, 254.0273, 254.0279, 254.0293, 254.0314, 
    254.0306, 254.032, 254.0323, 254.0301, 254.0315, 254.0271, 254.0278, 
    254.0274, 254.0258, 254.0307, 254.0282, 254.0329, 254.0315, 254.0355, 
    254.0335, 254.0374, 254.039, 254.0407, 254.0425, 254.027, 254.0265, 
    254.0274, 254.0287, 254.03, 254.0316, 254.0318, 254.0321, 254.0329, 
    254.0336, 254.0322, 254.0337, 254.0279, 254.031, 254.0262, 254.0276, 
    254.0287, 254.0282, 254.0305, 254.031, 254.0331, 254.0321, 254.0386, 
    254.0357, 254.0439, 254.0416, 254.0263, 254.027, 254.0295, 254.0283, 
    254.0317, 254.0325, 254.0332, 254.0341, 254.0342, 254.0347, 254.0339, 
    254.0347, 254.0316, 254.033, 254.0292, 254.0301, 254.0297, 254.0293, 
    254.0307, 254.0322, 254.0322, 254.0327, 254.034, 254.0317, 254.0389, 
    254.0344, 254.0278, 254.0291, 254.0294, 254.0288, 254.0325, 254.0312, 
    254.0347, 254.0338, 254.0353, 254.0345, 254.0344, 254.0334, 254.0328, 
    254.0312, 254.0299, 254.0289, 254.0292, 254.0303, 254.0323, 254.0342, 
    254.0338, 254.0352, 254.0315, 254.033, 254.0324, 254.034, 254.0305, 
    254.0334, 254.0298, 254.0301, 254.0311, 254.0331, 254.0336, 254.0341, 
    254.0338, 254.0323, 254.0321, 254.0311, 254.0308, 254.0301, 254.0294, 
    254.03, 254.0306, 254.0323, 254.0339, 254.0356, 254.036, 254.038, 
    254.0363, 254.039, 254.0367, 254.0407, 254.0336, 254.0367, 254.0312, 
    254.0318, 254.0328, 254.0353, 254.034, 254.0355, 254.0321, 254.0303, 
    254.0298, 254.029, 254.0299, 254.0298, 254.0307, 254.0304, 254.0324, 
    254.0313, 254.0344, 254.0355, 254.0388, 254.0407, 254.0428, 254.0437, 
    254.0439, 254.0441 ;

 THBOT =
  256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 256.2044, 
    256.2044, 256.2044 ;

 TKE1 =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TLAI =
  0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122, 0.001143122, 0.001143122, 
    0.001143122, 0.001143122, 0.001143122 ;

 TLAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TOTCOLC =
  18.24, 18.23998, 18.23999, 18.23998, 18.23998, 18.23997, 18.24, 18.23998, 
    18.23999, 18.24, 18.23996, 18.23998, 18.23993, 18.23995, 18.23991, 
    18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23988, 18.2399, 
    18.23987, 18.23989, 18.23988, 18.2399, 18.23997, 18.23996, 18.23997, 
    18.23997, 18.23997, 18.23998, 18.23999, 18.24, 18.24, 18.23999, 18.23997, 
    18.23998, 18.23996, 18.23996, 18.23994, 18.23995, 18.23992, 18.23993, 
    18.2399, 18.23991, 18.2399, 18.2399, 18.2399, 18.23991, 18.23991, 
    18.23992, 18.23995, 18.23994, 18.23997, 18.23998, 18.24, 18.24, 18.24, 
    18.24, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 18.23994, 
    18.23994, 18.23992, 18.23992, 18.23992, 18.23991, 18.2399, 18.2399, 
    18.2399, 18.23992, 18.2399, 18.23992, 18.23992, 18.23996, 18.23997, 
    18.23998, 18.23999, 18.24, 18.23999, 18.24, 18.23999, 18.23998, 18.23998, 
    18.23997, 18.23997, 18.23993, 18.23995, 18.23991, 18.23992, 18.23991, 
    18.23991, 18.2399, 18.23991, 18.2399, 18.23989, 18.23989, 18.23989, 
    18.23991, 18.2399, 18.23998, 18.23998, 18.23998, 18.23999, 18.23999, 
    18.24, 18.23999, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 
    18.23995, 18.23993, 18.23992, 18.23991, 18.23992, 18.23991, 18.23992, 
    18.23992, 18.23989, 18.23991, 18.23989, 18.23989, 18.2399, 18.23989, 
    18.23998, 18.23999, 18.24, 18.23999, 18.24, 18.23999, 18.23999, 18.23997, 
    18.23997, 18.23997, 18.23996, 18.23995, 18.23993, 18.23992, 18.23991, 
    18.23991, 18.23991, 18.23991, 18.23991, 18.23991, 18.2399, 18.23991, 
    18.23989, 18.23989, 18.23989, 18.23989, 18.23998, 18.23998, 18.23998, 
    18.23998, 18.23998, 18.23997, 18.23996, 18.23994, 18.23995, 18.23994, 
    18.23995, 18.23995, 18.23994, 18.23995, 18.23992, 18.23994, 18.23991, 
    18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23989, 18.23988, 
    18.23988, 18.23987, 18.23997, 18.23997, 18.23997, 18.23996, 18.23996, 
    18.23995, 18.23993, 18.23994, 18.23993, 18.23992, 18.23994, 18.23993, 
    18.23996, 18.23996, 18.23996, 18.23997, 18.23993, 18.23995, 18.23992, 
    18.23993, 18.2399, 18.23991, 18.23989, 18.23987, 18.23986, 18.23985, 
    18.23996, 18.23997, 18.23996, 18.23995, 18.23994, 18.23993, 18.23993, 
    18.23993, 18.23992, 18.23991, 18.23993, 18.23991, 18.23996, 18.23993, 
    18.23997, 18.23996, 18.23995, 18.23995, 18.23994, 18.23993, 18.23992, 
    18.23993, 18.23988, 18.2399, 18.23984, 18.23985, 18.23997, 18.23996, 
    18.23994, 18.23995, 18.23993, 18.23992, 18.23992, 18.23991, 18.23991, 
    18.23991, 18.23991, 18.23991, 18.23993, 18.23992, 18.23995, 18.23994, 
    18.23994, 18.23995, 18.23994, 18.23993, 18.23992, 18.23992, 18.23991, 
    18.23993, 18.23987, 18.23991, 18.23996, 18.23995, 18.23995, 18.23995, 
    18.23992, 18.23993, 18.23991, 18.23991, 18.2399, 18.23991, 18.23991, 
    18.23992, 18.23992, 18.23993, 18.23994, 18.23995, 18.23995, 18.23994, 
    18.23992, 18.23991, 18.23991, 18.2399, 18.23993, 18.23992, 18.23992, 
    18.23991, 18.23994, 18.23991, 18.23994, 18.23994, 18.23993, 18.23992, 
    18.23991, 18.23991, 18.23991, 18.23992, 18.23993, 18.23993, 18.23993, 
    18.23994, 18.23995, 18.23994, 18.23994, 18.23992, 18.23991, 18.2399, 
    18.23989, 18.23988, 18.23989, 18.23987, 18.23989, 18.23986, 18.23991, 
    18.23989, 18.23993, 18.23993, 18.23992, 18.2399, 18.23991, 18.2399, 
    18.23993, 18.23994, 18.23994, 18.23995, 18.23994, 18.23994, 18.23994, 
    18.23994, 18.23992, 18.23993, 18.23991, 18.2399, 18.23987, 18.23986, 
    18.23985, 18.23984, 18.23984, 18.23984 ;

 TOTCOLCH4 =
  1.383695e-05, 1.375052e-05, 1.37672e-05, 1.369838e-05, 1.373644e-05, 
    1.369155e-05, 1.381931e-05, 1.374711e-05, 1.379308e-05, 1.382912e-05, 
    1.356773e-05, 1.369534e-05, 1.35157e-05, 1.360669e-05, 1.338289e-05, 
    1.352968e-05, 1.335414e-05, 1.338706e-05, 1.328913e-05, 1.331685e-05, 
    1.319507e-05, 1.327642e-05, 1.313404e-05, 1.32143e-05, 1.320158e-05, 
    1.327914e-05, 1.366938e-05, 1.358341e-05, 1.367452e-05, 1.366215e-05, 
    1.36677e-05, 1.373564e-05, 1.377025e-05, 1.384364e-05, 1.383024e-05, 
    1.377638e-05, 1.36566e-05, 1.369692e-05, 1.359603e-05, 1.359829e-05, 
    1.357288e-05, 1.363001e-05, 1.342194e-05, 1.347973e-05, 1.331569e-05, 
    1.33561e-05, 1.331757e-05, 1.33292e-05, 1.331742e-05, 1.337692e-05, 
    1.335127e-05, 1.340418e-05, 1.361923e-05, 1.355453e-05, 1.364105e-05, 
    1.374541e-05, 1.381612e-05, 1.386693e-05, 1.385971e-05, 1.384598e-05, 
    1.377607e-05, 1.37113e-05, 1.366254e-05, 1.363022e-05, 1.359861e-05, 
    1.359106e-05, 1.35342e-05, 1.341038e-05, 1.343238e-05, 1.339521e-05, 
    1.336015e-05, 1.330218e-05, 1.331165e-05, 1.328639e-05, 1.33962e-05, 
    1.332275e-05, 1.344498e-05, 1.341105e-05, 1.358998e-05, 1.368601e-05, 
    1.372739e-05, 1.376399e-05, 1.385417e-05, 1.37917e-05, 1.381623e-05, 
    1.375811e-05, 1.372154e-05, 1.373959e-05, 1.362934e-05, 1.367188e-05, 
    1.353086e-05, 1.363912e-05, 1.336422e-05, 1.342786e-05, 1.334917e-05, 
    1.338907e-05, 1.332102e-05, 1.338219e-05, 1.327705e-05, 1.325464e-05, 
    1.326993e-05, 1.321168e-05, 1.338562e-05, 1.331756e-05, 1.37401e-05, 
    1.373715e-05, 1.372344e-05, 1.3784e-05, 1.378774e-05, 1.384401e-05, 
    1.379391e-05, 1.377273e-05, 1.371944e-05, 1.368819e-05, 1.365868e-05, 
    1.35945e-05, 1.361394e-05, 1.350186e-05, 1.342369e-05, 1.337238e-05, 
    1.340374e-05, 1.337604e-05, 1.340702e-05, 1.342166e-05, 1.326301e-05, 
    1.335103e-05, 1.321998e-05, 1.322708e-05, 1.328578e-05, 1.322628e-05, 
    1.373508e-05, 1.375207e-05, 1.381152e-05, 1.376493e-05, 1.385018e-05, 
    1.380226e-05, 1.377492e-05, 1.367097e-05, 1.364847e-05, 1.362768e-05, 
    1.358693e-05, 1.362706e-05, 1.352344e-05, 1.343591e-05, 1.335813e-05, 
    1.336376e-05, 1.336178e-05, 1.334464e-05, 1.338725e-05, 1.333771e-05, 
    1.332947e-05, 1.335105e-05, 1.322803e-05, 1.326264e-05, 1.322723e-05, 
    1.324971e-05, 1.374654e-05, 1.371802e-05, 1.373341e-05, 1.370452e-05, 
    1.372485e-05, 1.363512e-05, 1.360857e-05, 1.357042e-05, 1.362824e-05, 
    1.353672e-05, 1.361883e-05, 1.360413e-05, 1.353374e-05, 1.361435e-05, 
    1.344066e-05, 1.355737e-05, 1.334398e-05, 1.345685e-05, 1.333705e-05, 
    1.335846e-05, 1.33231e-05, 1.329178e-05, 1.325287e-05, 1.318244e-05, 
    1.319859e-05, 1.314073e-05, 1.367585e-05, 1.363946e-05, 1.364267e-05, 
    1.360489e-05, 1.357716e-05, 1.360668e-05, 1.349818e-05, 1.353856e-05, 
    1.346483e-05, 1.345022e-05, 1.356241e-05, 1.349305e-05, 1.361529e-05, 
    1.358303e-05, 1.360222e-05, 1.367296e-05, 1.352919e-05, 1.35634e-05, 
    1.342241e-05, 1.349034e-05, 1.329622e-05, 1.339118e-05, 1.320752e-05, 
    1.31325e-05, 1.306383e-05, 1.298569e-05, 1.361975e-05, 1.364433e-05, 
    1.360043e-05, 1.363314e-05, 1.356925e-05, 1.348615e-05, 1.347777e-05, 
    1.346248e-05, 1.342323e-05, 1.33906e-05, 1.345764e-05, 1.338248e-05, 
    1.357555e-05, 1.351808e-05, 1.365364e-05, 1.358855e-05, 1.363726e-05, 
    1.356345e-05, 1.354322e-05, 1.351625e-05, 1.340898e-05, 1.346399e-05, 
    1.315081e-05, 1.328518e-05, 1.292779e-05, 1.30229e-05, 1.365294e-05, 
    1.361984e-05, 1.359372e-05, 1.356007e-05, 1.348068e-05, 1.343891e-05, 
    1.340538e-05, 1.336302e-05, 1.335849e-05, 1.333372e-05, 1.337442e-05, 
    1.333532e-05, 1.348597e-05, 1.341773e-05, 1.360863e-05, 1.356111e-05, 
    1.358289e-05, 1.360694e-05, 1.353328e-05, 1.345657e-05, 1.345498e-05, 
    1.343078e-05, 1.336356e-05, 1.347999e-05, 1.313389e-05, 1.334267e-05, 
    1.358402e-05, 1.361107e-05, 1.360078e-05, 1.362883e-05, 1.344307e-05, 
    1.350915e-05, 1.333432e-05, 1.338059e-05, 1.330516e-05, 1.33424e-05, 
    1.334792e-05, 1.339655e-05, 1.342721e-05, 1.350609e-05, 1.357173e-05, 
    1.362475e-05, 1.361235e-05, 1.355437e-05, 1.345195e-05, 1.335807e-05, 
    1.337838e-05, 1.331083e-05, 1.349309e-05, 1.341532e-05, 1.344514e-05, 
    1.336799e-05, 1.353964e-05, 1.339279e-05, 1.357827e-05, 1.356158e-05, 
    1.351048e-05, 1.341009e-05, 1.338836e-05, 1.336527e-05, 1.33795e-05, 
    1.344939e-05, 1.346101e-05, 1.351172e-05, 1.352585e-05, 1.356521e-05, 
    1.359814e-05, 1.356803e-05, 1.35367e-05, 1.344937e-05, 1.337271e-05, 
    1.329133e-05, 1.327177e-05, 1.318009e-05, 1.325445e-05, 1.313276e-05, 
    1.323582e-05, 1.305986e-05, 1.338453e-05, 1.323897e-05, 1.350818e-05, 
    1.347801e-05, 1.342414e-05, 1.330414e-05, 1.336835e-05, 1.329341e-05, 
    1.346147e-05, 1.355238e-05, 1.357635e-05, 1.36215e-05, 1.357533e-05, 
    1.357906e-05, 1.353542e-05, 1.354939e-05, 1.344652e-05, 1.350136e-05, 
    1.334805e-05, 1.3294e-05, 1.314673e-05, 1.306022e-05, 1.297504e-05, 
    1.293828e-05, 1.29272e-05, 1.292258e-05 ;

 TOTCOLN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTECOSYSC =
  18.24, 18.23998, 18.23999, 18.23998, 18.23998, 18.23997, 18.24, 18.23998, 
    18.23999, 18.24, 18.23996, 18.23998, 18.23993, 18.23995, 18.23991, 
    18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23988, 18.2399, 
    18.23987, 18.23989, 18.23988, 18.2399, 18.23997, 18.23996, 18.23997, 
    18.23997, 18.23997, 18.23998, 18.23999, 18.24, 18.24, 18.23999, 18.23997, 
    18.23998, 18.23996, 18.23996, 18.23994, 18.23995, 18.23992, 18.23993, 
    18.2399, 18.23991, 18.2399, 18.2399, 18.2399, 18.23991, 18.23991, 
    18.23992, 18.23995, 18.23994, 18.23997, 18.23998, 18.24, 18.24, 18.24, 
    18.24, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 18.23994, 
    18.23994, 18.23992, 18.23992, 18.23992, 18.23991, 18.2399, 18.2399, 
    18.2399, 18.23992, 18.2399, 18.23992, 18.23992, 18.23996, 18.23997, 
    18.23998, 18.23999, 18.24, 18.23999, 18.24, 18.23999, 18.23998, 18.23998, 
    18.23997, 18.23997, 18.23993, 18.23995, 18.23991, 18.23992, 18.23991, 
    18.23991, 18.2399, 18.23991, 18.2399, 18.23989, 18.23989, 18.23989, 
    18.23991, 18.2399, 18.23998, 18.23998, 18.23998, 18.23999, 18.23999, 
    18.24, 18.23999, 18.23999, 18.23998, 18.23997, 18.23997, 18.23996, 
    18.23995, 18.23993, 18.23992, 18.23991, 18.23992, 18.23991, 18.23992, 
    18.23992, 18.23989, 18.23991, 18.23989, 18.23989, 18.2399, 18.23989, 
    18.23998, 18.23999, 18.24, 18.23999, 18.24, 18.23999, 18.23999, 18.23997, 
    18.23997, 18.23997, 18.23996, 18.23995, 18.23993, 18.23992, 18.23991, 
    18.23991, 18.23991, 18.23991, 18.23991, 18.23991, 18.2399, 18.23991, 
    18.23989, 18.23989, 18.23989, 18.23989, 18.23998, 18.23998, 18.23998, 
    18.23998, 18.23998, 18.23997, 18.23996, 18.23994, 18.23995, 18.23994, 
    18.23995, 18.23995, 18.23994, 18.23995, 18.23992, 18.23994, 18.23991, 
    18.23993, 18.23991, 18.23991, 18.2399, 18.2399, 18.23989, 18.23988, 
    18.23988, 18.23987, 18.23997, 18.23997, 18.23997, 18.23996, 18.23996, 
    18.23995, 18.23993, 18.23994, 18.23993, 18.23992, 18.23994, 18.23993, 
    18.23996, 18.23996, 18.23996, 18.23997, 18.23993, 18.23995, 18.23992, 
    18.23993, 18.2399, 18.23991, 18.23989, 18.23987, 18.23986, 18.23985, 
    18.23996, 18.23997, 18.23996, 18.23995, 18.23994, 18.23993, 18.23993, 
    18.23993, 18.23992, 18.23991, 18.23993, 18.23991, 18.23996, 18.23993, 
    18.23997, 18.23996, 18.23995, 18.23995, 18.23994, 18.23993, 18.23992, 
    18.23993, 18.23988, 18.2399, 18.23984, 18.23985, 18.23997, 18.23996, 
    18.23994, 18.23995, 18.23993, 18.23992, 18.23992, 18.23991, 18.23991, 
    18.23991, 18.23991, 18.23991, 18.23993, 18.23992, 18.23995, 18.23994, 
    18.23994, 18.23995, 18.23994, 18.23993, 18.23992, 18.23992, 18.23991, 
    18.23993, 18.23987, 18.23991, 18.23996, 18.23995, 18.23995, 18.23995, 
    18.23992, 18.23993, 18.23991, 18.23991, 18.2399, 18.23991, 18.23991, 
    18.23992, 18.23992, 18.23993, 18.23994, 18.23995, 18.23995, 18.23994, 
    18.23992, 18.23991, 18.23991, 18.2399, 18.23993, 18.23992, 18.23992, 
    18.23991, 18.23994, 18.23991, 18.23994, 18.23994, 18.23993, 18.23992, 
    18.23991, 18.23991, 18.23991, 18.23992, 18.23993, 18.23993, 18.23993, 
    18.23994, 18.23995, 18.23994, 18.23994, 18.23992, 18.23991, 18.2399, 
    18.23989, 18.23988, 18.23989, 18.23987, 18.23989, 18.23986, 18.23991, 
    18.23989, 18.23993, 18.23993, 18.23992, 18.2399, 18.23991, 18.2399, 
    18.23993, 18.23994, 18.23994, 18.23995, 18.23994, 18.23994, 18.23994, 
    18.23994, 18.23992, 18.23993, 18.23991, 18.2399, 18.23987, 18.23986, 
    18.23985, 18.23984, 18.23984, 18.23984 ;

 TOTECOSYSN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTLITC =
  6.210311e-05, 6.210295e-05, 6.210298e-05, 6.210285e-05, 6.210292e-05, 
    6.210284e-05, 6.210307e-05, 6.210294e-05, 6.210303e-05, 6.210309e-05, 
    6.21026e-05, 6.210284e-05, 6.210235e-05, 6.21025e-05, 6.210212e-05, 
    6.210238e-05, 6.210207e-05, 6.210212e-05, 6.210195e-05, 6.2102e-05, 
    6.210178e-05, 6.210193e-05, 6.210166e-05, 6.210181e-05, 6.210179e-05, 
    6.210194e-05, 6.210279e-05, 6.210263e-05, 6.21028e-05, 6.210278e-05, 
    6.210279e-05, 6.210292e-05, 6.210298e-05, 6.210311e-05, 6.210309e-05, 
    6.210299e-05, 6.210277e-05, 6.210284e-05, 6.210266e-05, 6.210266e-05, 
    6.210245e-05, 6.210255e-05, 6.210219e-05, 6.210229e-05, 6.2102e-05, 
    6.210207e-05, 6.2102e-05, 6.210202e-05, 6.2102e-05, 6.210211e-05, 
    6.210207e-05, 6.210216e-05, 6.210252e-05, 6.210242e-05, 6.210274e-05, 
    6.210294e-05, 6.210306e-05, 6.210316e-05, 6.210314e-05, 6.210312e-05, 
    6.210299e-05, 6.210287e-05, 6.210278e-05, 6.210272e-05, 6.210266e-05, 
    6.210248e-05, 6.210239e-05, 6.210217e-05, 6.21022e-05, 6.210214e-05, 
    6.210208e-05, 6.210197e-05, 6.210199e-05, 6.210194e-05, 6.210215e-05, 
    6.210202e-05, 6.210223e-05, 6.210217e-05, 6.210264e-05, 6.210282e-05, 
    6.21029e-05, 6.210297e-05, 6.210314e-05, 6.210302e-05, 6.210306e-05, 
    6.210296e-05, 6.210289e-05, 6.210292e-05, 6.210272e-05, 6.21028e-05, 
    6.210238e-05, 6.210256e-05, 6.210209e-05, 6.21022e-05, 6.210206e-05, 
    6.210213e-05, 6.210201e-05, 6.210212e-05, 6.210193e-05, 6.210188e-05, 
    6.210191e-05, 6.21018e-05, 6.210212e-05, 6.2102e-05, 6.210292e-05, 
    6.210292e-05, 6.21029e-05, 6.2103e-05, 6.210301e-05, 6.210311e-05, 
    6.210303e-05, 6.210298e-05, 6.210289e-05, 6.210283e-05, 6.210277e-05, 
    6.210266e-05, 6.210252e-05, 6.210233e-05, 6.210219e-05, 6.21021e-05, 
    6.210215e-05, 6.210211e-05, 6.210216e-05, 6.210219e-05, 6.21019e-05, 
    6.210207e-05, 6.210182e-05, 6.210183e-05, 6.210194e-05, 6.210183e-05, 
    6.210292e-05, 6.210295e-05, 6.210306e-05, 6.210297e-05, 6.210313e-05, 
    6.210304e-05, 6.210299e-05, 6.210279e-05, 6.210276e-05, 6.210271e-05, 
    6.210264e-05, 6.210254e-05, 6.210236e-05, 6.210221e-05, 6.210207e-05, 
    6.210209e-05, 6.210208e-05, 6.210205e-05, 6.210212e-05, 6.210204e-05, 
    6.210202e-05, 6.210207e-05, 6.210183e-05, 6.21019e-05, 6.210183e-05, 
    6.210188e-05, 6.210294e-05, 6.210289e-05, 6.210291e-05, 6.210286e-05, 
    6.21029e-05, 6.210273e-05, 6.210268e-05, 6.210244e-05, 6.210254e-05, 
    6.210239e-05, 6.210252e-05, 6.21025e-05, 6.210238e-05, 6.210252e-05, 
    6.210222e-05, 6.210242e-05, 6.210205e-05, 6.210225e-05, 6.210204e-05, 
    6.210207e-05, 6.210202e-05, 6.210196e-05, 6.210188e-05, 6.210175e-05, 
    6.210178e-05, 6.210167e-05, 6.210281e-05, 6.210274e-05, 6.210274e-05, 
    6.210267e-05, 6.210262e-05, 6.21025e-05, 6.210232e-05, 6.210239e-05, 
    6.210226e-05, 6.210224e-05, 6.210243e-05, 6.210231e-05, 6.210269e-05, 
    6.210263e-05, 6.210267e-05, 6.21028e-05, 6.210237e-05, 6.210259e-05, 
    6.210219e-05, 6.210231e-05, 6.210196e-05, 6.210213e-05, 6.21018e-05, 
    6.210165e-05, 6.210152e-05, 6.210136e-05, 6.21027e-05, 6.210275e-05, 
    6.210266e-05, 6.210255e-05, 6.210244e-05, 6.21023e-05, 6.210228e-05, 
    6.210226e-05, 6.210219e-05, 6.210213e-05, 6.210225e-05, 6.210212e-05, 
    6.210262e-05, 6.210236e-05, 6.210276e-05, 6.210264e-05, 6.210255e-05, 
    6.210259e-05, 6.21024e-05, 6.210235e-05, 6.210217e-05, 6.210226e-05, 
    6.210169e-05, 6.210194e-05, 6.210124e-05, 6.210144e-05, 6.210276e-05, 
    6.21027e-05, 6.210248e-05, 6.210259e-05, 6.210229e-05, 6.210222e-05, 
    6.210216e-05, 6.210208e-05, 6.210207e-05, 6.210203e-05, 6.21021e-05, 
    6.210204e-05, 6.21023e-05, 6.210218e-05, 6.210251e-05, 6.210243e-05, 
    6.210247e-05, 6.21025e-05, 6.210238e-05, 6.210225e-05, 6.210225e-05, 
    6.21022e-05, 6.210209e-05, 6.210229e-05, 6.210166e-05, 6.210204e-05, 
    6.210263e-05, 6.210251e-05, 6.21025e-05, 6.210254e-05, 6.210223e-05, 
    6.210234e-05, 6.210203e-05, 6.210212e-05, 6.210198e-05, 6.210204e-05, 
    6.210206e-05, 6.210215e-05, 6.21022e-05, 6.210234e-05, 6.210244e-05, 
    6.210253e-05, 6.210252e-05, 6.210242e-05, 6.210224e-05, 6.210207e-05, 
    6.210211e-05, 6.210199e-05, 6.210231e-05, 6.210218e-05, 6.210223e-05, 
    6.21021e-05, 6.210239e-05, 6.210214e-05, 6.210246e-05, 6.210243e-05, 
    6.210234e-05, 6.210217e-05, 6.210213e-05, 6.210209e-05, 6.210212e-05, 
    6.210223e-05, 6.210226e-05, 6.210234e-05, 6.210237e-05, 6.210244e-05, 
    6.210249e-05, 6.210244e-05, 6.210239e-05, 6.210223e-05, 6.21021e-05, 
    6.210196e-05, 6.210192e-05, 6.210175e-05, 6.210188e-05, 6.210166e-05, 
    6.210186e-05, 6.210151e-05, 6.210212e-05, 6.210186e-05, 6.210234e-05, 
    6.210228e-05, 6.210219e-05, 6.210198e-05, 6.21021e-05, 6.210196e-05, 
    6.210226e-05, 6.210242e-05, 6.210245e-05, 6.210253e-05, 6.210245e-05, 
    6.210246e-05, 6.210239e-05, 6.210241e-05, 6.210223e-05, 6.210233e-05, 
    6.210206e-05, 6.210196e-05, 6.210168e-05, 6.210151e-05, 6.210134e-05, 
    6.210127e-05, 6.210124e-05, 6.210123e-05 ;

 TOTLITC_1m =
  6.210311e-05, 6.210295e-05, 6.210298e-05, 6.210285e-05, 6.210292e-05, 
    6.210284e-05, 6.210307e-05, 6.210294e-05, 6.210303e-05, 6.210309e-05, 
    6.21026e-05, 6.210284e-05, 6.210235e-05, 6.21025e-05, 6.210212e-05, 
    6.210238e-05, 6.210207e-05, 6.210212e-05, 6.210195e-05, 6.2102e-05, 
    6.210178e-05, 6.210193e-05, 6.210166e-05, 6.210181e-05, 6.210179e-05, 
    6.210194e-05, 6.210279e-05, 6.210263e-05, 6.21028e-05, 6.210278e-05, 
    6.210279e-05, 6.210292e-05, 6.210298e-05, 6.210311e-05, 6.210309e-05, 
    6.210299e-05, 6.210277e-05, 6.210284e-05, 6.210266e-05, 6.210266e-05, 
    6.210245e-05, 6.210255e-05, 6.210219e-05, 6.210229e-05, 6.2102e-05, 
    6.210207e-05, 6.2102e-05, 6.210202e-05, 6.2102e-05, 6.210211e-05, 
    6.210207e-05, 6.210216e-05, 6.210252e-05, 6.210242e-05, 6.210274e-05, 
    6.210294e-05, 6.210306e-05, 6.210316e-05, 6.210314e-05, 6.210312e-05, 
    6.210299e-05, 6.210287e-05, 6.210278e-05, 6.210272e-05, 6.210266e-05, 
    6.210248e-05, 6.210239e-05, 6.210217e-05, 6.21022e-05, 6.210214e-05, 
    6.210208e-05, 6.210197e-05, 6.210199e-05, 6.210194e-05, 6.210215e-05, 
    6.210202e-05, 6.210223e-05, 6.210217e-05, 6.210264e-05, 6.210282e-05, 
    6.21029e-05, 6.210297e-05, 6.210314e-05, 6.210302e-05, 6.210306e-05, 
    6.210296e-05, 6.210289e-05, 6.210292e-05, 6.210272e-05, 6.21028e-05, 
    6.210238e-05, 6.210256e-05, 6.210209e-05, 6.21022e-05, 6.210206e-05, 
    6.210213e-05, 6.210201e-05, 6.210212e-05, 6.210193e-05, 6.210188e-05, 
    6.210191e-05, 6.21018e-05, 6.210212e-05, 6.2102e-05, 6.210292e-05, 
    6.210292e-05, 6.21029e-05, 6.2103e-05, 6.210301e-05, 6.210311e-05, 
    6.210303e-05, 6.210298e-05, 6.210289e-05, 6.210283e-05, 6.210277e-05, 
    6.210266e-05, 6.210252e-05, 6.210233e-05, 6.210219e-05, 6.21021e-05, 
    6.210215e-05, 6.210211e-05, 6.210216e-05, 6.210219e-05, 6.21019e-05, 
    6.210207e-05, 6.210182e-05, 6.210183e-05, 6.210194e-05, 6.210183e-05, 
    6.210292e-05, 6.210295e-05, 6.210306e-05, 6.210297e-05, 6.210313e-05, 
    6.210304e-05, 6.210299e-05, 6.210279e-05, 6.210276e-05, 6.210271e-05, 
    6.210264e-05, 6.210254e-05, 6.210236e-05, 6.210221e-05, 6.210207e-05, 
    6.210209e-05, 6.210208e-05, 6.210205e-05, 6.210212e-05, 6.210204e-05, 
    6.210202e-05, 6.210207e-05, 6.210183e-05, 6.21019e-05, 6.210183e-05, 
    6.210188e-05, 6.210294e-05, 6.210289e-05, 6.210291e-05, 6.210286e-05, 
    6.21029e-05, 6.210273e-05, 6.210268e-05, 6.210244e-05, 6.210254e-05, 
    6.210239e-05, 6.210252e-05, 6.21025e-05, 6.210238e-05, 6.210252e-05, 
    6.210222e-05, 6.210242e-05, 6.210205e-05, 6.210225e-05, 6.210204e-05, 
    6.210207e-05, 6.210202e-05, 6.210196e-05, 6.210188e-05, 6.210175e-05, 
    6.210178e-05, 6.210167e-05, 6.210281e-05, 6.210274e-05, 6.210274e-05, 
    6.210267e-05, 6.210262e-05, 6.21025e-05, 6.210232e-05, 6.210239e-05, 
    6.210226e-05, 6.210224e-05, 6.210243e-05, 6.210231e-05, 6.210269e-05, 
    6.210263e-05, 6.210267e-05, 6.21028e-05, 6.210237e-05, 6.210259e-05, 
    6.210219e-05, 6.210231e-05, 6.210196e-05, 6.210213e-05, 6.21018e-05, 
    6.210165e-05, 6.210152e-05, 6.210136e-05, 6.21027e-05, 6.210275e-05, 
    6.210266e-05, 6.210255e-05, 6.210244e-05, 6.21023e-05, 6.210228e-05, 
    6.210226e-05, 6.210219e-05, 6.210213e-05, 6.210225e-05, 6.210212e-05, 
    6.210262e-05, 6.210236e-05, 6.210276e-05, 6.210264e-05, 6.210255e-05, 
    6.210259e-05, 6.21024e-05, 6.210235e-05, 6.210217e-05, 6.210226e-05, 
    6.210169e-05, 6.210194e-05, 6.210124e-05, 6.210144e-05, 6.210276e-05, 
    6.21027e-05, 6.210248e-05, 6.210259e-05, 6.210229e-05, 6.210222e-05, 
    6.210216e-05, 6.210208e-05, 6.210207e-05, 6.210203e-05, 6.21021e-05, 
    6.210204e-05, 6.21023e-05, 6.210218e-05, 6.210251e-05, 6.210243e-05, 
    6.210247e-05, 6.21025e-05, 6.210238e-05, 6.210225e-05, 6.210225e-05, 
    6.21022e-05, 6.210209e-05, 6.210229e-05, 6.210166e-05, 6.210204e-05, 
    6.210263e-05, 6.210251e-05, 6.21025e-05, 6.210254e-05, 6.210223e-05, 
    6.210234e-05, 6.210203e-05, 6.210212e-05, 6.210198e-05, 6.210204e-05, 
    6.210206e-05, 6.210215e-05, 6.21022e-05, 6.210234e-05, 6.210244e-05, 
    6.210253e-05, 6.210252e-05, 6.210242e-05, 6.210224e-05, 6.210207e-05, 
    6.210211e-05, 6.210199e-05, 6.210231e-05, 6.210218e-05, 6.210223e-05, 
    6.21021e-05, 6.210239e-05, 6.210214e-05, 6.210246e-05, 6.210243e-05, 
    6.210234e-05, 6.210217e-05, 6.210213e-05, 6.210209e-05, 6.210212e-05, 
    6.210223e-05, 6.210226e-05, 6.210234e-05, 6.210237e-05, 6.210244e-05, 
    6.210249e-05, 6.210244e-05, 6.210239e-05, 6.210223e-05, 6.21021e-05, 
    6.210196e-05, 6.210192e-05, 6.210175e-05, 6.210188e-05, 6.210166e-05, 
    6.210186e-05, 6.210151e-05, 6.210212e-05, 6.210186e-05, 6.210234e-05, 
    6.210228e-05, 6.210219e-05, 6.210198e-05, 6.21021e-05, 6.210196e-05, 
    6.210226e-05, 6.210242e-05, 6.210245e-05, 6.210253e-05, 6.210245e-05, 
    6.210246e-05, 6.210239e-05, 6.210241e-05, 6.210223e-05, 6.210233e-05, 
    6.210206e-05, 6.210196e-05, 6.210168e-05, 6.210151e-05, 6.210134e-05, 
    6.210127e-05, 6.210124e-05, 6.210123e-05 ;

 TOTLITN =
  1.429818e-06, 1.429813e-06, 1.429814e-06, 1.429811e-06, 1.429813e-06, 
    1.42981e-06, 1.429817e-06, 1.429813e-06, 1.429816e-06, 1.429818e-06, 
    1.429804e-06, 1.429811e-06, 1.429797e-06, 1.429801e-06, 1.42979e-06, 
    1.429797e-06, 1.429789e-06, 1.42979e-06, 1.429785e-06, 1.429787e-06, 
    1.42978e-06, 1.429785e-06, 1.429777e-06, 1.429781e-06, 1.429781e-06, 
    1.429785e-06, 1.429809e-06, 1.429805e-06, 1.429809e-06, 1.429809e-06, 
    1.429809e-06, 1.429813e-06, 1.429814e-06, 1.429818e-06, 1.429818e-06, 
    1.429815e-06, 1.429809e-06, 1.429811e-06, 1.429805e-06, 1.429805e-06, 
    1.429799e-06, 1.429802e-06, 1.429792e-06, 1.429795e-06, 1.429787e-06, 
    1.429789e-06, 1.429787e-06, 1.429788e-06, 1.429787e-06, 1.42979e-06, 
    1.429789e-06, 1.429791e-06, 1.429802e-06, 1.429799e-06, 1.429808e-06, 
    1.429813e-06, 1.429817e-06, 1.429819e-06, 1.429819e-06, 1.429818e-06, 
    1.429815e-06, 1.429811e-06, 1.429809e-06, 1.429807e-06, 1.429805e-06, 
    1.4298e-06, 1.429798e-06, 1.429792e-06, 1.429793e-06, 1.429791e-06, 
    1.429789e-06, 1.429786e-06, 1.429787e-06, 1.429785e-06, 1.429791e-06, 
    1.429787e-06, 1.429793e-06, 1.429792e-06, 1.429805e-06, 1.42981e-06, 
    1.429812e-06, 1.429814e-06, 1.429819e-06, 1.429816e-06, 1.429817e-06, 
    1.429814e-06, 1.429812e-06, 1.429813e-06, 1.429807e-06, 1.429809e-06, 
    1.429798e-06, 1.429803e-06, 1.429789e-06, 1.429793e-06, 1.429789e-06, 
    1.429791e-06, 1.429787e-06, 1.42979e-06, 1.429785e-06, 1.429784e-06, 
    1.429784e-06, 1.429781e-06, 1.42979e-06, 1.429787e-06, 1.429813e-06, 
    1.429813e-06, 1.429812e-06, 1.429815e-06, 1.429815e-06, 1.429818e-06, 
    1.429816e-06, 1.429815e-06, 1.429812e-06, 1.42981e-06, 1.429809e-06, 
    1.429805e-06, 1.429801e-06, 1.429796e-06, 1.429792e-06, 1.42979e-06, 
    1.429791e-06, 1.42979e-06, 1.429791e-06, 1.429792e-06, 1.429784e-06, 
    1.429789e-06, 1.429782e-06, 1.429782e-06, 1.429785e-06, 1.429782e-06, 
    1.429813e-06, 1.429814e-06, 1.429817e-06, 1.429814e-06, 1.429819e-06, 
    1.429816e-06, 1.429815e-06, 1.429809e-06, 1.429808e-06, 1.429807e-06, 
    1.429805e-06, 1.429802e-06, 1.429797e-06, 1.429793e-06, 1.429789e-06, 
    1.429789e-06, 1.429789e-06, 1.429788e-06, 1.42979e-06, 1.429788e-06, 
    1.429788e-06, 1.429789e-06, 1.429782e-06, 1.429784e-06, 1.429782e-06, 
    1.429783e-06, 1.429813e-06, 1.429812e-06, 1.429813e-06, 1.429811e-06, 
    1.429812e-06, 1.429807e-06, 1.429806e-06, 1.429799e-06, 1.429802e-06, 
    1.429798e-06, 1.429802e-06, 1.429801e-06, 1.429798e-06, 1.429801e-06, 
    1.429793e-06, 1.429799e-06, 1.429788e-06, 1.429794e-06, 1.429788e-06, 
    1.429789e-06, 1.429787e-06, 1.429786e-06, 1.429784e-06, 1.42978e-06, 
    1.429781e-06, 1.429778e-06, 1.42981e-06, 1.429808e-06, 1.429808e-06, 
    1.429806e-06, 1.429804e-06, 1.429801e-06, 1.429796e-06, 1.429798e-06, 
    1.429794e-06, 1.429794e-06, 1.429799e-06, 1.429796e-06, 1.429806e-06, 
    1.429805e-06, 1.429806e-06, 1.429809e-06, 1.429797e-06, 1.429804e-06, 
    1.429792e-06, 1.429796e-06, 1.429786e-06, 1.429791e-06, 1.429781e-06, 
    1.429777e-06, 1.429773e-06, 1.429769e-06, 1.429807e-06, 1.429808e-06, 
    1.429806e-06, 1.429802e-06, 1.429799e-06, 1.429795e-06, 1.429795e-06, 
    1.429794e-06, 1.429792e-06, 1.429791e-06, 1.429794e-06, 1.42979e-06, 
    1.429804e-06, 1.429797e-06, 1.429808e-06, 1.429805e-06, 1.429803e-06, 
    1.429804e-06, 1.429798e-06, 1.429797e-06, 1.429791e-06, 1.429794e-06, 
    1.429778e-06, 1.429785e-06, 1.429766e-06, 1.429771e-06, 1.429808e-06, 
    1.429807e-06, 1.4298e-06, 1.429803e-06, 1.429795e-06, 1.429793e-06, 
    1.429791e-06, 1.429789e-06, 1.429789e-06, 1.429788e-06, 1.42979e-06, 
    1.429788e-06, 1.429795e-06, 1.429792e-06, 1.429801e-06, 1.429799e-06, 
    1.4298e-06, 1.429801e-06, 1.429798e-06, 1.429794e-06, 1.429794e-06, 
    1.429793e-06, 1.429789e-06, 1.429795e-06, 1.429777e-06, 1.429788e-06, 
    1.429805e-06, 1.429801e-06, 1.429801e-06, 1.429802e-06, 1.429793e-06, 
    1.429796e-06, 1.429788e-06, 1.42979e-06, 1.429786e-06, 1.429788e-06, 
    1.429788e-06, 1.429791e-06, 1.429792e-06, 1.429796e-06, 1.429799e-06, 
    1.429802e-06, 1.429801e-06, 1.429799e-06, 1.429794e-06, 1.429789e-06, 
    1.42979e-06, 1.429787e-06, 1.429796e-06, 1.429792e-06, 1.429793e-06, 
    1.429789e-06, 1.429798e-06, 1.429791e-06, 1.4298e-06, 1.429799e-06, 
    1.429796e-06, 1.429792e-06, 1.42979e-06, 1.429789e-06, 1.42979e-06, 
    1.429794e-06, 1.429794e-06, 1.429797e-06, 1.429797e-06, 1.429799e-06, 
    1.429801e-06, 1.429799e-06, 1.429798e-06, 1.429794e-06, 1.42979e-06, 
    1.429786e-06, 1.429785e-06, 1.42978e-06, 1.429784e-06, 1.429777e-06, 
    1.429783e-06, 1.429773e-06, 1.42979e-06, 1.429783e-06, 1.429796e-06, 
    1.429795e-06, 1.429792e-06, 1.429786e-06, 1.429789e-06, 1.429786e-06, 
    1.429794e-06, 1.429799e-06, 1.4298e-06, 1.429802e-06, 1.4298e-06, 
    1.4298e-06, 1.429798e-06, 1.429798e-06, 1.429793e-06, 1.429796e-06, 
    1.429788e-06, 1.429786e-06, 1.429778e-06, 1.429773e-06, 1.429768e-06, 
    1.429766e-06, 1.429765e-06, 1.429765e-06 ;

 TOTLITN_1m =
  1.429818e-06, 1.429813e-06, 1.429814e-06, 1.429811e-06, 1.429813e-06, 
    1.42981e-06, 1.429817e-06, 1.429813e-06, 1.429816e-06, 1.429818e-06, 
    1.429804e-06, 1.429811e-06, 1.429797e-06, 1.429801e-06, 1.42979e-06, 
    1.429797e-06, 1.429789e-06, 1.42979e-06, 1.429785e-06, 1.429787e-06, 
    1.42978e-06, 1.429785e-06, 1.429777e-06, 1.429781e-06, 1.429781e-06, 
    1.429785e-06, 1.429809e-06, 1.429805e-06, 1.429809e-06, 1.429809e-06, 
    1.429809e-06, 1.429813e-06, 1.429814e-06, 1.429818e-06, 1.429818e-06, 
    1.429815e-06, 1.429809e-06, 1.429811e-06, 1.429805e-06, 1.429805e-06, 
    1.429799e-06, 1.429802e-06, 1.429792e-06, 1.429795e-06, 1.429787e-06, 
    1.429789e-06, 1.429787e-06, 1.429788e-06, 1.429787e-06, 1.42979e-06, 
    1.429789e-06, 1.429791e-06, 1.429802e-06, 1.429799e-06, 1.429808e-06, 
    1.429813e-06, 1.429817e-06, 1.429819e-06, 1.429819e-06, 1.429818e-06, 
    1.429815e-06, 1.429811e-06, 1.429809e-06, 1.429807e-06, 1.429805e-06, 
    1.4298e-06, 1.429798e-06, 1.429792e-06, 1.429793e-06, 1.429791e-06, 
    1.429789e-06, 1.429786e-06, 1.429787e-06, 1.429785e-06, 1.429791e-06, 
    1.429787e-06, 1.429793e-06, 1.429792e-06, 1.429805e-06, 1.42981e-06, 
    1.429812e-06, 1.429814e-06, 1.429819e-06, 1.429816e-06, 1.429817e-06, 
    1.429814e-06, 1.429812e-06, 1.429813e-06, 1.429807e-06, 1.429809e-06, 
    1.429798e-06, 1.429803e-06, 1.429789e-06, 1.429793e-06, 1.429789e-06, 
    1.429791e-06, 1.429787e-06, 1.42979e-06, 1.429785e-06, 1.429784e-06, 
    1.429784e-06, 1.429781e-06, 1.42979e-06, 1.429787e-06, 1.429813e-06, 
    1.429813e-06, 1.429812e-06, 1.429815e-06, 1.429815e-06, 1.429818e-06, 
    1.429816e-06, 1.429815e-06, 1.429812e-06, 1.42981e-06, 1.429809e-06, 
    1.429805e-06, 1.429801e-06, 1.429796e-06, 1.429792e-06, 1.42979e-06, 
    1.429791e-06, 1.42979e-06, 1.429791e-06, 1.429792e-06, 1.429784e-06, 
    1.429789e-06, 1.429782e-06, 1.429782e-06, 1.429785e-06, 1.429782e-06, 
    1.429813e-06, 1.429814e-06, 1.429817e-06, 1.429814e-06, 1.429819e-06, 
    1.429816e-06, 1.429815e-06, 1.429809e-06, 1.429808e-06, 1.429807e-06, 
    1.429805e-06, 1.429802e-06, 1.429797e-06, 1.429793e-06, 1.429789e-06, 
    1.429789e-06, 1.429789e-06, 1.429788e-06, 1.42979e-06, 1.429788e-06, 
    1.429788e-06, 1.429789e-06, 1.429782e-06, 1.429784e-06, 1.429782e-06, 
    1.429783e-06, 1.429813e-06, 1.429812e-06, 1.429813e-06, 1.429811e-06, 
    1.429812e-06, 1.429807e-06, 1.429806e-06, 1.429799e-06, 1.429802e-06, 
    1.429798e-06, 1.429802e-06, 1.429801e-06, 1.429798e-06, 1.429801e-06, 
    1.429793e-06, 1.429799e-06, 1.429788e-06, 1.429794e-06, 1.429788e-06, 
    1.429789e-06, 1.429787e-06, 1.429786e-06, 1.429784e-06, 1.42978e-06, 
    1.429781e-06, 1.429778e-06, 1.42981e-06, 1.429808e-06, 1.429808e-06, 
    1.429806e-06, 1.429804e-06, 1.429801e-06, 1.429796e-06, 1.429798e-06, 
    1.429794e-06, 1.429794e-06, 1.429799e-06, 1.429796e-06, 1.429806e-06, 
    1.429805e-06, 1.429806e-06, 1.429809e-06, 1.429797e-06, 1.429804e-06, 
    1.429792e-06, 1.429796e-06, 1.429786e-06, 1.429791e-06, 1.429781e-06, 
    1.429777e-06, 1.429773e-06, 1.429769e-06, 1.429807e-06, 1.429808e-06, 
    1.429806e-06, 1.429802e-06, 1.429799e-06, 1.429795e-06, 1.429795e-06, 
    1.429794e-06, 1.429792e-06, 1.429791e-06, 1.429794e-06, 1.42979e-06, 
    1.429804e-06, 1.429797e-06, 1.429808e-06, 1.429805e-06, 1.429803e-06, 
    1.429804e-06, 1.429798e-06, 1.429797e-06, 1.429791e-06, 1.429794e-06, 
    1.429778e-06, 1.429785e-06, 1.429766e-06, 1.429771e-06, 1.429808e-06, 
    1.429807e-06, 1.4298e-06, 1.429803e-06, 1.429795e-06, 1.429793e-06, 
    1.429791e-06, 1.429789e-06, 1.429789e-06, 1.429788e-06, 1.42979e-06, 
    1.429788e-06, 1.429795e-06, 1.429792e-06, 1.429801e-06, 1.429799e-06, 
    1.4298e-06, 1.429801e-06, 1.429798e-06, 1.429794e-06, 1.429794e-06, 
    1.429793e-06, 1.429789e-06, 1.429795e-06, 1.429777e-06, 1.429788e-06, 
    1.429805e-06, 1.429801e-06, 1.429801e-06, 1.429802e-06, 1.429793e-06, 
    1.429796e-06, 1.429788e-06, 1.42979e-06, 1.429786e-06, 1.429788e-06, 
    1.429788e-06, 1.429791e-06, 1.429792e-06, 1.429796e-06, 1.429799e-06, 
    1.429802e-06, 1.429801e-06, 1.429799e-06, 1.429794e-06, 1.429789e-06, 
    1.42979e-06, 1.429787e-06, 1.429796e-06, 1.429792e-06, 1.429793e-06, 
    1.429789e-06, 1.429798e-06, 1.429791e-06, 1.4298e-06, 1.429799e-06, 
    1.429796e-06, 1.429792e-06, 1.42979e-06, 1.429789e-06, 1.42979e-06, 
    1.429794e-06, 1.429794e-06, 1.429797e-06, 1.429797e-06, 1.429799e-06, 
    1.429801e-06, 1.429799e-06, 1.429798e-06, 1.429794e-06, 1.42979e-06, 
    1.429786e-06, 1.429785e-06, 1.42978e-06, 1.429784e-06, 1.429777e-06, 
    1.429783e-06, 1.429773e-06, 1.42979e-06, 1.429783e-06, 1.429796e-06, 
    1.429795e-06, 1.429792e-06, 1.429786e-06, 1.429789e-06, 1.429786e-06, 
    1.429794e-06, 1.429799e-06, 1.4298e-06, 1.429802e-06, 1.4298e-06, 
    1.4298e-06, 1.429798e-06, 1.429798e-06, 1.429793e-06, 1.429796e-06, 
    1.429788e-06, 1.429786e-06, 1.429778e-06, 1.429773e-06, 1.429768e-06, 
    1.429766e-06, 1.429765e-06, 1.429765e-06 ;

 TOTPFTC =
  0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174 ;

 TOTPFTN =
  0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255 ;

 TOTPRODC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTPRODN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTSOMC =
  17.34462, 17.3446, 17.34461, 17.3446, 17.3446, 17.34459, 17.34462, 17.3446, 
    17.34461, 17.34462, 17.34457, 17.3446, 17.34455, 17.34457, 17.34453, 
    17.34455, 17.34453, 17.34453, 17.34452, 17.34452, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.3445, 17.34452, 17.34459, 17.34458, 17.34459, 
    17.34459, 17.34459, 17.3446, 17.34461, 17.34462, 17.34462, 17.34461, 
    17.34459, 17.3446, 17.34458, 17.34458, 17.34456, 17.34457, 17.34454, 
    17.34455, 17.34452, 17.34453, 17.34452, 17.34452, 17.34452, 17.34453, 
    17.34453, 17.34454, 17.34457, 17.34456, 17.34459, 17.3446, 17.34462, 
    17.34462, 17.34462, 17.34462, 17.34461, 17.3446, 17.34459, 17.34459, 
    17.34458, 17.34456, 17.34455, 17.34454, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34452, 17.34453, 17.34452, 17.34454, 17.34454, 
    17.34458, 17.34459, 17.3446, 17.34461, 17.34462, 17.34461, 17.34462, 
    17.34461, 17.3446, 17.3446, 17.34459, 17.34459, 17.34455, 17.34457, 
    17.34453, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34451, 17.34451, 17.34451, 17.34453, 17.34452, 17.3446, 17.3446, 
    17.3446, 17.34461, 17.34461, 17.34462, 17.34461, 17.34461, 17.3446, 
    17.34459, 17.34459, 17.34458, 17.34457, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34454, 17.34454, 17.34451, 17.34453, 17.34451, 
    17.34451, 17.34452, 17.34451, 17.3446, 17.3446, 17.34461, 17.34461, 
    17.34462, 17.34461, 17.34461, 17.34459, 17.34459, 17.34459, 17.34458, 
    17.34457, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 17.34453, 
    17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 17.34451, 17.34451, 
    17.34451, 17.3446, 17.3446, 17.3446, 17.3446, 17.3446, 17.34459, 
    17.34458, 17.34456, 17.34457, 17.34456, 17.34457, 17.34457, 17.34455, 
    17.34457, 17.34454, 17.34456, 17.34453, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34451, 17.3445, 17.3445, 17.34449, 17.34459, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34457, 17.34455, 17.34456, 
    17.34455, 17.34454, 17.34456, 17.34455, 17.34458, 17.34458, 17.34458, 
    17.34459, 17.34455, 17.34457, 17.34454, 17.34455, 17.34452, 17.34453, 
    17.34451, 17.34449, 17.34448, 17.34447, 17.34458, 17.34459, 17.34458, 
    17.34457, 17.34456, 17.34455, 17.34455, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34458, 17.34455, 17.34459, 17.34458, 17.34457, 
    17.34457, 17.34456, 17.34455, 17.34454, 17.34455, 17.3445, 17.34452, 
    17.34446, 17.34447, 17.34459, 17.34458, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34455, 17.34454, 17.34457, 17.34456, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34454, 17.34453, 17.34455, 17.34449, 17.34453, 
    17.34458, 17.34457, 17.34457, 17.34457, 17.34454, 17.34455, 17.34452, 
    17.34453, 17.34452, 17.34453, 17.34453, 17.34453, 17.34454, 17.34455, 
    17.34456, 17.34457, 17.34457, 17.34456, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34455, 17.34454, 17.34454, 17.34453, 17.34456, 17.34453, 
    17.34456, 17.34456, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 
    17.34454, 17.34455, 17.34455, 17.34455, 17.34456, 17.34456, 17.34456, 
    17.34456, 17.34454, 17.34453, 17.34452, 17.34451, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.34448, 17.34453, 17.34451, 17.34455, 17.34455, 
    17.34454, 17.34452, 17.34453, 17.34452, 17.34455, 17.34456, 17.34456, 
    17.34457, 17.34456, 17.34456, 17.34456, 17.34456, 17.34454, 17.34455, 
    17.34453, 17.34452, 17.34449, 17.34448, 17.34446, 17.34446, 17.34446, 
    17.34445 ;

 TOTSOMC_1m =
  17.34462, 17.3446, 17.34461, 17.3446, 17.3446, 17.34459, 17.34462, 17.3446, 
    17.34461, 17.34462, 17.34457, 17.3446, 17.34455, 17.34457, 17.34453, 
    17.34455, 17.34453, 17.34453, 17.34452, 17.34452, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.3445, 17.34452, 17.34459, 17.34458, 17.34459, 
    17.34459, 17.34459, 17.3446, 17.34461, 17.34462, 17.34462, 17.34461, 
    17.34459, 17.3446, 17.34458, 17.34458, 17.34456, 17.34457, 17.34454, 
    17.34455, 17.34452, 17.34453, 17.34452, 17.34452, 17.34452, 17.34453, 
    17.34453, 17.34454, 17.34457, 17.34456, 17.34459, 17.3446, 17.34462, 
    17.34462, 17.34462, 17.34462, 17.34461, 17.3446, 17.34459, 17.34459, 
    17.34458, 17.34456, 17.34455, 17.34454, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34452, 17.34453, 17.34452, 17.34454, 17.34454, 
    17.34458, 17.34459, 17.3446, 17.34461, 17.34462, 17.34461, 17.34462, 
    17.34461, 17.3446, 17.3446, 17.34459, 17.34459, 17.34455, 17.34457, 
    17.34453, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34451, 17.34451, 17.34451, 17.34453, 17.34452, 17.3446, 17.3446, 
    17.3446, 17.34461, 17.34461, 17.34462, 17.34461, 17.34461, 17.3446, 
    17.34459, 17.34459, 17.34458, 17.34457, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34454, 17.34454, 17.34451, 17.34453, 17.34451, 
    17.34451, 17.34452, 17.34451, 17.3446, 17.3446, 17.34461, 17.34461, 
    17.34462, 17.34461, 17.34461, 17.34459, 17.34459, 17.34459, 17.34458, 
    17.34457, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 17.34453, 
    17.34453, 17.34453, 17.34452, 17.34453, 17.34451, 17.34451, 17.34451, 
    17.34451, 17.3446, 17.3446, 17.3446, 17.3446, 17.3446, 17.34459, 
    17.34458, 17.34456, 17.34457, 17.34456, 17.34457, 17.34457, 17.34455, 
    17.34457, 17.34454, 17.34456, 17.34453, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34452, 17.34451, 17.3445, 17.3445, 17.34449, 17.34459, 
    17.34459, 17.34459, 17.34458, 17.34458, 17.34457, 17.34455, 17.34456, 
    17.34455, 17.34454, 17.34456, 17.34455, 17.34458, 17.34458, 17.34458, 
    17.34459, 17.34455, 17.34457, 17.34454, 17.34455, 17.34452, 17.34453, 
    17.34451, 17.34449, 17.34448, 17.34447, 17.34458, 17.34459, 17.34458, 
    17.34457, 17.34456, 17.34455, 17.34455, 17.34455, 17.34454, 17.34453, 
    17.34454, 17.34453, 17.34458, 17.34455, 17.34459, 17.34458, 17.34457, 
    17.34457, 17.34456, 17.34455, 17.34454, 17.34455, 17.3445, 17.34452, 
    17.34446, 17.34447, 17.34459, 17.34458, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34453, 17.34453, 17.34452, 17.34453, 17.34452, 
    17.34455, 17.34454, 17.34457, 17.34456, 17.34456, 17.34457, 17.34455, 
    17.34454, 17.34454, 17.34454, 17.34453, 17.34455, 17.34449, 17.34453, 
    17.34458, 17.34457, 17.34457, 17.34457, 17.34454, 17.34455, 17.34452, 
    17.34453, 17.34452, 17.34453, 17.34453, 17.34453, 17.34454, 17.34455, 
    17.34456, 17.34457, 17.34457, 17.34456, 17.34454, 17.34453, 17.34453, 
    17.34452, 17.34455, 17.34454, 17.34454, 17.34453, 17.34456, 17.34453, 
    17.34456, 17.34456, 17.34455, 17.34454, 17.34453, 17.34453, 17.34453, 
    17.34454, 17.34455, 17.34455, 17.34455, 17.34456, 17.34456, 17.34456, 
    17.34456, 17.34454, 17.34453, 17.34452, 17.34451, 17.3445, 17.34451, 
    17.34449, 17.34451, 17.34448, 17.34453, 17.34451, 17.34455, 17.34455, 
    17.34454, 17.34452, 17.34453, 17.34452, 17.34455, 17.34456, 17.34456, 
    17.34457, 17.34456, 17.34456, 17.34456, 17.34456, 17.34454, 17.34455, 
    17.34453, 17.34452, 17.34449, 17.34448, 17.34446, 17.34446, 17.34446, 
    17.34445 ;

 TOTSOMN =
  1.773759, 1.773758, 1.773758, 1.773756, 1.773757, 1.773756, 1.773759, 
    1.773757, 1.773759, 1.773759, 1.773753, 1.773756, 1.77375, 1.773752, 
    1.773747, 1.773751, 1.773747, 1.773747, 1.773745, 1.773746, 1.773743, 
    1.773745, 1.773742, 1.773744, 1.773743, 1.773745, 1.773756, 1.773754, 
    1.773756, 1.773756, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773758, 1.773755, 1.773756, 1.773754, 1.773754, 1.773751, 1.773753, 
    1.773748, 1.773749, 1.773746, 1.773747, 1.773746, 1.773746, 1.773746, 
    1.773747, 1.773747, 1.773748, 1.773752, 1.773751, 1.773755, 1.773757, 
    1.773759, 1.77376, 1.77376, 1.77376, 1.773758, 1.773757, 1.773756, 
    1.773755, 1.773754, 1.773752, 1.773751, 1.773748, 1.773749, 1.773748, 
    1.773747, 1.773746, 1.773746, 1.773745, 1.773748, 1.773746, 1.773749, 
    1.773748, 1.773754, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773759, 1.773758, 1.773757, 1.773757, 1.773755, 1.773756, 1.773751, 
    1.773753, 1.773747, 1.773748, 1.773747, 1.773748, 1.773746, 1.773747, 
    1.773745, 1.773744, 1.773745, 1.773744, 1.773747, 1.773746, 1.773757, 
    1.773757, 1.773757, 1.773758, 1.773758, 1.77376, 1.773759, 1.773758, 
    1.773757, 1.773756, 1.773755, 1.773754, 1.773752, 1.77375, 1.773748, 
    1.773747, 1.773748, 1.773747, 1.773748, 1.773748, 1.773745, 1.773747, 
    1.773744, 1.773744, 1.773745, 1.773744, 1.773757, 1.773758, 1.773759, 
    1.773758, 1.77376, 1.773759, 1.773758, 1.773756, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.77375, 1.773749, 1.773747, 1.773747, 1.773747, 
    1.773747, 1.773747, 1.773746, 1.773746, 1.773747, 1.773744, 1.773745, 
    1.773744, 1.773744, 1.773757, 1.773757, 1.773757, 1.773757, 1.773757, 
    1.773755, 1.773754, 1.773751, 1.773753, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773752, 1.773749, 1.773751, 1.773746, 1.773749, 1.773746, 
    1.773747, 1.773746, 1.773745, 1.773744, 1.773743, 1.773743, 1.773742, 
    1.773756, 1.773755, 1.773755, 1.773754, 1.773754, 1.773752, 1.77375, 
    1.773751, 1.773749, 1.773749, 1.773751, 1.77375, 1.773754, 1.773754, 
    1.773754, 1.773756, 1.773751, 1.773753, 1.773748, 1.77375, 1.773745, 
    1.773748, 1.773743, 1.773742, 1.77374, 1.773738, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.773751, 1.77375, 1.773749, 1.773749, 1.773748, 
    1.773748, 1.773749, 1.773747, 1.773754, 1.77375, 1.773755, 1.773754, 
    1.773753, 1.773753, 1.773751, 1.77375, 1.773748, 1.773749, 1.773742, 
    1.773745, 1.773736, 1.773739, 1.773755, 1.773755, 1.773752, 1.773753, 
    1.773749, 1.773749, 1.773748, 1.773747, 1.773747, 1.773746, 1.773747, 
    1.773746, 1.77375, 1.773748, 1.773752, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773749, 1.773749, 1.773748, 1.773747, 1.773749, 1.773742, 
    1.773746, 1.773754, 1.773752, 1.773752, 1.773753, 1.773749, 1.77375, 
    1.773746, 1.773747, 1.773746, 1.773746, 1.773747, 1.773748, 1.773748, 
    1.77375, 1.773751, 1.773753, 1.773752, 1.773751, 1.773749, 1.773747, 
    1.773747, 1.773746, 1.77375, 1.773748, 1.773749, 1.773747, 1.773751, 
    1.773748, 1.773752, 1.773751, 1.77375, 1.773748, 1.773748, 1.773747, 
    1.773747, 1.773749, 1.773749, 1.77375, 1.77375, 1.773751, 1.773752, 
    1.773751, 1.773751, 1.773749, 1.773747, 1.773745, 1.773745, 1.773743, 
    1.773744, 1.773742, 1.773744, 1.77374, 1.773747, 1.773744, 1.77375, 
    1.773749, 1.773748, 1.773746, 1.773747, 1.773745, 1.773749, 1.773751, 
    1.773751, 1.773752, 1.773751, 1.773752, 1.773751, 1.773751, 1.773749, 
    1.77375, 1.773747, 1.773745, 1.773742, 1.77374, 1.773738, 1.773737, 
    1.773736, 1.773736 ;

 TOTSOMN_1m =
  1.773759, 1.773758, 1.773758, 1.773756, 1.773757, 1.773756, 1.773759, 
    1.773757, 1.773759, 1.773759, 1.773753, 1.773756, 1.77375, 1.773752, 
    1.773747, 1.773751, 1.773747, 1.773747, 1.773745, 1.773746, 1.773743, 
    1.773745, 1.773742, 1.773744, 1.773743, 1.773745, 1.773756, 1.773754, 
    1.773756, 1.773756, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773758, 1.773755, 1.773756, 1.773754, 1.773754, 1.773751, 1.773753, 
    1.773748, 1.773749, 1.773746, 1.773747, 1.773746, 1.773746, 1.773746, 
    1.773747, 1.773747, 1.773748, 1.773752, 1.773751, 1.773755, 1.773757, 
    1.773759, 1.77376, 1.77376, 1.77376, 1.773758, 1.773757, 1.773756, 
    1.773755, 1.773754, 1.773752, 1.773751, 1.773748, 1.773749, 1.773748, 
    1.773747, 1.773746, 1.773746, 1.773745, 1.773748, 1.773746, 1.773749, 
    1.773748, 1.773754, 1.773756, 1.773757, 1.773758, 1.77376, 1.773759, 
    1.773759, 1.773758, 1.773757, 1.773757, 1.773755, 1.773756, 1.773751, 
    1.773753, 1.773747, 1.773748, 1.773747, 1.773748, 1.773746, 1.773747, 
    1.773745, 1.773744, 1.773745, 1.773744, 1.773747, 1.773746, 1.773757, 
    1.773757, 1.773757, 1.773758, 1.773758, 1.77376, 1.773759, 1.773758, 
    1.773757, 1.773756, 1.773755, 1.773754, 1.773752, 1.77375, 1.773748, 
    1.773747, 1.773748, 1.773747, 1.773748, 1.773748, 1.773745, 1.773747, 
    1.773744, 1.773744, 1.773745, 1.773744, 1.773757, 1.773758, 1.773759, 
    1.773758, 1.77376, 1.773759, 1.773758, 1.773756, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.77375, 1.773749, 1.773747, 1.773747, 1.773747, 
    1.773747, 1.773747, 1.773746, 1.773746, 1.773747, 1.773744, 1.773745, 
    1.773744, 1.773744, 1.773757, 1.773757, 1.773757, 1.773757, 1.773757, 
    1.773755, 1.773754, 1.773751, 1.773753, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773752, 1.773749, 1.773751, 1.773746, 1.773749, 1.773746, 
    1.773747, 1.773746, 1.773745, 1.773744, 1.773743, 1.773743, 1.773742, 
    1.773756, 1.773755, 1.773755, 1.773754, 1.773754, 1.773752, 1.77375, 
    1.773751, 1.773749, 1.773749, 1.773751, 1.77375, 1.773754, 1.773754, 
    1.773754, 1.773756, 1.773751, 1.773753, 1.773748, 1.77375, 1.773745, 
    1.773748, 1.773743, 1.773742, 1.77374, 1.773738, 1.773755, 1.773755, 
    1.773754, 1.773753, 1.773751, 1.77375, 1.773749, 1.773749, 1.773748, 
    1.773748, 1.773749, 1.773747, 1.773754, 1.77375, 1.773755, 1.773754, 
    1.773753, 1.773753, 1.773751, 1.77375, 1.773748, 1.773749, 1.773742, 
    1.773745, 1.773736, 1.773739, 1.773755, 1.773755, 1.773752, 1.773753, 
    1.773749, 1.773749, 1.773748, 1.773747, 1.773747, 1.773746, 1.773747, 
    1.773746, 1.77375, 1.773748, 1.773752, 1.773751, 1.773752, 1.773752, 
    1.773751, 1.773749, 1.773749, 1.773748, 1.773747, 1.773749, 1.773742, 
    1.773746, 1.773754, 1.773752, 1.773752, 1.773753, 1.773749, 1.77375, 
    1.773746, 1.773747, 1.773746, 1.773746, 1.773747, 1.773748, 1.773748, 
    1.77375, 1.773751, 1.773753, 1.773752, 1.773751, 1.773749, 1.773747, 
    1.773747, 1.773746, 1.77375, 1.773748, 1.773749, 1.773747, 1.773751, 
    1.773748, 1.773752, 1.773751, 1.77375, 1.773748, 1.773748, 1.773747, 
    1.773747, 1.773749, 1.773749, 1.77375, 1.77375, 1.773751, 1.773752, 
    1.773751, 1.773751, 1.773749, 1.773747, 1.773745, 1.773745, 1.773743, 
    1.773744, 1.773742, 1.773744, 1.77374, 1.773747, 1.773744, 1.77375, 
    1.773749, 1.773748, 1.773746, 1.773747, 1.773745, 1.773749, 1.773751, 
    1.773751, 1.773752, 1.773751, 1.773752, 1.773751, 1.773751, 1.773749, 
    1.77375, 1.773747, 1.773745, 1.773742, 1.77374, 1.773738, 1.773737, 
    1.773736, 1.773736 ;

 TOTVEGC =
  0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 0.8953174, 
    0.8953174, 0.8953174 ;

 TOTVEGN =
  0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 0.03250255, 
    0.03250255, 0.03250255 ;

 TREFMNAV =
  243.0864, 243.0896, 243.089, 243.0916, 243.0902, 243.0918, 243.0871, 
    243.0897, 243.088, 243.0867, 243.0965, 243.0917, 243.1017, 243.0986, 
    243.1064, 243.1012, 243.1074, 243.1063, 243.1098, 243.1088, 243.1133, 
    243.1103, 243.1157, 243.1126, 243.1131, 243.1102, 243.0927, 243.0959, 
    243.0925, 243.093, 243.0928, 243.0902, 243.0888, 243.0862, 243.0867, 
    243.0886, 243.0932, 243.0917, 243.0956, 243.0955, 243.0997, 243.0978, 
    243.105, 243.103, 243.1089, 243.1074, 243.1088, 243.1084, 243.1088, 
    243.1066, 243.1076, 243.1057, 243.0982, 243.1004, 243.0938, 243.0897, 
    243.0872, 243.0853, 243.0856, 243.086, 243.0887, 243.0911, 243.093, 
    243.0942, 243.0955, 243.099, 243.101, 243.1054, 243.1047, 243.1059, 
    243.1072, 243.1094, 243.109, 243.1099, 243.1059, 243.1086, 243.1042, 
    243.1054, 243.0956, 243.0921, 243.0904, 243.0891, 243.0858, 243.0881, 
    243.0872, 243.0894, 243.0907, 243.0901, 243.0943, 243.0926, 243.1012, 
    243.0975, 243.1071, 243.1048, 243.1077, 243.1062, 243.1087, 243.1065, 
    243.1103, 243.1111, 243.1105, 243.1127, 243.1063, 243.1088, 243.09, 
    243.0901, 243.0907, 243.0883, 243.0882, 243.0861, 243.088, 243.0888, 
    243.0908, 243.092, 243.0931, 243.0956, 243.0983, 243.1022, 243.105, 
    243.1068, 243.1057, 243.1067, 243.1056, 243.1051, 243.1108, 243.1076, 
    243.1124, 243.1122, 243.1099, 243.1122, 243.0902, 243.0896, 243.0873, 
    243.0891, 243.0859, 243.0877, 243.0887, 243.0926, 243.0935, 243.0943, 
    243.0959, 243.0979, 243.1014, 243.1045, 243.1073, 243.1071, 243.1072, 
    243.1078, 243.1063, 243.1081, 243.1083, 243.1076, 243.1121, 243.1108, 
    243.1122, 243.1113, 243.0898, 243.0909, 243.0903, 243.0914, 243.0906, 
    243.094, 243.095, 243.0998, 243.0979, 243.101, 243.0982, 243.0987, 
    243.101, 243.0984, 243.1043, 243.1002, 243.1078, 243.1037, 243.1081, 
    243.1073, 243.1086, 243.1097, 243.1112, 243.1138, 243.1132, 243.1154, 
    243.0925, 243.0939, 243.0938, 243.0952, 243.0963, 243.0986, 243.1023, 
    243.101, 243.1035, 243.104, 243.1001, 243.1025, 243.0948, 243.096, 
    243.0953, 243.0926, 243.1012, 243.0968, 243.105, 243.1026, 243.1096, 
    243.1061, 243.1129, 243.1157, 243.1185, 243.1215, 243.0946, 243.0937, 
    243.0954, 243.0977, 243.0999, 243.1028, 243.1031, 243.1036, 243.105, 
    243.1062, 243.1037, 243.1064, 243.0962, 243.1016, 243.0933, 243.0958, 
    243.0976, 243.0968, 243.1008, 243.1017, 243.1055, 243.1035, 243.115, 
    243.1099, 243.124, 243.1201, 243.0934, 243.0947, 243.099, 243.097, 
    243.103, 243.1044, 243.1056, 243.1071, 243.1073, 243.1082, 243.1067, 
    243.1082, 243.1028, 243.1052, 243.0986, 243.1002, 243.0994, 243.0986, 
    243.1011, 243.1037, 243.1039, 243.1047, 243.1069, 243.103, 243.1155, 
    243.1077, 243.096, 243.0984, 243.0988, 243.0979, 243.1043, 243.102, 
    243.1082, 243.1065, 243.1093, 243.1079, 243.1077, 243.1059, 243.1048, 
    243.1021, 243.0998, 243.098, 243.0984, 243.1004, 243.1039, 243.1073, 
    243.1066, 243.1091, 243.1025, 243.1052, 243.1042, 243.107, 243.1009, 
    243.1059, 243.0996, 243.1002, 243.1019, 243.1054, 243.1062, 243.107, 
    243.1066, 243.104, 243.1036, 243.1019, 243.1014, 243.1001, 243.0989, 
    243.0999, 243.101, 243.104, 243.1068, 243.1097, 243.1105, 243.1138, 
    243.111, 243.1155, 243.1116, 243.1185, 243.1063, 243.1116, 243.102, 
    243.1031, 243.1049, 243.1092, 243.1069, 243.1096, 243.1036, 243.1004, 
    243.0997, 243.0981, 243.0997, 243.0996, 243.1011, 243.1006, 243.1042, 
    243.1022, 243.1077, 243.1096, 243.1152, 243.1185, 243.1221, 243.1236, 
    243.124, 243.1242 ;

 TREFMNAV_R =
  243.0864, 243.0896, 243.089, 243.0916, 243.0902, 243.0918, 243.0871, 
    243.0897, 243.088, 243.0867, 243.0965, 243.0917, 243.1017, 243.0986, 
    243.1064, 243.1012, 243.1074, 243.1063, 243.1098, 243.1088, 243.1133, 
    243.1103, 243.1157, 243.1126, 243.1131, 243.1102, 243.0927, 243.0959, 
    243.0925, 243.093, 243.0928, 243.0902, 243.0888, 243.0862, 243.0867, 
    243.0886, 243.0932, 243.0917, 243.0956, 243.0955, 243.0997, 243.0978, 
    243.105, 243.103, 243.1089, 243.1074, 243.1088, 243.1084, 243.1088, 
    243.1066, 243.1076, 243.1057, 243.0982, 243.1004, 243.0938, 243.0897, 
    243.0872, 243.0853, 243.0856, 243.086, 243.0887, 243.0911, 243.093, 
    243.0942, 243.0955, 243.099, 243.101, 243.1054, 243.1047, 243.1059, 
    243.1072, 243.1094, 243.109, 243.1099, 243.1059, 243.1086, 243.1042, 
    243.1054, 243.0956, 243.0921, 243.0904, 243.0891, 243.0858, 243.0881, 
    243.0872, 243.0894, 243.0907, 243.0901, 243.0943, 243.0926, 243.1012, 
    243.0975, 243.1071, 243.1048, 243.1077, 243.1062, 243.1087, 243.1065, 
    243.1103, 243.1111, 243.1105, 243.1127, 243.1063, 243.1088, 243.09, 
    243.0901, 243.0907, 243.0883, 243.0882, 243.0861, 243.088, 243.0888, 
    243.0908, 243.092, 243.0931, 243.0956, 243.0983, 243.1022, 243.105, 
    243.1068, 243.1057, 243.1067, 243.1056, 243.1051, 243.1108, 243.1076, 
    243.1124, 243.1122, 243.1099, 243.1122, 243.0902, 243.0896, 243.0873, 
    243.0891, 243.0859, 243.0877, 243.0887, 243.0926, 243.0935, 243.0943, 
    243.0959, 243.0979, 243.1014, 243.1045, 243.1073, 243.1071, 243.1072, 
    243.1078, 243.1063, 243.1081, 243.1083, 243.1076, 243.1121, 243.1108, 
    243.1122, 243.1113, 243.0898, 243.0909, 243.0903, 243.0914, 243.0906, 
    243.094, 243.095, 243.0998, 243.0979, 243.101, 243.0982, 243.0987, 
    243.101, 243.0984, 243.1043, 243.1002, 243.1078, 243.1037, 243.1081, 
    243.1073, 243.1086, 243.1097, 243.1112, 243.1138, 243.1132, 243.1154, 
    243.0925, 243.0939, 243.0938, 243.0952, 243.0963, 243.0986, 243.1023, 
    243.101, 243.1035, 243.104, 243.1001, 243.1025, 243.0948, 243.096, 
    243.0953, 243.0926, 243.1012, 243.0968, 243.105, 243.1026, 243.1096, 
    243.1061, 243.1129, 243.1157, 243.1185, 243.1215, 243.0946, 243.0937, 
    243.0954, 243.0977, 243.0999, 243.1028, 243.1031, 243.1036, 243.105, 
    243.1062, 243.1037, 243.1064, 243.0962, 243.1016, 243.0933, 243.0958, 
    243.0976, 243.0968, 243.1008, 243.1017, 243.1055, 243.1035, 243.115, 
    243.1099, 243.124, 243.1201, 243.0934, 243.0947, 243.099, 243.097, 
    243.103, 243.1044, 243.1056, 243.1071, 243.1073, 243.1082, 243.1067, 
    243.1082, 243.1028, 243.1052, 243.0986, 243.1002, 243.0994, 243.0986, 
    243.1011, 243.1037, 243.1039, 243.1047, 243.1069, 243.103, 243.1155, 
    243.1077, 243.096, 243.0984, 243.0988, 243.0979, 243.1043, 243.102, 
    243.1082, 243.1065, 243.1093, 243.1079, 243.1077, 243.1059, 243.1048, 
    243.1021, 243.0998, 243.098, 243.0984, 243.1004, 243.1039, 243.1073, 
    243.1066, 243.1091, 243.1025, 243.1052, 243.1042, 243.107, 243.1009, 
    243.1059, 243.0996, 243.1002, 243.1019, 243.1054, 243.1062, 243.107, 
    243.1066, 243.104, 243.1036, 243.1019, 243.1014, 243.1001, 243.0989, 
    243.0999, 243.101, 243.104, 243.1068, 243.1097, 243.1105, 243.1138, 
    243.111, 243.1155, 243.1116, 243.1185, 243.1063, 243.1116, 243.102, 
    243.1031, 243.1049, 243.1092, 243.1069, 243.1096, 243.1036, 243.1004, 
    243.0997, 243.0981, 243.0997, 243.0996, 243.1011, 243.1006, 243.1042, 
    243.1022, 243.1077, 243.1096, 243.1152, 243.1185, 243.1221, 243.1236, 
    243.124, 243.1242 ;

 TREFMNAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TREFMXAV =
  270.7704, 270.7683, 270.7687, 270.767, 270.7679, 270.7668, 270.77, 
    270.7682, 270.7693, 270.7702, 270.7638, 270.7669, 270.7603, 270.7624, 
    270.7572, 270.7607, 270.7565, 270.7573, 270.7549, 270.7556, 270.7526, 
    270.7545, 270.7509, 270.753, 270.7527, 270.7546, 270.7663, 270.7642, 
    270.7664, 270.7661, 270.7662, 270.7679, 270.7688, 270.7706, 270.7702, 
    270.769, 270.766, 270.7669, 270.7644, 270.7644, 270.7616, 270.7629, 
    270.7581, 270.7595, 270.7555, 270.7565, 270.7556, 270.7559, 270.7556, 
    270.757, 270.7564, 270.7577, 270.7627, 270.7612, 270.7656, 270.7682, 
    270.7699, 270.7711, 270.771, 270.7706, 270.769, 270.7673, 270.7661, 
    270.7653, 270.7645, 270.7621, 270.7608, 270.7579, 270.7584, 270.7575, 
    270.7566, 270.7552, 270.7554, 270.7548, 270.7575, 270.7557, 270.7586, 
    270.7578, 270.7644, 270.7667, 270.7678, 270.7686, 270.7708, 270.7693, 
    270.7699, 270.7685, 270.7676, 270.768, 270.7652, 270.7663, 270.7607, 
    270.7631, 270.7567, 270.7582, 270.7563, 270.7573, 270.7557, 270.7571, 
    270.7546, 270.754, 270.7544, 270.7529, 270.7572, 270.7556, 270.768, 
    270.7679, 270.7676, 270.7691, 270.7692, 270.7706, 270.7693, 270.7689, 
    270.7675, 270.7667, 270.766, 270.7644, 270.7626, 270.76, 270.7581, 
    270.7569, 270.7577, 270.757, 270.7578, 270.7581, 270.7542, 270.7564, 
    270.7531, 270.7533, 270.7548, 270.7533, 270.7679, 270.7683, 270.7698, 
    270.7686, 270.7707, 270.7696, 270.7689, 270.7663, 270.7657, 270.7652, 
    270.7642, 270.7628, 270.7605, 270.7585, 270.7566, 270.7567, 270.7567, 
    270.7563, 270.7573, 270.7561, 270.7559, 270.7564, 270.7534, 270.7542, 
    270.7533, 270.7539, 270.7682, 270.7675, 270.7679, 270.7672, 270.7677, 
    270.7654, 270.7648, 270.7616, 270.7628, 270.7608, 270.7626, 270.7623, 
    270.7608, 270.7625, 270.7586, 270.7613, 270.7562, 270.759, 270.7561, 
    270.7566, 270.7557, 270.7549, 270.754, 270.7522, 270.7526, 270.7511, 
    270.7664, 270.7655, 270.7656, 270.7646, 270.7639, 270.7624, 270.7599, 
    270.7608, 270.7591, 270.7588, 270.7614, 270.7598, 270.7649, 270.7641, 
    270.7646, 270.7664, 270.7607, 270.7636, 270.7581, 270.7597, 270.7551, 
    270.7574, 270.7528, 270.7509, 270.7491, 270.747, 270.765, 270.7656, 
    270.7645, 270.763, 270.7615, 270.7596, 270.7594, 270.7591, 270.7581, 
    270.7574, 270.759, 270.7571, 270.764, 270.7604, 270.7659, 270.7643, 
    270.7631, 270.7636, 270.7609, 270.7603, 270.7578, 270.7591, 270.7514, 
    270.7548, 270.7453, 270.748, 270.7658, 270.765, 270.7621, 270.7635, 
    270.7595, 270.7585, 270.7577, 270.7567, 270.7566, 270.756, 270.757, 
    270.756, 270.7596, 270.758, 270.7624, 270.7614, 270.7618, 270.7624, 
    270.7607, 270.759, 270.7589, 270.7583, 270.7569, 270.7595, 270.7511, 
    270.7563, 270.7641, 270.7625, 270.7622, 270.7628, 270.7586, 270.7602, 
    270.756, 270.7571, 270.7553, 270.7562, 270.7563, 270.7575, 270.7582, 
    270.7601, 270.7616, 270.7628, 270.7625, 270.7612, 270.7589, 270.7566, 
    270.7571, 270.7554, 270.7598, 270.758, 270.7587, 270.7568, 270.7609, 
    270.7575, 270.7617, 270.7614, 270.7602, 270.7579, 270.7573, 270.7568, 
    270.7571, 270.7588, 270.759, 270.7602, 270.7606, 270.7614, 270.7622, 
    270.7615, 270.7608, 270.7588, 270.7569, 270.7549, 270.7545, 270.7522, 
    270.7541, 270.7511, 270.7537, 270.7491, 270.7573, 270.7537, 270.7601, 
    270.7594, 270.7582, 270.7553, 270.7568, 270.755, 270.759, 270.7612, 
    270.7617, 270.7627, 270.7617, 270.7617, 270.7607, 270.761, 270.7587, 
    270.7599, 270.7563, 270.755, 270.7513, 270.749, 270.7466, 270.7456, 
    270.7453, 270.7451 ;

 TREFMXAV_R =
  270.7704, 270.7683, 270.7687, 270.767, 270.7679, 270.7668, 270.77, 
    270.7682, 270.7693, 270.7702, 270.7638, 270.7669, 270.7603, 270.7624, 
    270.7572, 270.7607, 270.7565, 270.7573, 270.7549, 270.7556, 270.7526, 
    270.7545, 270.7509, 270.753, 270.7527, 270.7546, 270.7663, 270.7642, 
    270.7664, 270.7661, 270.7662, 270.7679, 270.7688, 270.7706, 270.7702, 
    270.769, 270.766, 270.7669, 270.7644, 270.7644, 270.7616, 270.7629, 
    270.7581, 270.7595, 270.7555, 270.7565, 270.7556, 270.7559, 270.7556, 
    270.757, 270.7564, 270.7577, 270.7627, 270.7612, 270.7656, 270.7682, 
    270.7699, 270.7711, 270.771, 270.7706, 270.769, 270.7673, 270.7661, 
    270.7653, 270.7645, 270.7621, 270.7608, 270.7579, 270.7584, 270.7575, 
    270.7566, 270.7552, 270.7554, 270.7548, 270.7575, 270.7557, 270.7586, 
    270.7578, 270.7644, 270.7667, 270.7678, 270.7686, 270.7708, 270.7693, 
    270.7699, 270.7685, 270.7676, 270.768, 270.7652, 270.7663, 270.7607, 
    270.7631, 270.7567, 270.7582, 270.7563, 270.7573, 270.7557, 270.7571, 
    270.7546, 270.754, 270.7544, 270.7529, 270.7572, 270.7556, 270.768, 
    270.7679, 270.7676, 270.7691, 270.7692, 270.7706, 270.7693, 270.7689, 
    270.7675, 270.7667, 270.766, 270.7644, 270.7626, 270.76, 270.7581, 
    270.7569, 270.7577, 270.757, 270.7578, 270.7581, 270.7542, 270.7564, 
    270.7531, 270.7533, 270.7548, 270.7533, 270.7679, 270.7683, 270.7698, 
    270.7686, 270.7707, 270.7696, 270.7689, 270.7663, 270.7657, 270.7652, 
    270.7642, 270.7628, 270.7605, 270.7585, 270.7566, 270.7567, 270.7567, 
    270.7563, 270.7573, 270.7561, 270.7559, 270.7564, 270.7534, 270.7542, 
    270.7533, 270.7539, 270.7682, 270.7675, 270.7679, 270.7672, 270.7677, 
    270.7654, 270.7648, 270.7616, 270.7628, 270.7608, 270.7626, 270.7623, 
    270.7608, 270.7625, 270.7586, 270.7613, 270.7562, 270.759, 270.7561, 
    270.7566, 270.7557, 270.7549, 270.754, 270.7522, 270.7526, 270.7511, 
    270.7664, 270.7655, 270.7656, 270.7646, 270.7639, 270.7624, 270.7599, 
    270.7608, 270.7591, 270.7588, 270.7614, 270.7598, 270.7649, 270.7641, 
    270.7646, 270.7664, 270.7607, 270.7636, 270.7581, 270.7597, 270.7551, 
    270.7574, 270.7528, 270.7509, 270.7491, 270.747, 270.765, 270.7656, 
    270.7645, 270.763, 270.7615, 270.7596, 270.7594, 270.7591, 270.7581, 
    270.7574, 270.759, 270.7571, 270.764, 270.7604, 270.7659, 270.7643, 
    270.7631, 270.7636, 270.7609, 270.7603, 270.7578, 270.7591, 270.7514, 
    270.7548, 270.7453, 270.748, 270.7658, 270.765, 270.7621, 270.7635, 
    270.7595, 270.7585, 270.7577, 270.7567, 270.7566, 270.756, 270.757, 
    270.756, 270.7596, 270.758, 270.7624, 270.7614, 270.7618, 270.7624, 
    270.7607, 270.759, 270.7589, 270.7583, 270.7569, 270.7595, 270.7511, 
    270.7563, 270.7641, 270.7625, 270.7622, 270.7628, 270.7586, 270.7602, 
    270.756, 270.7571, 270.7553, 270.7562, 270.7563, 270.7575, 270.7582, 
    270.7601, 270.7616, 270.7628, 270.7625, 270.7612, 270.7589, 270.7566, 
    270.7571, 270.7554, 270.7598, 270.758, 270.7587, 270.7568, 270.7609, 
    270.7575, 270.7617, 270.7614, 270.7602, 270.7579, 270.7573, 270.7568, 
    270.7571, 270.7588, 270.759, 270.7602, 270.7606, 270.7614, 270.7622, 
    270.7615, 270.7608, 270.7588, 270.7569, 270.7549, 270.7545, 270.7522, 
    270.7541, 270.7511, 270.7537, 270.7491, 270.7573, 270.7537, 270.7601, 
    270.7594, 270.7582, 270.7553, 270.7568, 270.755, 270.759, 270.7612, 
    270.7617, 270.7627, 270.7617, 270.7617, 270.7607, 270.761, 270.7587, 
    270.7599, 270.7563, 270.755, 270.7513, 270.749, 270.7466, 270.7456, 
    270.7453, 270.7451 ;

 TREFMXAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSA =
  255.2069, 255.2067, 255.2068, 255.2066, 255.2067, 255.2066, 255.2069, 
    255.2067, 255.2068, 255.2069, 255.2064, 255.2066, 255.2061, 255.2063, 
    255.2059, 255.2061, 255.2058, 255.2059, 255.2057, 255.2057, 255.2055, 
    255.2056, 255.2054, 255.2055, 255.2055, 255.2056, 255.2066, 255.2064, 
    255.2066, 255.2066, 255.2066, 255.2067, 255.2068, 255.2069, 255.2069, 
    255.2068, 255.2066, 255.2066, 255.2064, 255.2064, 255.2062, 255.2063, 
    255.2059, 255.206, 255.2057, 255.2058, 255.2057, 255.2057, 255.2057, 
    255.2058, 255.2058, 255.2059, 255.2063, 255.2062, 255.2065, 255.2067, 
    255.2069, 255.207, 255.2069, 255.2069, 255.2068, 255.2067, 255.2066, 
    255.2065, 255.2064, 255.2063, 255.2061, 255.2059, 255.2059, 255.2059, 
    255.2058, 255.2057, 255.2057, 255.2057, 255.2059, 255.2057, 255.206, 
    255.2059, 255.2064, 255.2066, 255.2067, 255.2068, 255.2069, 255.2068, 
    255.2069, 255.2067, 255.2067, 255.2067, 255.2065, 255.2066, 255.2061, 
    255.2063, 255.2058, 255.2059, 255.2058, 255.2059, 255.2057, 255.2059, 
    255.2056, 255.2056, 255.2056, 255.2055, 255.2059, 255.2057, 255.2067, 
    255.2067, 255.2067, 255.2068, 255.2068, 255.2069, 255.2068, 255.2068, 
    255.2067, 255.2066, 255.2066, 255.2064, 255.2063, 255.2061, 255.2059, 
    255.2058, 255.2059, 255.2058, 255.2059, 255.2059, 255.2056, 255.2058, 
    255.2055, 255.2055, 255.2057, 255.2055, 255.2067, 255.2067, 255.2068, 
    255.2068, 255.2069, 255.2068, 255.2068, 255.2066, 255.2065, 255.2065, 
    255.2064, 255.2063, 255.2061, 255.206, 255.2058, 255.2058, 255.2058, 
    255.2058, 255.2059, 255.2058, 255.2057, 255.2058, 255.2056, 255.2056, 
    255.2055, 255.2056, 255.2067, 255.2067, 255.2067, 255.2066, 255.2067, 
    255.2065, 255.2065, 255.2062, 255.2063, 255.2061, 255.2063, 255.2063, 
    255.2061, 255.2063, 255.206, 255.2062, 255.2058, 255.206, 255.2058, 
    255.2058, 255.2057, 255.2057, 255.2056, 255.2055, 255.2055, 255.2054, 
    255.2066, 255.2065, 255.2065, 255.2065, 255.2064, 255.2063, 255.2061, 
    255.2061, 255.206, 255.206, 255.2062, 255.2061, 255.2065, 255.2064, 
    255.2065, 255.2066, 255.2061, 255.2064, 255.2059, 255.2061, 255.2057, 
    255.2059, 255.2055, 255.2054, 255.2052, 255.205, 255.2065, 255.2065, 
    255.2064, 255.2063, 255.2062, 255.2061, 255.206, 255.206, 255.2059, 
    255.2059, 255.206, 255.2059, 255.2064, 255.2061, 255.2065, 255.2064, 
    255.2063, 255.2064, 255.2062, 255.2061, 255.2059, 255.206, 255.2054, 
    255.2057, 255.2049, 255.2051, 255.2065, 255.2065, 255.2063, 255.2064, 
    255.206, 255.206, 255.2059, 255.2058, 255.2058, 255.2058, 255.2058, 
    255.2058, 255.2061, 255.2059, 255.2063, 255.2062, 255.2062, 255.2063, 
    255.2061, 255.206, 255.206, 255.2059, 255.2058, 255.206, 255.2054, 
    255.2058, 255.2064, 255.2063, 255.2063, 255.2063, 255.206, 255.2061, 
    255.2058, 255.2059, 255.2057, 255.2058, 255.2058, 255.2059, 255.2059, 
    255.2061, 255.2062, 255.2063, 255.2063, 255.2062, 255.206, 255.2058, 
    255.2058, 255.2057, 255.2061, 255.2059, 255.206, 255.2058, 255.2061, 
    255.2059, 255.2062, 255.2062, 255.2061, 255.2059, 255.2059, 255.2058, 
    255.2058, 255.206, 255.206, 255.2061, 255.2061, 255.2062, 255.2063, 
    255.2062, 255.2061, 255.206, 255.2058, 255.2057, 255.2056, 255.2055, 
    255.2056, 255.2054, 255.2056, 255.2052, 255.2059, 255.2056, 255.2061, 
    255.206, 255.2059, 255.2057, 255.2058, 255.2057, 255.206, 255.2062, 
    255.2062, 255.2063, 255.2062, 255.2062, 255.2061, 255.2062, 255.206, 
    255.2061, 255.2058, 255.2057, 255.2054, 255.2052, 255.205, 255.2049, 
    255.2049, 255.2049 ;

 TSAI =
  0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 0.4323173, 
    0.4323173, 0.4323173 ;

 TSA_R =
  255.2069, 255.2067, 255.2068, 255.2066, 255.2067, 255.2066, 255.2069, 
    255.2067, 255.2068, 255.2069, 255.2064, 255.2066, 255.2061, 255.2063, 
    255.2059, 255.2061, 255.2058, 255.2059, 255.2057, 255.2057, 255.2055, 
    255.2056, 255.2054, 255.2055, 255.2055, 255.2056, 255.2066, 255.2064, 
    255.2066, 255.2066, 255.2066, 255.2067, 255.2068, 255.2069, 255.2069, 
    255.2068, 255.2066, 255.2066, 255.2064, 255.2064, 255.2062, 255.2063, 
    255.2059, 255.206, 255.2057, 255.2058, 255.2057, 255.2057, 255.2057, 
    255.2058, 255.2058, 255.2059, 255.2063, 255.2062, 255.2065, 255.2067, 
    255.2069, 255.207, 255.2069, 255.2069, 255.2068, 255.2067, 255.2066, 
    255.2065, 255.2064, 255.2063, 255.2061, 255.2059, 255.2059, 255.2059, 
    255.2058, 255.2057, 255.2057, 255.2057, 255.2059, 255.2057, 255.206, 
    255.2059, 255.2064, 255.2066, 255.2067, 255.2068, 255.2069, 255.2068, 
    255.2069, 255.2067, 255.2067, 255.2067, 255.2065, 255.2066, 255.2061, 
    255.2063, 255.2058, 255.2059, 255.2058, 255.2059, 255.2057, 255.2059, 
    255.2056, 255.2056, 255.2056, 255.2055, 255.2059, 255.2057, 255.2067, 
    255.2067, 255.2067, 255.2068, 255.2068, 255.2069, 255.2068, 255.2068, 
    255.2067, 255.2066, 255.2066, 255.2064, 255.2063, 255.2061, 255.2059, 
    255.2058, 255.2059, 255.2058, 255.2059, 255.2059, 255.2056, 255.2058, 
    255.2055, 255.2055, 255.2057, 255.2055, 255.2067, 255.2067, 255.2068, 
    255.2068, 255.2069, 255.2068, 255.2068, 255.2066, 255.2065, 255.2065, 
    255.2064, 255.2063, 255.2061, 255.206, 255.2058, 255.2058, 255.2058, 
    255.2058, 255.2059, 255.2058, 255.2057, 255.2058, 255.2056, 255.2056, 
    255.2055, 255.2056, 255.2067, 255.2067, 255.2067, 255.2066, 255.2067, 
    255.2065, 255.2065, 255.2062, 255.2063, 255.2061, 255.2063, 255.2063, 
    255.2061, 255.2063, 255.206, 255.2062, 255.2058, 255.206, 255.2058, 
    255.2058, 255.2057, 255.2057, 255.2056, 255.2055, 255.2055, 255.2054, 
    255.2066, 255.2065, 255.2065, 255.2065, 255.2064, 255.2063, 255.2061, 
    255.2061, 255.206, 255.206, 255.2062, 255.2061, 255.2065, 255.2064, 
    255.2065, 255.2066, 255.2061, 255.2064, 255.2059, 255.2061, 255.2057, 
    255.2059, 255.2055, 255.2054, 255.2052, 255.205, 255.2065, 255.2065, 
    255.2064, 255.2063, 255.2062, 255.2061, 255.206, 255.206, 255.2059, 
    255.2059, 255.206, 255.2059, 255.2064, 255.2061, 255.2065, 255.2064, 
    255.2063, 255.2064, 255.2062, 255.2061, 255.2059, 255.206, 255.2054, 
    255.2057, 255.2049, 255.2051, 255.2065, 255.2065, 255.2063, 255.2064, 
    255.206, 255.206, 255.2059, 255.2058, 255.2058, 255.2058, 255.2058, 
    255.2058, 255.2061, 255.2059, 255.2063, 255.2062, 255.2062, 255.2063, 
    255.2061, 255.206, 255.206, 255.2059, 255.2058, 255.206, 255.2054, 
    255.2058, 255.2064, 255.2063, 255.2063, 255.2063, 255.206, 255.2061, 
    255.2058, 255.2059, 255.2057, 255.2058, 255.2058, 255.2059, 255.2059, 
    255.2061, 255.2062, 255.2063, 255.2063, 255.2062, 255.206, 255.2058, 
    255.2058, 255.2057, 255.2061, 255.2059, 255.206, 255.2058, 255.2061, 
    255.2059, 255.2062, 255.2062, 255.2061, 255.2059, 255.2059, 255.2058, 
    255.2058, 255.206, 255.206, 255.2061, 255.2061, 255.2062, 255.2063, 
    255.2062, 255.2061, 255.206, 255.2058, 255.2057, 255.2056, 255.2055, 
    255.2056, 255.2054, 255.2056, 255.2052, 255.2059, 255.2056, 255.2061, 
    255.206, 255.2059, 255.2057, 255.2058, 255.2057, 255.206, 255.2062, 
    255.2062, 255.2063, 255.2062, 255.2062, 255.2061, 255.2062, 255.206, 
    255.2061, 255.2058, 255.2057, 255.2054, 255.2052, 255.205, 255.2049, 
    255.2049, 255.2049 ;

 TSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSOI =
  253.6968, 253.6987, 253.6983, 253.6998, 253.699, 253.7, 253.6972, 253.6987, 
    253.6978, 253.697, 253.7027, 253.6999, 253.7057, 253.7039, 253.7085, 
    253.7054, 253.7091, 253.7084, 253.7106, 253.71, 253.7126, 253.7109, 
    253.7141, 253.7122, 253.7125, 253.7108, 253.7005, 253.7023, 253.7004, 
    253.7006, 253.7005, 253.699, 253.6982, 253.6967, 253.697, 253.6981, 
    253.7007, 253.6999, 253.7021, 253.7021, 253.7046, 253.7035, 253.7077, 
    253.7065, 253.71, 253.7091, 253.7099, 253.7097, 253.7099, 253.7086, 
    253.7092, 253.7081, 253.7037, 253.705, 253.7011, 253.6987, 253.6973, 
    253.6962, 253.6963, 253.6966, 253.6981, 253.6996, 253.7007, 253.7014, 
    253.7021, 253.7042, 253.7054, 253.7079, 253.7075, 253.7083, 253.709, 
    253.7103, 253.7101, 253.7106, 253.7083, 253.7098, 253.7072, 253.7079, 
    253.7022, 253.7001, 253.6991, 253.6984, 253.6964, 253.6978, 253.6972, 
    253.6985, 253.6993, 253.6989, 253.7014, 253.7004, 253.7054, 253.7033, 
    253.7089, 253.7076, 253.7093, 253.7084, 253.7099, 253.7086, 253.7108, 
    253.7113, 253.711, 253.7123, 253.7085, 253.7099, 253.6989, 253.699, 
    253.6993, 253.6979, 253.6979, 253.6967, 253.6977, 253.6982, 253.6994, 
    253.7001, 253.7007, 253.7022, 253.7038, 253.706, 253.7077, 253.7088, 
    253.7081, 253.7087, 253.708, 253.7077, 253.7111, 253.7092, 253.7121, 
    253.712, 253.7106, 253.712, 253.699, 253.6987, 253.6974, 253.6984, 
    253.6965, 253.6975, 253.6981, 253.7004, 253.701, 253.7014, 253.7023, 
    253.7035, 253.7056, 253.7074, 253.7091, 253.709, 253.709, 253.7094, 
    253.7085, 253.7095, 253.7097, 253.7092, 253.7119, 253.7112, 253.712, 
    253.7115, 253.6988, 253.6994, 253.6991, 253.6997, 253.6992, 253.7012, 
    253.7018, 253.7046, 253.7035, 253.7053, 253.7037, 253.704, 253.7053, 
    253.7038, 253.7073, 253.7049, 253.7094, 253.7069, 253.7095, 253.7091, 
    253.7098, 253.7105, 253.7114, 253.713, 253.7126, 253.7139, 253.7003, 
    253.7011, 253.7011, 253.702, 253.7026, 253.7039, 253.7061, 253.7053, 
    253.7068, 253.7071, 253.7048, 253.7062, 253.7017, 253.7024, 253.702, 
    253.7004, 253.7055, 253.7029, 253.7077, 253.7063, 253.7104, 253.7083, 
    253.7124, 253.7141, 253.7157, 253.7176, 253.7016, 253.701, 253.7021, 
    253.7034, 253.7047, 253.7064, 253.7066, 253.7069, 253.7077, 253.7084, 
    253.7069, 253.7086, 253.7025, 253.7057, 253.7008, 253.7023, 253.7033, 
    253.7029, 253.7052, 253.7058, 253.708, 253.7068, 253.7136, 253.7106, 
    253.7191, 253.7167, 253.7009, 253.7016, 253.7042, 253.703, 253.7065, 
    253.7074, 253.7081, 253.709, 253.7091, 253.7096, 253.7087, 253.7096, 
    253.7064, 253.7078, 253.7039, 253.7048, 253.7044, 253.7039, 253.7054, 
    253.707, 253.707, 253.7075, 253.7088, 253.7065, 253.7139, 253.7093, 
    253.7024, 253.7038, 253.7041, 253.7035, 253.7073, 253.7059, 253.7096, 
    253.7086, 253.7102, 253.7094, 253.7093, 253.7083, 253.7076, 253.706, 
    253.7046, 253.7036, 253.7038, 253.705, 253.7071, 253.7091, 253.7086, 
    253.7101, 253.7062, 253.7078, 253.7072, 253.7088, 253.7053, 253.7082, 
    253.7045, 253.7048, 253.7059, 253.7079, 253.7084, 253.7089, 253.7086, 
    253.7071, 253.7069, 253.7059, 253.7056, 253.7048, 253.7041, 253.7047, 
    253.7053, 253.7071, 253.7087, 253.7105, 253.711, 253.7129, 253.7113, 
    253.714, 253.7116, 253.7157, 253.7084, 253.7116, 253.7059, 253.7066, 
    253.7076, 253.7102, 253.7088, 253.7104, 253.7069, 253.705, 253.7045, 
    253.7036, 253.7046, 253.7045, 253.7054, 253.7051, 253.7072, 253.7061, 
    253.7093, 253.7104, 253.7138, 253.7158, 253.7179, 253.7188, 253.7191, 
    253.7192,
  255.228, 255.2297, 255.2294, 255.2308, 255.23, 255.2309, 255.2283, 
    255.2298, 255.2289, 255.2282, 255.2335, 255.2309, 255.2363, 255.2346, 
    255.2389, 255.236, 255.2395, 255.2388, 255.2408, 255.2403, 255.2428, 
    255.2411, 255.2441, 255.2424, 255.2426, 255.241, 255.2314, 255.2331, 
    255.2313, 255.2316, 255.2314, 255.23, 255.2293, 255.2279, 255.2281, 
    255.2292, 255.2317, 255.2309, 255.233, 255.2329, 255.2352, 255.2342, 
    255.2381, 255.237, 255.2403, 255.2395, 255.2402, 255.24, 255.2402, 
    255.239, 255.2395, 255.2385, 255.2344, 255.2356, 255.232, 255.2298, 
    255.2284, 255.2274, 255.2276, 255.2278, 255.2292, 255.2305, 255.2316, 
    255.2322, 255.2329, 255.2348, 255.2359, 255.2384, 255.2379, 255.2387, 
    255.2394, 255.2406, 255.2404, 255.2409, 255.2387, 255.2401, 255.2377, 
    255.2384, 255.233, 255.2311, 255.2302, 255.2295, 255.2277, 255.2289, 
    255.2284, 255.2296, 255.2303, 255.23, 255.2323, 255.2314, 255.236, 
    255.234, 255.2393, 255.238, 255.2396, 255.2388, 255.2402, 255.2389, 
    255.2411, 255.2415, 255.2412, 255.2424, 255.2389, 255.2402, 255.23, 
    255.23, 255.2303, 255.229, 255.229, 255.2279, 255.2289, 255.2293, 
    255.2304, 255.231, 255.2316, 255.233, 255.2345, 255.2366, 255.2381, 
    255.2391, 255.2385, 255.2391, 255.2384, 255.2382, 255.2413, 255.2395, 
    255.2423, 255.2421, 255.2409, 255.2421, 255.2301, 255.2297, 255.2285, 
    255.2295, 255.2277, 255.2287, 255.2292, 255.2314, 255.2319, 255.2323, 
    255.2332, 255.2343, 255.2362, 255.2379, 255.2394, 255.2393, 255.2393, 
    255.2397, 255.2388, 255.2398, 255.24, 255.2396, 255.2421, 255.2414, 
    255.2421, 255.2417, 255.2298, 255.2304, 255.2301, 255.2307, 255.2303, 
    255.2321, 255.2327, 255.2353, 255.2342, 255.2359, 255.2344, 255.2347, 
    255.2359, 255.2345, 255.2377, 255.2355, 255.2397, 255.2374, 255.2398, 
    255.2394, 255.2401, 255.2408, 255.2416, 255.2431, 255.2427, 255.244, 
    255.2313, 255.232, 255.232, 255.2328, 255.2334, 255.2346, 255.2367, 
    255.2359, 255.2373, 255.2376, 255.2355, 255.2368, 255.2325, 255.2332, 
    255.2328, 255.2313, 255.2361, 255.2336, 255.2381, 255.2368, 255.2407, 
    255.2387, 255.2425, 255.2441, 255.2457, 255.2474, 255.2325, 255.2319, 
    255.2329, 255.2341, 255.2353, 255.2369, 255.2371, 255.2374, 255.2381, 
    255.2388, 255.2374, 255.2389, 255.2333, 255.2363, 255.2317, 255.2331, 
    255.234, 255.2336, 255.2358, 255.2363, 255.2384, 255.2373, 255.2437, 
    255.2409, 255.2488, 255.2466, 255.2318, 255.2325, 255.2348, 255.2337, 
    255.237, 255.2378, 255.2385, 255.2393, 255.2394, 255.2399, 255.2391, 
    255.2399, 255.2369, 255.2382, 255.2346, 255.2355, 255.2351, 255.2346, 
    255.236, 255.2374, 255.2375, 255.238, 255.2392, 255.237, 255.244, 
    255.2396, 255.2332, 255.2345, 255.2347, 255.2342, 255.2377, 255.2365, 
    255.2399, 255.239, 255.2405, 255.2397, 255.2396, 255.2386, 255.238, 
    255.2365, 255.2353, 255.2343, 255.2345, 255.2356, 255.2375, 255.2394, 
    255.239, 255.2404, 255.2368, 255.2383, 255.2377, 255.2392, 255.2359, 
    255.2386, 255.2352, 255.2355, 255.2364, 255.2383, 255.2388, 255.2393, 
    255.239, 255.2376, 255.2374, 255.2364, 255.2361, 255.2354, 255.2348, 
    255.2354, 255.2359, 255.2376, 255.2391, 255.2408, 255.2412, 255.2431, 
    255.2415, 255.244, 255.2418, 255.2457, 255.2388, 255.2418, 255.2365, 
    255.2371, 255.2381, 255.2405, 255.2392, 255.2407, 255.2374, 255.2356, 
    255.2352, 255.2344, 255.2352, 255.2352, 255.236, 255.2357, 255.2377, 
    255.2366, 255.2396, 255.2407, 255.2438, 255.2457, 255.2477, 255.2486, 
    255.2489, 255.249,
  257.293, 257.2944, 257.2942, 257.2953, 257.2947, 257.2954, 257.2933, 
    257.2945, 257.2937, 257.2932, 257.2974, 257.2953, 257.2997, 257.2984, 
    257.3018, 257.2995, 257.3023, 257.3018, 257.3034, 257.3029, 257.305, 
    257.3036, 257.3061, 257.3047, 257.3049, 257.3036, 257.2958, 257.2971, 
    257.2957, 257.2959, 257.2958, 257.2947, 257.2941, 257.2929, 257.2932, 
    257.294, 257.296, 257.2953, 257.297, 257.297, 257.2989, 257.298, 
    257.3012, 257.3003, 257.303, 257.3023, 257.3029, 257.3028, 257.3029, 
    257.3019, 257.3024, 257.3015, 257.2982, 257.2992, 257.2962, 257.2945, 
    257.2934, 257.2926, 257.2927, 257.2929, 257.294, 257.2951, 257.2959, 
    257.2964, 257.297, 257.2986, 257.2994, 257.3014, 257.3011, 257.3016, 
    257.3022, 257.3032, 257.303, 257.3035, 257.3016, 257.3029, 257.3009, 
    257.3014, 257.2971, 257.2955, 257.2948, 257.2942, 257.2928, 257.2938, 
    257.2934, 257.2943, 257.2949, 257.2946, 257.2964, 257.2957, 257.2995, 
    257.2979, 257.3022, 257.3011, 257.3024, 257.3018, 257.3029, 257.3019, 
    257.3036, 257.304, 257.3037, 257.3047, 257.3018, 257.3029, 257.2946, 
    257.2946, 257.2949, 257.2939, 257.2938, 257.2929, 257.2937, 257.2941, 
    257.295, 257.2955, 257.296, 257.2971, 257.2982, 257.3, 257.3012, 257.302, 
    257.3015, 257.302, 257.3015, 257.3012, 257.3039, 257.3024, 257.3046, 
    257.3045, 257.3035, 257.3045, 257.2947, 257.2944, 257.2935, 257.2942, 
    257.2928, 257.2936, 257.294, 257.2957, 257.2961, 257.2965, 257.2972, 
    257.2981, 257.2996, 257.301, 257.3023, 257.3022, 257.3022, 257.3025, 
    257.3018, 257.3026, 257.3027, 257.3024, 257.3045, 257.3039, 257.3045, 
    257.3041, 257.2945, 257.295, 257.2947, 257.2952, 257.2949, 257.2963, 
    257.2968, 257.2989, 257.298, 257.2994, 257.2982, 257.2984, 257.2994, 
    257.2982, 257.3009, 257.2991, 257.3025, 257.3006, 257.3026, 257.3023, 
    257.3029, 257.3034, 257.304, 257.3052, 257.305, 257.306, 257.2957, 
    257.2963, 257.2962, 257.2969, 257.2973, 257.2984, 257.3, 257.2994, 
    257.3006, 257.3008, 257.299, 257.3001, 257.2967, 257.2972, 257.2969, 
    257.2957, 257.2995, 257.2975, 257.3012, 257.3001, 257.3033, 257.3017, 
    257.3048, 257.3061, 257.3074, 257.3089, 257.2966, 257.2962, 257.2969, 
    257.2979, 257.2989, 257.3002, 257.3004, 257.3006, 257.3012, 257.3017, 
    257.3007, 257.3019, 257.2973, 257.2997, 257.2961, 257.2971, 257.2979, 
    257.2976, 257.2993, 257.2997, 257.3014, 257.3006, 257.3058, 257.3035, 
    257.31, 257.3082, 257.2961, 257.2966, 257.2986, 257.2976, 257.3003, 
    257.301, 257.3015, 257.3022, 257.3023, 257.3027, 257.302, 257.3026, 
    257.3002, 257.3013, 257.2983, 257.299, 257.2987, 257.2984, 257.2995, 
    257.3007, 257.3007, 257.3011, 257.3021, 257.3003, 257.306, 257.3025, 
    257.2972, 257.2983, 257.2985, 257.298, 257.3009, 257.2999, 257.3027, 
    257.3019, 257.3032, 257.3025, 257.3024, 257.3016, 257.3011, 257.2999, 
    257.2989, 257.2981, 257.2983, 257.2992, 257.3008, 257.3022, 257.3019, 
    257.3031, 257.3001, 257.3013, 257.3008, 257.3021, 257.2994, 257.3016, 
    257.2988, 257.2991, 257.2998, 257.3014, 257.3018, 257.3022, 257.3019, 
    257.3008, 257.3006, 257.2998, 257.2996, 257.299, 257.2985, 257.299, 
    257.2994, 257.3008, 257.302, 257.3034, 257.3037, 257.3052, 257.304, 
    257.3061, 257.3042, 257.3074, 257.3018, 257.3042, 257.2999, 257.3004, 
    257.3012, 257.3031, 257.3021, 257.3033, 257.3006, 257.2992, 257.2988, 
    257.2982, 257.2989, 257.2988, 257.2995, 257.2993, 257.3008, 257.3, 
    257.3024, 257.3033, 257.3059, 257.3075, 257.3091, 257.3098, 257.31, 
    257.3101,
  259.7986, 259.7994, 259.7992, 259.7999, 259.7995, 259.7999, 259.7987, 
    259.7994, 259.799, 259.7986, 259.8011, 259.7999, 259.8025, 259.8017, 
    259.8037, 259.8023, 259.804, 259.8037, 259.8047, 259.8044, 259.8056, 
    259.8048, 259.8063, 259.8055, 259.8056, 259.8048, 259.8001, 259.801, 
    259.8001, 259.8002, 259.8002, 259.7995, 259.7992, 259.7985, 259.7986, 
    259.7991, 259.8003, 259.7999, 259.8009, 259.8009, 259.802, 259.8015, 
    259.8034, 259.8028, 259.8044, 259.804, 259.8044, 259.8043, 259.8044, 
    259.8038, 259.804, 259.8036, 259.8016, 259.8021, 259.8004, 259.7994, 
    259.7987, 259.7983, 259.7983, 259.7985, 259.7991, 259.7997, 259.8002, 
    259.8005, 259.8008, 259.8018, 259.8023, 259.8035, 259.8033, 259.8036, 
    259.804, 259.8046, 259.8045, 259.8047, 259.8036, 259.8044, 259.8032, 
    259.8035, 259.8009, 259.8, 259.7996, 259.7992, 259.7984, 259.799, 
    259.7987, 259.7993, 259.7997, 259.7995, 259.8005, 259.8001, 259.8023, 
    259.8014, 259.8039, 259.8033, 259.8041, 259.8037, 259.8044, 259.8038, 
    259.8048, 259.805, 259.8049, 259.8055, 259.8037, 259.8044, 259.7995, 
    259.7995, 259.7996, 259.799, 259.799, 259.7985, 259.799, 259.7992, 
    259.7997, 259.8, 259.8003, 259.8009, 259.8016, 259.8026, 259.8033, 
    259.8039, 259.8036, 259.8038, 259.8035, 259.8034, 259.805, 259.804, 
    259.8054, 259.8053, 259.8047, 259.8053, 259.7995, 259.7993, 259.7988, 
    259.7992, 259.7984, 259.7989, 259.7991, 259.8001, 259.8004, 259.8006, 
    259.801, 259.8015, 259.8024, 259.8032, 259.804, 259.804, 259.804, 
    259.8041, 259.8037, 259.8042, 259.8043, 259.8041, 259.8053, 259.805, 
    259.8053, 259.8051, 259.7994, 259.7997, 259.7995, 259.7998, 259.7996, 
    259.8005, 259.8008, 259.802, 259.8015, 259.8023, 259.8016, 259.8017, 
    259.8023, 259.8016, 259.8032, 259.8021, 259.8041, 259.803, 259.8042, 
    259.804, 259.8044, 259.8047, 259.8051, 259.8058, 259.8056, 259.8062, 
    259.8001, 259.8004, 259.8004, 259.8008, 259.8011, 259.8017, 259.8026, 
    259.8023, 259.803, 259.8031, 259.8021, 259.8027, 259.8007, 259.801, 
    259.8008, 259.8001, 259.8024, 259.8012, 259.8034, 259.8027, 259.8046, 
    259.8036, 259.8055, 259.8063, 259.8071, 259.808, 259.8006, 259.8004, 
    259.8008, 259.8014, 259.802, 259.8028, 259.8029, 259.803, 259.8034, 
    259.8037, 259.803, 259.8038, 259.8011, 259.8025, 259.8003, 259.8009, 
    259.8014, 259.8012, 259.8022, 259.8025, 259.8035, 259.803, 259.8061, 
    259.8047, 259.8087, 259.8076, 259.8003, 259.8007, 259.8018, 259.8012, 
    259.8028, 259.8032, 259.8035, 259.804, 259.804, 259.8042, 259.8038, 
    259.8042, 259.8028, 259.8034, 259.8017, 259.8021, 259.8019, 259.8017, 
    259.8023, 259.803, 259.8031, 259.8033, 259.8039, 259.8028, 259.8063, 
    259.8041, 259.801, 259.8016, 259.8017, 259.8015, 259.8032, 259.8026, 
    259.8042, 259.8038, 259.8045, 259.8041, 259.8041, 259.8036, 259.8033, 
    259.8026, 259.802, 259.8015, 259.8016, 259.8021, 259.8031, 259.804, 
    259.8038, 259.8045, 259.8027, 259.8034, 259.8032, 259.8039, 259.8023, 
    259.8036, 259.8019, 259.8021, 259.8026, 259.8035, 259.8037, 259.8039, 
    259.8038, 259.8031, 259.803, 259.8025, 259.8024, 259.8021, 259.8018, 
    259.802, 259.8023, 259.8031, 259.8038, 259.8047, 259.8049, 259.8058, 
    259.805, 259.8063, 259.8052, 259.8071, 259.8037, 259.8052, 259.8026, 
    259.8029, 259.8033, 259.8045, 259.8039, 259.8046, 259.803, 259.8022, 
    259.8019, 259.8015, 259.802, 259.8019, 259.8023, 259.8022, 259.8031, 
    259.8026, 259.8041, 259.8046, 259.8062, 259.8071, 259.8081, 259.8086, 
    259.8087, 259.8088,
  262.0124, 262.0125, 262.0125, 262.0127, 262.0126, 262.0127, 262.0124, 
    262.0126, 262.0125, 262.0124, 262.013, 262.0127, 262.0134, 262.0132, 
    262.0137, 262.0133, 262.0138, 262.0137, 262.014, 262.0139, 262.0143, 
    262.014, 262.0144, 262.0142, 262.0142, 262.014, 262.0128, 262.013, 
    262.0127, 262.0128, 262.0128, 262.0126, 262.0125, 262.0123, 262.0124, 
    262.0125, 262.0128, 262.0127, 262.0129, 262.0129, 262.0132, 262.0131, 
    262.0136, 262.0135, 262.0139, 262.0138, 262.0139, 262.0139, 262.0139, 
    262.0137, 262.0138, 262.0137, 262.0131, 262.0133, 262.0128, 262.0126, 
    262.0124, 262.0123, 262.0123, 262.0123, 262.0125, 262.0126, 262.0128, 
    262.0128, 262.0129, 262.0132, 262.0133, 262.0136, 262.0136, 262.0137, 
    262.0138, 262.0139, 262.0139, 262.014, 262.0137, 262.0139, 262.0135, 
    262.0136, 262.0129, 262.0127, 262.0126, 262.0125, 262.0123, 262.0125, 
    262.0124, 262.0125, 262.0126, 262.0126, 262.0128, 262.0128, 262.0133, 
    262.0131, 262.0138, 262.0136, 262.0138, 262.0137, 262.0139, 262.0137, 
    262.014, 262.0141, 262.014, 262.0142, 262.0137, 262.0139, 262.0126, 
    262.0126, 262.0126, 262.0125, 262.0125, 262.0123, 262.0125, 262.0125, 
    262.0126, 262.0127, 262.0128, 262.0129, 262.0131, 262.0134, 262.0136, 
    262.0137, 262.0137, 262.0137, 262.0136, 262.0136, 262.014, 262.0138, 
    262.0142, 262.0142, 262.014, 262.0142, 262.0126, 262.0125, 262.0124, 
    262.0125, 262.0123, 262.0124, 262.0125, 262.0128, 262.0128, 262.0128, 
    262.013, 262.0131, 262.0133, 262.0136, 262.0138, 262.0138, 262.0138, 
    262.0138, 262.0137, 262.0138, 262.0139, 262.0138, 262.0142, 262.0141, 
    262.0142, 262.0141, 262.0126, 262.0126, 262.0126, 262.0127, 262.0126, 
    262.0128, 262.0129, 262.0132, 262.0131, 262.0133, 262.0131, 262.0132, 
    262.0133, 262.0131, 262.0135, 262.0133, 262.0138, 262.0135, 262.0139, 
    262.0138, 262.0139, 262.014, 262.0141, 262.0143, 262.0143, 262.0144, 
    262.0127, 262.0128, 262.0128, 262.0129, 262.013, 262.0132, 262.0134, 
    262.0133, 262.0135, 262.0135, 262.0132, 262.0134, 262.0129, 262.013, 
    262.0129, 262.0128, 262.0133, 262.013, 262.0136, 262.0134, 262.0139, 
    262.0137, 262.0142, 262.0144, 262.0147, 262.015, 262.0129, 262.0128, 
    262.0129, 262.0131, 262.0132, 262.0135, 262.0135, 262.0135, 262.0136, 
    262.0137, 262.0135, 262.0137, 262.013, 262.0134, 262.0128, 262.013, 
    262.0131, 262.013, 262.0133, 262.0134, 262.0136, 262.0135, 262.0144, 
    262.014, 262.0152, 262.0148, 262.0128, 262.0129, 262.0132, 262.013, 
    262.0135, 262.0136, 262.0136, 262.0138, 262.0138, 262.0139, 262.0137, 
    262.0139, 262.0135, 262.0136, 262.0132, 262.0132, 262.0132, 262.0132, 
    262.0133, 262.0135, 262.0135, 262.0136, 262.0138, 262.0135, 262.0144, 
    262.0138, 262.013, 262.0131, 262.0132, 262.0131, 262.0135, 262.0134, 
    262.0139, 262.0137, 262.0139, 262.0138, 262.0138, 262.0137, 262.0136, 
    262.0134, 262.0132, 262.0131, 262.0132, 262.0133, 262.0135, 262.0138, 
    262.0137, 262.0139, 262.0134, 262.0136, 262.0135, 262.0138, 262.0133, 
    262.0137, 262.0132, 262.0132, 262.0134, 262.0136, 262.0137, 262.0138, 
    262.0137, 262.0135, 262.0135, 262.0134, 262.0133, 262.0132, 262.0132, 
    262.0132, 262.0133, 262.0135, 262.0137, 262.014, 262.014, 262.0143, 
    262.0141, 262.0144, 262.0141, 262.0147, 262.0137, 262.0141, 262.0134, 
    262.0135, 262.0136, 262.0139, 262.0138, 262.0139, 262.0135, 262.0133, 
    262.0132, 262.0131, 262.0132, 262.0132, 262.0133, 262.0133, 262.0135, 
    262.0134, 262.0138, 262.0139, 262.0144, 262.0147, 262.015, 262.0151, 
    262.0152, 262.0152,
  262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 262.9993, 
    262.9993, 262.9993,
  263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 263.1448, 
    263.1448, 263.1448,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15 ;

 TSOI_10CM =
  263.1089, 263.1212, 263.1189, 263.1288, 263.1233, 263.1298, 263.1115, 
    263.1217, 263.1152, 263.1101, 263.1478, 263.1292, 263.1672, 263.1554, 
    263.1851, 263.1653, 263.189, 263.1846, 263.1981, 263.1942, 263.2114, 
    263.1999, 263.2203, 263.2086, 263.2105, 263.1995, 263.133, 263.1455, 
    263.1322, 263.134, 263.1332, 263.1234, 263.1184, 263.108, 263.1099, 
    263.1176, 263.1348, 263.129, 263.1437, 263.1434, 263.1598, 263.1524, 
    263.1798, 263.1721, 263.1944, 263.1888, 263.1941, 263.1925, 263.1941, 
    263.1859, 263.1895, 263.1823, 263.1537, 263.1621, 263.1371, 263.1219, 
    263.1119, 263.1047, 263.1057, 263.1077, 263.1176, 263.1269, 263.134, 
    263.1387, 263.1433, 263.1573, 263.1648, 263.1814, 263.1784, 263.1834, 
    263.1882, 263.1962, 263.1949, 263.1984, 263.1833, 263.1934, 263.1767, 
    263.1813, 263.1445, 263.1306, 263.1245, 263.1193, 263.1065, 263.1154, 
    263.1119, 263.1202, 263.1254, 263.1228, 263.1388, 263.1326, 263.1652, 
    263.1512, 263.1877, 263.179, 263.1897, 263.1843, 263.1936, 263.1852, 
    263.1998, 263.2029, 263.2007, 263.209, 263.1848, 263.1941, 263.1228, 
    263.1232, 263.1252, 263.1165, 263.1159, 263.108, 263.1151, 263.1181, 
    263.1258, 263.1302, 263.1346, 263.144, 263.1544, 263.1691, 263.1796, 
    263.1866, 263.1823, 263.1861, 263.1819, 263.1799, 263.2017, 263.1895, 
    263.2079, 263.2068, 263.1985, 263.207, 263.1235, 263.1211, 263.1125, 
    263.1192, 263.1071, 263.1139, 263.1177, 263.1327, 263.136, 263.1391, 
    263.1451, 263.1527, 263.1662, 263.1779, 263.1885, 263.1877, 263.188, 
    263.1904, 263.1845, 263.1913, 263.1924, 263.1895, 263.2067, 263.2018, 
    263.2068, 263.2036, 263.1219, 263.1259, 263.1237, 263.1279, 263.125, 
    263.1379, 263.1418, 263.16, 263.1526, 263.1645, 263.1538, 263.1557, 
    263.1648, 263.1544, 263.1772, 263.1617, 263.1905, 263.175, 263.1914, 
    263.1885, 263.1933, 263.1977, 263.2032, 263.2133, 263.2109, 263.2194, 
    263.132, 263.1373, 263.1369, 263.1424, 263.1465, 263.1554, 263.1696, 
    263.1642, 263.174, 263.176, 263.1611, 263.1703, 263.1409, 263.1456, 
    263.1428, 263.1324, 263.1654, 263.1485, 263.1797, 263.1706, 263.1971, 
    263.184, 263.2097, 263.2206, 263.2309, 263.2428, 263.1402, 263.1367, 
    263.1431, 263.1519, 263.1602, 263.1712, 263.1723, 263.1743, 263.1797, 
    263.1841, 263.175, 263.1852, 263.1467, 263.1669, 263.1353, 263.1448, 
    263.1514, 263.1485, 263.1636, 263.1672, 263.1816, 263.1742, 263.2178, 
    263.1986, 263.252, 263.2371, 263.1354, 263.1402, 263.157, 263.149, 
    263.1719, 263.1775, 263.1821, 263.1878, 263.1884, 263.1919, 263.1863, 
    263.1917, 263.1712, 263.1804, 263.1551, 263.1613, 263.1584, 263.1554, 
    263.1649, 263.1751, 263.1754, 263.1786, 263.1877, 263.172, 263.2203, 
    263.1905, 263.1455, 263.1548, 263.1561, 263.1525, 263.1769, 263.1681, 
    263.1918, 263.1855, 263.1958, 263.1907, 263.1899, 263.1833, 263.1791, 
    263.1685, 263.1599, 263.1531, 263.1547, 263.1622, 263.1758, 263.1885, 
    263.1857, 263.195, 263.1703, 263.1807, 263.1766, 263.1872, 263.1641, 
    263.1837, 263.1591, 263.1612, 263.1679, 263.1814, 263.1844, 263.1875, 
    263.1856, 263.1761, 263.1746, 263.1678, 263.1659, 263.1608, 263.1565, 
    263.1604, 263.1645, 263.1761, 263.1865, 263.1978, 263.2005, 263.2135, 
    263.2029, 263.2204, 263.2054, 263.2314, 263.1848, 263.2051, 263.1683, 
    263.1723, 263.1795, 263.1959, 263.1871, 263.1974, 263.1745, 263.1624, 
    263.1593, 263.1535, 263.1595, 263.159, 263.1647, 263.1628, 263.1765, 
    263.1692, 263.1899, 263.1974, 263.2185, 263.2314, 263.2445, 263.2503, 
    263.2521, 263.2528 ;

 TSOI_ICE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TV =
  253.595, 253.5958, 253.5956, 253.5963, 253.5959, 253.5963, 253.5952, 
    253.5958, 253.5954, 253.5951, 253.5975, 253.5963, 253.5988, 253.598, 
    253.6, 253.5987, 253.6002, 253.5999, 253.6008, 253.6006, 253.6017, 
    253.601, 253.6023, 253.6015, 253.6017, 253.6009, 253.5966, 253.5974, 
    253.5965, 253.5966, 253.5966, 253.5959, 253.5956, 253.5949, 253.595, 
    253.5955, 253.5967, 253.5963, 253.5973, 253.5973, 253.5983, 253.5978, 
    253.5996, 253.5991, 253.6006, 253.6002, 253.6006, 253.6005, 253.6006, 
    253.6, 253.6003, 253.5998, 253.5979, 253.5985, 253.5968, 253.5958, 
    253.5952, 253.5947, 253.5948, 253.5949, 253.5956, 253.5962, 253.5966, 
    253.5969, 253.5972, 253.5981, 253.5986, 253.5997, 253.5995, 253.5999, 
    253.6002, 253.6007, 253.6006, 253.6009, 253.5999, 253.6005, 253.5994, 
    253.5997, 253.5973, 253.5964, 253.596, 253.5957, 253.5948, 253.5954, 
    253.5952, 253.5957, 253.5961, 253.5959, 253.597, 253.5965, 253.5987, 
    253.5978, 253.6002, 253.5996, 253.6003, 253.5999, 253.6005, 253.6, 
    253.601, 253.6012, 253.601, 253.6016, 253.6, 253.6006, 253.5959, 
    253.5959, 253.5961, 253.5955, 253.5954, 253.5949, 253.5954, 253.5956, 
    253.5961, 253.5964, 253.5967, 253.5973, 253.598, 253.5989, 253.5996, 
    253.6001, 253.5998, 253.6001, 253.5998, 253.5996, 253.6011, 253.6003, 
    253.6015, 253.6014, 253.6009, 253.6014, 253.5959, 253.5958, 253.5952, 
    253.5957, 253.5949, 253.5953, 253.5956, 253.5965, 253.5968, 253.597, 
    253.5974, 253.5979, 253.5987, 253.5995, 253.6002, 253.6002, 253.6002, 
    253.6003, 253.5999, 253.6004, 253.6005, 253.6003, 253.6014, 253.6011, 
    253.6014, 253.6012, 253.5958, 253.5961, 253.596, 253.5962, 253.596, 
    253.5969, 253.5971, 253.5983, 253.5979, 253.5986, 253.5979, 253.5981, 
    253.5986, 253.598, 253.5995, 253.5984, 253.6003, 253.5993, 253.6004, 
    253.6002, 253.6005, 253.6008, 253.6012, 253.6019, 253.6017, 253.6023, 
    253.5965, 253.5968, 253.5968, 253.5972, 253.5975, 253.598, 253.599, 
    253.5986, 253.5993, 253.5994, 253.5984, 253.599, 253.5971, 253.5974, 
    253.5972, 253.5965, 253.5987, 253.5976, 253.5996, 253.599, 253.6008, 
    253.5999, 253.6016, 253.6023, 253.603, 253.6038, 253.597, 253.5968, 
    253.5972, 253.5978, 253.5984, 253.5991, 253.5992, 253.5993, 253.5996, 
    253.5999, 253.5993, 253.6, 253.5974, 253.5988, 253.5967, 253.5973, 
    253.5978, 253.5976, 253.5986, 253.5988, 253.5997, 253.5993, 253.6021, 
    253.6009, 253.6044, 253.6034, 253.5967, 253.597, 253.5981, 253.5976, 
    253.5991, 253.5995, 253.5998, 253.6002, 253.6002, 253.6004, 253.6001, 
    253.6004, 253.5991, 253.5997, 253.598, 253.5984, 253.5983, 253.598, 
    253.5987, 253.5993, 253.5993, 253.5995, 253.6001, 253.5991, 253.6023, 
    253.6003, 253.5974, 253.598, 253.5981, 253.5979, 253.5994, 253.5989, 
    253.6004, 253.6, 253.6007, 253.6004, 253.6003, 253.5999, 253.5996, 
    253.5989, 253.5983, 253.5979, 253.598, 253.5985, 253.5994, 253.6002, 
    253.6, 253.6006, 253.599, 253.5997, 253.5994, 253.6001, 253.5986, 
    253.5999, 253.5983, 253.5984, 253.5989, 253.5997, 253.5999, 253.6001, 
    253.6, 253.5994, 253.5993, 253.5988, 253.5987, 253.5984, 253.5981, 
    253.5984, 253.5986, 253.5994, 253.6001, 253.6008, 253.601, 253.6019, 
    253.6012, 253.6023, 253.6013, 253.603, 253.5999, 253.6013, 253.5989, 
    253.5992, 253.5996, 253.6007, 253.6001, 253.6008, 253.5993, 253.5985, 
    253.5983, 253.5979, 253.5983, 253.5983, 253.5986, 253.5985, 253.5994, 
    253.5989, 253.6003, 253.6008, 253.6022, 253.6031, 253.6039, 253.6043, 
    253.6044, 253.6045 ;

 TWS =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 T_SCALAR =
  0.1457035, 0.1457024, 0.1457026, 0.1457018, 0.1457022, 0.1457017, 
    0.1457033, 0.1457024, 0.1457029, 0.1457034, 0.1457002, 0.1457017, 
    0.1456987, 0.1456996, 0.1456974, 0.1456989, 0.1456971, 0.1456974, 
    0.1456965, 0.1456967, 0.1456956, 0.1456964, 0.145695, 0.1456958, 
    0.1456957, 0.1456964, 0.1457014, 0.1457004, 0.1457015, 0.1457013, 
    0.1457014, 0.1457022, 0.1457027, 0.1457036, 0.1457034, 0.1457027, 
    0.1457013, 0.1457018, 0.1457005, 0.1457006, 0.1456993, 0.1456999, 
    0.1456978, 0.1456984, 0.1456967, 0.1456971, 0.1456967, 0.1456968, 
    0.1456967, 0.1456973, 0.1456971, 0.1456976, 0.1456998, 0.1456991, 
    0.1457011, 0.1457024, 0.1457032, 0.1457038, 0.1457037, 0.1457036, 
    0.1457027, 0.1457019, 0.1457013, 0.145701, 0.1457006, 0.1456995, 
    0.1456989, 0.1456976, 0.1456978, 0.1456975, 0.1456971, 0.1456966, 
    0.1456967, 0.1456964, 0.1456975, 0.1456968, 0.145698, 0.1456977, 
    0.1457005, 0.1457016, 0.1457021, 0.1457026, 0.1457037, 0.1457029, 
    0.1457032, 0.1457025, 0.145702, 0.1457023, 0.1457009, 0.1457015, 
    0.1456989, 0.1457, 0.1456972, 0.1456978, 0.145697, 0.1456974, 0.1456968, 
    0.1456974, 0.1456964, 0.1456961, 0.1456963, 0.1456957, 0.1456974, 
    0.1456967, 0.1457023, 0.1457022, 0.1457021, 0.1457028, 0.1457029, 
    0.1457036, 0.1457029, 0.1457027, 0.145702, 0.1457016, 0.1457013, 
    0.1457005, 0.1456997, 0.1456986, 0.1456978, 0.1456973, 0.1456976, 
    0.1456973, 0.1456976, 0.1456977, 0.1456962, 0.1456971, 0.1456958, 
    0.1456959, 0.1456964, 0.1456959, 0.1457022, 0.1457024, 0.1457032, 
    0.1457026, 0.1457036, 0.145703, 0.1457027, 0.1457015, 0.1457012, 
    0.1457009, 0.1457004, 0.1456998, 0.1456988, 0.1456979, 0.1456971, 
    0.1456972, 0.1456972, 0.145697, 0.1456974, 0.1456969, 0.1456969, 
    0.1456971, 0.1456959, 0.1456962, 0.1456959, 0.1456961, 0.1457024, 
    0.145702, 0.1457022, 0.1457019, 0.1457021, 0.145701, 0.1457007, 
    0.1456993, 0.1456998, 0.1456989, 0.1456998, 0.1456996, 0.1456989, 
    0.1456997, 0.145698, 0.1456991, 0.145697, 0.1456981, 0.1456969, 
    0.1456971, 0.1456968, 0.1456965, 0.1456961, 0.1456955, 0.1456956, 
    0.1456951, 0.1457015, 0.1457011, 0.1457011, 0.1457007, 0.1457003, 
    0.1456996, 0.1456985, 0.1456989, 0.1456982, 0.145698, 0.1456992, 
    0.1456985, 0.1457008, 0.1457004, 0.1457006, 0.1457015, 0.1456989, 
    0.1457002, 0.1456978, 0.1456985, 0.1456965, 0.1456975, 0.1456957, 
    0.145695, 0.1456944, 0.1456938, 0.1457008, 0.1457011, 0.1457006, 
    0.1456999, 0.1456992, 0.1456984, 0.1456983, 0.1456982, 0.1456978, 
    0.1456974, 0.1456981, 0.1456974, 0.1457003, 0.1456987, 0.1457012, 
    0.1457005, 0.1456999, 0.1457002, 0.145699, 0.1456987, 0.1456976, 
    0.1456982, 0.1456952, 0.1456964, 0.1456933, 0.1456941, 0.1457012, 
    0.1457008, 0.1456995, 0.1457001, 0.1456984, 0.1456979, 0.1456976, 
    0.1456972, 0.1456971, 0.1456969, 0.1456973, 0.1456969, 0.1456984, 
    0.1456977, 0.1456997, 0.1456992, 0.1456994, 0.1456996, 0.1456989, 
    0.1456981, 0.1456981, 0.1456978, 0.1456972, 0.1456984, 0.1456951, 
    0.145697, 0.1457004, 0.1456997, 0.1456996, 0.1456999, 0.145698, 
    0.1456987, 0.1456969, 0.1456974, 0.1456966, 0.145697, 0.145697, 
    0.1456975, 0.1456978, 0.1456986, 0.1456993, 0.1456998, 0.1456997, 
    0.1456991, 0.1456981, 0.1456971, 0.1456973, 0.1456967, 0.1456985, 
    0.1456977, 0.145698, 0.1456972, 0.1456989, 0.1456975, 0.1456993, 
    0.1456992, 0.1456987, 0.1456976, 0.1456974, 0.1456972, 0.1456973, 
    0.145698, 0.1456982, 0.1456987, 0.1456988, 0.1456992, 0.1456995, 
    0.1456992, 0.1456989, 0.145698, 0.1456973, 0.1456965, 0.1456963, 
    0.1456955, 0.1456961, 0.145695, 0.145696, 0.1456944, 0.1456974, 0.145696, 
    0.1456986, 0.1456983, 0.1456978, 0.1456966, 0.1456972, 0.1456965, 
    0.1456982, 0.1456991, 0.1456993, 0.1456998, 0.1456993, 0.1456994, 
    0.1456989, 0.1456991, 0.145698, 0.1456986, 0.145697, 0.1456965, 
    0.1456952, 0.1456944, 0.1456937, 0.1456934, 0.1456933, 0.1456933,
  0.1513279, 0.1513324, 0.1513316, 0.1513352, 0.1513332, 0.1513356, 
    0.1513288, 0.1513326, 0.1513302, 0.1513283, 0.1513422, 0.1513354, 
    0.1513497, 0.1513453, 0.1513565, 0.151349, 0.1513581, 0.1513564, 
    0.1513617, 0.1513602, 0.1513669, 0.1513624, 0.1513705, 0.1513658, 
    0.1513665, 0.1513623, 0.1513368, 0.1513413, 0.1513366, 0.1513372, 
    0.1513369, 0.1513332, 0.1513313, 0.1513276, 0.1513283, 0.1513311, 
    0.1513375, 0.1513353, 0.1513409, 0.1513408, 0.1513469, 0.1513442, 
    0.1513546, 0.1513516, 0.1513603, 0.1513581, 0.1513601, 0.1513595, 
    0.1513602, 0.1513569, 0.1513583, 0.1513555, 0.1513447, 0.1513478, 
    0.1513384, 0.1513326, 0.151329, 0.1513264, 0.1513267, 0.1513274, 
    0.1513311, 0.1513346, 0.1513372, 0.151339, 0.1513408, 0.1513459, 
    0.1513488, 0.1513551, 0.151354, 0.1513559, 0.1513578, 0.151361, 
    0.1513605, 0.1513618, 0.1513559, 0.1513598, 0.1513534, 0.1513551, 
    0.151341, 0.1513359, 0.1513336, 0.1513317, 0.151327, 0.1513302, 0.151329, 
    0.1513321, 0.151334, 0.1513331, 0.1513391, 0.1513367, 0.1513489, 
    0.1513437, 0.1513576, 0.1513543, 0.1513584, 0.1513563, 0.1513599, 
    0.1513567, 0.1513624, 0.1513636, 0.1513627, 0.151366, 0.1513565, 
    0.1513601, 0.151333, 0.1513332, 0.1513339, 0.1513306, 0.1513305, 
    0.1513275, 0.1513302, 0.1513313, 0.1513342, 0.1513358, 0.1513374, 
    0.151341, 0.1513449, 0.1513505, 0.1513545, 0.1513572, 0.1513555, 
    0.151357, 0.1513554, 0.1513546, 0.1513631, 0.1513583, 0.1513656, 
    0.1513652, 0.1513619, 0.1513652, 0.1513333, 0.1513324, 0.1513292, 
    0.1513317, 0.1513272, 0.1513297, 0.1513311, 0.1513367, 0.151338, 
    0.1513391, 0.1513414, 0.1513443, 0.1513494, 0.1513538, 0.151358, 
    0.1513577, 0.1513578, 0.1513587, 0.1513564, 0.1513591, 0.1513595, 
    0.1513583, 0.1513651, 0.1513632, 0.1513652, 0.1513639, 0.1513327, 
    0.1513342, 0.1513334, 0.1513349, 0.1513338, 0.1513387, 0.1513401, 
    0.151347, 0.1513442, 0.1513487, 0.1513447, 0.1513454, 0.1513487, 
    0.1513449, 0.1513535, 0.1513476, 0.1513587, 0.1513526, 0.1513591, 
    0.1513579, 0.1513599, 0.1513615, 0.1513637, 0.1513677, 0.1513668, 
    0.1513701, 0.1513365, 0.1513384, 0.1513383, 0.1513404, 0.1513419, 
    0.1513453, 0.1513507, 0.1513487, 0.1513524, 0.1513531, 0.1513475, 
    0.1513509, 0.1513398, 0.1513415, 0.1513405, 0.1513366, 0.1513491, 
    0.1513426, 0.1513546, 0.1513511, 0.1513613, 0.1513561, 0.1513662, 
    0.1513705, 0.1513747, 0.1513795, 0.1513396, 0.1513382, 0.1513407, 
    0.1513439, 0.1513471, 0.1513513, 0.1513517, 0.1513525, 0.1513545, 
    0.1513562, 0.1513527, 0.1513567, 0.1513418, 0.1513496, 0.1513377, 
    0.1513412, 0.1513438, 0.1513427, 0.1513484, 0.1513498, 0.1513552, 
    0.1513525, 0.1513694, 0.1513618, 0.1513832, 0.1513772, 0.1513378, 
    0.1513396, 0.1513459, 0.1513429, 0.1513516, 0.1513537, 0.1513555, 
    0.1513577, 0.1513579, 0.1513593, 0.1513571, 0.1513592, 0.1513513, 
    0.1513548, 0.1513452, 0.1513475, 0.1513465, 0.1513453, 0.1513489, 
    0.1513527, 0.1513529, 0.1513541, 0.1513574, 0.1513516, 0.1513702, 
    0.1513585, 0.1513416, 0.151345, 0.1513456, 0.1513442, 0.1513535, 
    0.1513501, 0.1513592, 0.1513568, 0.1513608, 0.1513588, 0.1513585, 
    0.1513559, 0.1513543, 0.1513503, 0.151347, 0.1513444, 0.151345, 
    0.1513478, 0.151353, 0.1513579, 0.1513568, 0.1513605, 0.1513509, 
    0.1513549, 0.1513533, 0.1513574, 0.1513486, 0.1513559, 0.1513467, 
    0.1513475, 0.1513501, 0.1513551, 0.1513564, 0.1513575, 0.1513568, 
    0.1513531, 0.1513526, 0.15135, 0.1513493, 0.1513474, 0.1513457, 
    0.1513472, 0.1513487, 0.1513532, 0.1513571, 0.1513616, 0.1513627, 
    0.1513677, 0.1513635, 0.1513703, 0.1513643, 0.1513747, 0.1513564, 
    0.1513643, 0.1513502, 0.1513517, 0.1513544, 0.1513608, 0.1513574, 
    0.1513614, 0.1513526, 0.1513479, 0.1513468, 0.1513446, 0.1513468, 
    0.1513467, 0.1513488, 0.1513481, 0.1513533, 0.1513505, 0.1513585, 
    0.1513614, 0.1513697, 0.1513749, 0.1513802, 0.1513826, 0.1513833, 
    0.1513836,
  0.1611694, 0.1611753, 0.1611742, 0.1611789, 0.1611763, 0.1611794, 
    0.1611706, 0.1611755, 0.1611724, 0.16117, 0.161188, 0.1611791, 0.1611977, 
    0.1611919, 0.1612066, 0.1611967, 0.1612086, 0.1612064, 0.1612133, 
    0.1612114, 0.1612201, 0.1612142, 0.1612248, 0.1612187, 0.1612196, 
    0.161214, 0.161181, 0.1611869, 0.1611806, 0.1611815, 0.1611811, 
    0.1611763, 0.1611739, 0.161169, 0.1611699, 0.1611735, 0.1611818, 
    0.1611791, 0.1611863, 0.1611861, 0.1611941, 0.1611905, 0.161204, 
    0.1612002, 0.1612114, 0.1612086, 0.1612113, 0.1612105, 0.1612113, 
    0.1612071, 0.1612089, 0.1612052, 0.1611911, 0.1611952, 0.161183, 
    0.1611755, 0.1611708, 0.1611675, 0.1611679, 0.1611688, 0.1611735, 
    0.1611781, 0.1611815, 0.1611838, 0.1611861, 0.1611927, 0.1611965, 
    0.1612048, 0.1612033, 0.1612058, 0.1612083, 0.1612124, 0.1612117, 
    0.1612135, 0.1612058, 0.1612109, 0.1612025, 0.1612048, 0.1611864, 
    0.1611798, 0.1611768, 0.1611744, 0.1611683, 0.1611725, 0.1611708, 
    0.1611748, 0.1611774, 0.1611761, 0.1611839, 0.1611808, 0.1611967, 
    0.1611899, 0.161208, 0.1612036, 0.1612091, 0.1612063, 0.161211, 
    0.1612068, 0.1612142, 0.1612158, 0.1612147, 0.161219, 0.1612065, 
    0.1612113, 0.1611761, 0.1611763, 0.1611772, 0.161173, 0.1611728, 
    0.161169, 0.1611724, 0.1611738, 0.1611775, 0.1611797, 0.1611817, 
    0.1611863, 0.1611914, 0.1611986, 0.1612039, 0.1612075, 0.1612053, 
    0.1612072, 0.1612051, 0.1612041, 0.1612151, 0.1612089, 0.1612183, 
    0.1612178, 0.1612135, 0.1612179, 0.1611764, 0.1611753, 0.1611712, 
    0.1611744, 0.1611686, 0.1611718, 0.1611736, 0.1611808, 0.1611825, 
    0.161184, 0.1611869, 0.1611907, 0.1611972, 0.1612031, 0.1612085, 
    0.1612081, 0.1612082, 0.1612094, 0.1612064, 0.1612099, 0.1612104, 
    0.1612089, 0.1612178, 0.1612152, 0.1612178, 0.1612162, 0.1611756, 
    0.1611776, 0.1611765, 0.1611785, 0.1611771, 0.1611833, 0.1611852, 
    0.1611941, 0.1611906, 0.1611964, 0.1611912, 0.1611921, 0.1611964, 
    0.1611915, 0.1612027, 0.161195, 0.1612094, 0.1612015, 0.1612099, 
    0.1612084, 0.1612109, 0.1612131, 0.1612159, 0.1612211, 0.1612199, 
    0.1612243, 0.1611806, 0.1611831, 0.1611829, 0.1611856, 0.1611876, 
    0.161192, 0.1611989, 0.1611963, 0.1612012, 0.1612021, 0.1611948, 
    0.1611992, 0.1611848, 0.1611871, 0.1611858, 0.1611807, 0.1611968, 
    0.1611885, 0.161204, 0.1611995, 0.1612128, 0.1612061, 0.1612193, 
    0.1612248, 0.1612303, 0.1612365, 0.1611845, 0.1611828, 0.1611859, 
    0.1611902, 0.1611943, 0.1611997, 0.1612003, 0.1612013, 0.161204, 
    0.1612062, 0.1612016, 0.1612068, 0.1611875, 0.1611976, 0.1611821, 
    0.1611867, 0.16119, 0.1611886, 0.161196, 0.1611978, 0.1612049, 0.1612012, 
    0.1612234, 0.1612135, 0.1612414, 0.1612335, 0.1611822, 0.1611845, 
    0.1611927, 0.1611888, 0.1612001, 0.1612029, 0.1612052, 0.1612081, 
    0.1612084, 0.1612101, 0.1612073, 0.16121, 0.1611997, 0.1612043, 
    0.1611919, 0.1611948, 0.1611935, 0.161192, 0.1611967, 0.1612016, 
    0.1612018, 0.1612034, 0.1612077, 0.1612002, 0.1612245, 0.1612092, 
    0.1611871, 0.1611916, 0.1611923, 0.1611906, 0.1612026, 0.1611982, 
    0.1612101, 0.1612069, 0.1612122, 0.1612095, 0.1612092, 0.1612058, 
    0.1612037, 0.1611984, 0.1611941, 0.1611908, 0.1611916, 0.1611953, 
    0.161202, 0.1612084, 0.161207, 0.1612118, 0.1611993, 0.1612045, 
    0.1612024, 0.1612078, 0.1611962, 0.1612057, 0.1611938, 0.1611948, 
    0.1611981, 0.1612047, 0.1612063, 0.1612079, 0.161207, 0.1612021, 
    0.1612014, 0.1611981, 0.1611971, 0.1611946, 0.1611925, 0.1611944, 
    0.1611964, 0.1612022, 0.1612074, 0.1612131, 0.1612146, 0.1612211, 
    0.1612156, 0.1612245, 0.1612168, 0.1612303, 0.1612064, 0.1612167, 
    0.1611983, 0.1612003, 0.1612038, 0.1612121, 0.1612077, 0.1612129, 
    0.1612014, 0.1611953, 0.1611939, 0.161191, 0.161194, 0.1611937, 
    0.1611965, 0.1611957, 0.1612024, 0.1611988, 0.1612091, 0.1612129, 
    0.1612238, 0.1612305, 0.1612375, 0.1612406, 0.1612415, 0.1612419,
  0.175368, 0.1753724, 0.1753715, 0.1753751, 0.1753731, 0.1753754, 0.1753689, 
    0.1753725, 0.1753702, 0.1753684, 0.175382, 0.1753753, 0.1753894, 
    0.175385, 0.1753962, 0.1753886, 0.1753978, 0.1753961, 0.1754015, 
    0.1753999, 0.1754067, 0.1754022, 0.1754104, 0.1754057, 0.1754064, 
    0.175402, 0.1753767, 0.1753811, 0.1753764, 0.175377, 0.1753768, 
    0.1753732, 0.1753713, 0.1753677, 0.1753684, 0.175371, 0.1753773, 
    0.1753752, 0.1753806, 0.1753805, 0.1753866, 0.1753839, 0.1753943, 
    0.1753913, 0.1754, 0.1753978, 0.1753999, 0.1753992, 0.1753999, 0.1753966, 
    0.175398, 0.1753952, 0.1753844, 0.1753875, 0.1753782, 0.1753725, 
    0.175369, 0.1753665, 0.1753669, 0.1753675, 0.1753711, 0.1753745, 
    0.1753771, 0.1753788, 0.1753805, 0.1753856, 0.1753885, 0.1753948, 
    0.1753937, 0.1753956, 0.1753976, 0.1754007, 0.1754002, 0.1754016, 
    0.1753956, 0.1753996, 0.1753931, 0.1753948, 0.1753807, 0.1753758, 
    0.1753735, 0.1753717, 0.1753671, 0.1753703, 0.175369, 0.175372, 
    0.1753739, 0.175373, 0.1753788, 0.1753765, 0.1753886, 0.1753834, 
    0.1753973, 0.175394, 0.1753982, 0.175396, 0.1753997, 0.1753964, 
    0.1754021, 0.1754034, 0.1754025, 0.1754059, 0.1753962, 0.1753998, 
    0.175373, 0.1753731, 0.1753738, 0.1753706, 0.1753705, 0.1753677, 
    0.1753702, 0.1753712, 0.175374, 0.1753757, 0.1753772, 0.1753807, 
    0.1753846, 0.1753901, 0.1753942, 0.1753969, 0.1753953, 0.1753967, 
    0.1753951, 0.1753943, 0.1754029, 0.175398, 0.1754054, 0.175405, 
    0.1754016, 0.175405, 0.1753732, 0.1753723, 0.1753693, 0.1753717, 
    0.1753674, 0.1753697, 0.1753711, 0.1753765, 0.1753778, 0.1753789, 
    0.1753811, 0.175384, 0.175389, 0.1753935, 0.1753977, 0.1753974, 
    0.1753975, 0.1753984, 0.1753961, 0.1753988, 0.1753992, 0.1753981, 
    0.1754049, 0.1754029, 0.175405, 0.1754037, 0.1753726, 0.1753741, 
    0.1753733, 0.1753748, 0.1753737, 0.1753784, 0.1753799, 0.1753867, 
    0.1753839, 0.1753884, 0.1753844, 0.1753851, 0.1753884, 0.1753846, 
    0.1753932, 0.1753873, 0.1753984, 0.1753923, 0.1753988, 0.1753977, 
    0.1753996, 0.1754013, 0.1754035, 0.1754075, 0.1754066, 0.17541, 
    0.1753763, 0.1753782, 0.1753781, 0.1753802, 0.1753817, 0.175385, 
    0.1753903, 0.1753883, 0.1753921, 0.1753928, 0.1753872, 0.1753906, 
    0.1753796, 0.1753813, 0.1753803, 0.1753765, 0.1753887, 0.1753824, 
    0.1753942, 0.1753907, 0.175401, 0.1753958, 0.1754061, 0.1754104, 
    0.1754148, 0.1754197, 0.1753793, 0.175378, 0.1753804, 0.1753836, 
    0.1753868, 0.1753909, 0.1753914, 0.1753922, 0.1753942, 0.1753959, 
    0.1753924, 0.1753964, 0.1753816, 0.1753893, 0.1753775, 0.175381, 
    0.1753835, 0.1753824, 0.1753881, 0.1753895, 0.1753949, 0.1753921, 
    0.1754093, 0.1754016, 0.1754236, 0.1754173, 0.1753776, 0.1753794, 
    0.1753856, 0.1753826, 0.1753912, 0.1753934, 0.1753952, 0.1753974, 
    0.1753976, 0.175399, 0.1753968, 0.1753989, 0.1753909, 0.1753945, 
    0.1753849, 0.1753872, 0.1753862, 0.175385, 0.1753886, 0.1753924, 
    0.1753926, 0.1753938, 0.1753971, 0.1753913, 0.1754102, 0.1753983, 
    0.1753813, 0.1753847, 0.1753853, 0.1753839, 0.1753931, 0.1753898, 
    0.1753989, 0.1753965, 0.1754006, 0.1753985, 0.1753982, 0.1753956, 
    0.175394, 0.1753899, 0.1753867, 0.1753841, 0.1753847, 0.1753875, 
    0.1753927, 0.1753976, 0.1753965, 0.1754003, 0.1753906, 0.1753946, 
    0.175393, 0.1753971, 0.1753883, 0.1753956, 0.1753864, 0.1753872, 
    0.1753897, 0.1753948, 0.1753961, 0.1753972, 0.1753965, 0.1753928, 
    0.1753922, 0.1753897, 0.1753889, 0.175387, 0.1753854, 0.1753869, 
    0.1753884, 0.1753928, 0.1753968, 0.1754013, 0.1754024, 0.1754075, 
    0.1754033, 0.1754102, 0.1754041, 0.1754148, 0.1753961, 0.1754041, 
    0.1753899, 0.1753914, 0.1753941, 0.1754005, 0.1753971, 0.1754011, 
    0.1753922, 0.1753876, 0.1753865, 0.1753843, 0.1753865, 0.1753863, 
    0.1753885, 0.1753878, 0.175393, 0.1753902, 0.1753982, 0.1754011, 
    0.1754096, 0.1754149, 0.1754205, 0.1754229, 0.1754237, 0.175424,
  0.1899665, 0.1899678, 0.1899675, 0.1899686, 0.189968, 0.1899687, 0.1899667, 
    0.1899678, 0.1899671, 0.1899666, 0.1899708, 0.1899687, 0.1899731, 
    0.1899717, 0.1899754, 0.1899729, 0.1899759, 0.1899754, 0.1899772, 
    0.1899767, 0.189979, 0.1899774, 0.1899803, 0.1899786, 0.1899789, 
    0.1899774, 0.1899691, 0.1899705, 0.189969, 0.1899692, 0.1899691, 
    0.189968, 0.1899675, 0.1899664, 0.1899666, 0.1899674, 0.1899693, 
    0.1899687, 0.1899703, 0.1899703, 0.1899723, 0.1899714, 0.1899748, 
    0.1899738, 0.1899767, 0.1899759, 0.1899766, 0.1899764, 0.1899766, 
    0.1899756, 0.189976, 0.1899751, 0.1899715, 0.1899725, 0.1899696, 
    0.1899678, 0.1899668, 0.189966, 0.1899661, 0.1899663, 0.1899674, 
    0.1899684, 0.1899692, 0.1899698, 0.1899703, 0.1899719, 0.1899728, 
    0.1899749, 0.1899746, 0.1899752, 0.1899759, 0.1899769, 0.1899768, 
    0.1899772, 0.1899752, 0.1899765, 0.1899744, 0.1899749, 0.1899704, 
    0.1899688, 0.1899681, 0.1899676, 0.1899662, 0.1899672, 0.1899668, 
    0.1899677, 0.1899683, 0.189968, 0.1899698, 0.1899691, 0.1899729, 
    0.1899712, 0.1899758, 0.1899747, 0.1899761, 0.1899754, 0.1899766, 
    0.1899755, 0.1899774, 0.1899778, 0.1899776, 0.1899787, 0.1899754, 
    0.1899766, 0.189968, 0.189968, 0.1899682, 0.1899673, 0.1899672, 
    0.1899664, 0.1899671, 0.1899675, 0.1899683, 0.1899688, 0.1899693, 
    0.1899704, 0.1899716, 0.1899734, 0.1899747, 0.1899756, 0.1899751, 
    0.1899756, 0.189975, 0.1899748, 0.1899777, 0.189976, 0.1899785, 
    0.1899784, 0.1899772, 0.1899784, 0.189968, 0.1899678, 0.1899669, 
    0.1899676, 0.1899663, 0.189967, 0.1899674, 0.1899691, 0.1899695, 
    0.1899698, 0.1899705, 0.1899714, 0.189973, 0.1899745, 0.1899759, 
    0.1899758, 0.1899758, 0.1899761, 0.1899754, 0.1899763, 0.1899764, 
    0.189976, 0.1899784, 0.1899777, 0.1899784, 0.189978, 0.1899679, 
    0.1899683, 0.1899681, 0.1899685, 0.1899682, 0.1899697, 0.1899701, 
    0.1899723, 0.1899714, 0.1899728, 0.1899715, 0.1899718, 0.1899728, 
    0.1899716, 0.1899744, 0.1899725, 0.1899762, 0.1899741, 0.1899763, 
    0.1899759, 0.1899766, 0.1899771, 0.1899779, 0.1899793, 0.189979, 
    0.1899802, 0.189969, 0.1899696, 0.1899696, 0.1899702, 0.1899707, 
    0.1899717, 0.1899735, 0.1899728, 0.189974, 0.1899743, 0.1899724, 
    0.1899735, 0.18997, 0.1899705, 0.1899702, 0.189969, 0.1899729, 0.1899709, 
    0.1899748, 0.1899736, 0.189977, 0.1899753, 0.1899788, 0.1899803, 
    0.1899819, 0.1899836, 0.1899699, 0.1899695, 0.1899703, 0.1899713, 
    0.1899723, 0.1899737, 0.1899738, 0.1899741, 0.1899747, 0.1899753, 
    0.1899741, 0.1899755, 0.1899706, 0.1899731, 0.1899694, 0.1899704, 
    0.1899712, 0.1899709, 0.1899727, 0.1899732, 0.189975, 0.189974, 
    0.1899799, 0.1899772, 0.1899851, 0.1899828, 0.1899694, 0.1899699, 
    0.1899719, 0.189971, 0.1899738, 0.1899745, 0.1899751, 0.1899758, 
    0.1899759, 0.1899763, 0.1899756, 0.1899763, 0.1899737, 0.1899748, 
    0.1899717, 0.1899724, 0.1899721, 0.1899717, 0.1899729, 0.1899741, 
    0.1899742, 0.1899746, 0.1899757, 0.1899738, 0.1899802, 0.1899761, 
    0.1899706, 0.1899716, 0.1899718, 0.1899714, 0.1899744, 0.1899733, 
    0.1899763, 0.1899755, 0.1899769, 0.1899762, 0.1899761, 0.1899752, 
    0.1899747, 0.1899733, 0.1899723, 0.1899715, 0.1899716, 0.1899725, 
    0.1899742, 0.1899759, 0.1899755, 0.1899768, 0.1899735, 0.1899749, 
    0.1899743, 0.1899757, 0.1899728, 0.1899752, 0.1899722, 0.1899724, 
    0.1899733, 0.1899749, 0.1899754, 0.1899758, 0.1899755, 0.1899743, 
    0.1899741, 0.1899733, 0.189973, 0.1899724, 0.1899719, 0.1899723, 
    0.1899728, 0.1899743, 0.1899756, 0.1899771, 0.1899775, 0.1899793, 
    0.1899778, 0.1899802, 0.1899781, 0.1899819, 0.1899754, 0.1899781, 
    0.1899733, 0.1899738, 0.1899747, 0.1899769, 0.1899757, 0.1899771, 
    0.1899741, 0.1899725, 0.1899722, 0.1899715, 0.1899722, 0.1899722, 
    0.1899729, 0.1899726, 0.1899743, 0.1899734, 0.1899761, 0.1899771, 
    0.18998, 0.1899819, 0.1899839, 0.1899848, 0.1899851, 0.1899852,
  0.1973253, 0.1973253, 0.1973253, 0.1973252, 0.1973253, 0.1973252, 
    0.1973253, 0.1973253, 0.1973253, 0.1973253, 0.1973252, 0.1973252, 
    0.1973251, 0.1973252, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973252, 0.1973251, 0.1973252, 0.1973252, 0.1973252, 0.1973252, 
    0.1973252, 0.1973252, 0.1973252, 0.1973252, 0.1973252, 0.1973252, 
    0.1973252, 0.1973253, 0.1973253, 0.1973253, 0.1973253, 0.1973253, 
    0.1973252, 0.1973252, 0.1973252, 0.1973252, 0.1973251, 0.1973252, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973252, 0.1973251, 
    0.1973252, 0.1973253, 0.1973253, 0.1973254, 0.1973253, 0.1973253, 
    0.1973253, 0.1973252, 0.1973252, 0.1973252, 0.1973252, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973252, 
    0.1973252, 0.1973252, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973252, 0.1973252, 0.1973252, 0.1973253, 0.1973253, 0.1973253, 
    0.1973253, 0.1973253, 0.1973252, 0.1973253, 0.1973252, 0.1973252, 
    0.1973251, 0.1973252, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973252, 0.1973252, 0.1973252, 0.1973252, 
    0.1973251, 0.1973251, 0.1973253, 0.1973253, 0.1973252, 0.1973253, 
    0.1973253, 0.1973253, 0.1973253, 0.1973253, 0.1973252, 0.1973252, 
    0.1973252, 0.1973252, 0.1973252, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973252, 0.1973251, 
    0.1973252, 0.1973252, 0.1973252, 0.1973252, 0.1973253, 0.1973253, 
    0.1973253, 0.1973253, 0.1973253, 0.1973253, 0.1973253, 0.1973252, 
    0.1973252, 0.1973252, 0.1973252, 0.1973252, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973252, 0.1973252, 0.1973252, 0.1973252, 
    0.1973253, 0.1973252, 0.1973253, 0.1973252, 0.1973252, 0.1973252, 
    0.1973252, 0.1973251, 0.1973252, 0.1973251, 0.1973252, 0.1973252, 
    0.1973251, 0.1973252, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973252, 0.1973252, 0.1973252, 
    0.1973252, 0.1973252, 0.1973252, 0.1973252, 0.1973252, 0.1973252, 
    0.1973252, 0.1973252, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973252, 0.1973252, 0.1973252, 0.1973252, 
    0.1973251, 0.1973252, 0.1973251, 0.1973251, 0.1973252, 0.1973251, 
    0.1973252, 0.1973252, 0.1973253, 0.1973254, 0.1973252, 0.1973252, 
    0.1973252, 0.1973252, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973252, 0.1973251, 
    0.1973252, 0.1973252, 0.1973252, 0.1973252, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973252, 0.1973252, 0.1973254, 0.1973253, 
    0.1973252, 0.1973252, 0.1973251, 0.1973252, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973252, 0.1973251, 0.1973251, 0.1973252, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973252, 0.1973251, 0.1973252, 0.1973252, 0.1973251, 0.1973252, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973252, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973252, 
    0.1973252, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973252, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973252, 
    0.1973252, 0.1973252, 0.1973252, 0.1973252, 0.1973252, 0.1973253, 
    0.1973251, 0.1973252, 0.1973251, 0.1973251, 0.1973251, 0.1973252, 
    0.1973251, 0.1973252, 0.1973251, 0.1973251, 0.1973251, 0.1973252, 
    0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 0.1973251, 
    0.1973251, 0.1973252, 0.1973252, 0.1973253, 0.1973254, 0.1973254, 
    0.1973254, 0.1973254,
  0.1984806, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 
    0.1984806, 0.1984805, 0.1984805, 0.1984806, 0.1984805, 0.1984805, 
    0.1984804, 0.1984805, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984803, 0.1984804, 0.1984803, 0.1984803, 
    0.1984803, 0.1984804, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 
    0.1984805, 0.1984805, 0.1984805, 0.1984806, 0.1984806, 0.1984805, 
    0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984804, 0.1984805, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984805, 0.1984804, 
    0.1984805, 0.1984805, 0.1984806, 0.1984806, 0.1984806, 0.1984806, 
    0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984806, 0.1984805, 
    0.1984806, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 
    0.1984804, 0.1984805, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984803, 
    0.1984804, 0.1984804, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 
    0.1984805, 0.1984806, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 
    0.1984805, 0.1984805, 0.1984805, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984803, 0.1984804, 0.1984804, 0.1984804, 0.1984805, 0.1984805, 
    0.1984806, 0.1984805, 0.1984806, 0.1984806, 0.1984805, 0.1984805, 
    0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 
    0.1984805, 0.1984804, 0.1984805, 0.1984804, 0.1984805, 0.1984805, 
    0.1984804, 0.1984805, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984803, 
    0.1984803, 0.1984803, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 
    0.1984805, 0.1984805, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 
    0.1984804, 0.1984805, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984803, 0.1984803, 0.1984803, 0.1984803, 0.1984805, 0.1984805, 
    0.1984805, 0.1984805, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984805, 0.1984804, 
    0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984803, 0.1984804, 0.1984803, 0.1984803, 
    0.1984805, 0.1984805, 0.1984805, 0.1984805, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984805, 0.1984804, 0.1984804, 0.1984805, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984803, 0.1984804, 0.1984805, 0.1984805, 0.1984805, 0.1984805, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984805, 
    0.1984805, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984805, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984803, 0.1984804, 0.1984803, 0.1984804, 0.1984803, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984805, 
    0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 0.1984804, 
    0.1984804, 0.1984804, 0.1984803, 0.1984803, 0.1984803, 0.1984803, 
    0.1984803, 0.1984803,
  0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 U10 =
  5.61174, 5.611793, 5.611783, 5.611824, 5.611802, 5.611828, 5.611751, 
    5.611794, 5.611767, 5.611745, 5.611903, 5.611826, 5.611987, 5.611938, 
    5.612066, 5.611979, 5.612084, 5.612064, 5.612125, 5.612108, 5.612183, 
    5.612134, 5.612223, 5.612172, 5.612179, 5.612132, 5.611843, 5.611893, 
    5.611839, 5.611847, 5.611844, 5.611802, 5.611779, 5.611737, 5.611744, 
    5.611776, 5.61185, 5.611826, 5.611889, 5.611887, 5.611956, 5.611925, 
    5.612043, 5.612009, 5.612109, 5.612083, 5.612107, 5.612101, 5.612108, 
    5.612071, 5.612086, 5.612054, 5.611931, 5.611966, 5.61186, 5.611794, 
    5.611753, 5.611722, 5.611727, 5.611734, 5.611777, 5.611817, 5.611847, 
    5.611867, 5.611887, 5.611944, 5.611977, 5.61205, 5.612037, 5.612059, 
    5.612081, 5.612117, 5.612111, 5.612127, 5.612059, 5.612104, 5.612029, 
    5.61205, 5.611888, 5.611833, 5.611805, 5.611784, 5.61173, 5.611767, 
    5.611753, 5.611788, 5.611811, 5.6118, 5.611868, 5.611841, 5.611979, 
    5.61192, 5.612079, 5.61204, 5.612088, 5.612064, 5.612105, 5.612068, 
    5.612133, 5.612146, 5.612137, 5.612174, 5.612066, 5.612107, 5.611799, 
    5.611801, 5.61181, 5.611772, 5.61177, 5.611736, 5.611766, 5.611779, 
    5.611812, 5.611831, 5.611849, 5.611889, 5.611933, 5.611995, 5.612042, 
    5.612074, 5.612055, 5.612072, 5.612052, 5.612044, 5.612141, 5.612086, 
    5.612169, 5.612164, 5.612127, 5.612165, 5.611803, 5.611792, 5.611755, 
    5.611784, 5.611732, 5.611761, 5.611777, 5.611841, 5.611856, 5.611868, 
    5.611894, 5.611927, 5.611983, 5.612034, 5.612082, 5.612079, 5.612081, 
    5.612091, 5.612064, 5.612095, 5.6121, 5.612087, 5.612164, 5.612142, 
    5.612164, 5.61215, 5.611795, 5.611813, 5.611804, 5.611821, 5.611808, 
    5.611863, 5.611879, 5.611957, 5.611926, 5.611976, 5.611931, 5.611939, 
    5.611976, 5.611934, 5.61203, 5.611963, 5.612091, 5.61202, 5.612095, 
    5.612082, 5.612104, 5.612123, 5.612148, 5.612192, 5.612182, 5.612219, 
    5.611839, 5.611861, 5.61186, 5.611883, 5.6119, 5.611938, 5.611998, 
    5.611976, 5.612017, 5.612025, 5.611963, 5.612, 5.611876, 5.611896, 
    5.611885, 5.61184, 5.61198, 5.611908, 5.612043, 5.612002, 5.612121, 
    5.612061, 5.612176, 5.612223, 5.61227, 5.612321, 5.611874, 5.611859, 
    5.611886, 5.611923, 5.611959, 5.612005, 5.61201, 5.612018, 5.612043, 
    5.612062, 5.61202, 5.612068, 5.611898, 5.611986, 5.611852, 5.611892, 
    5.611921, 5.611909, 5.611973, 5.611988, 5.612051, 5.612018, 5.612211, 
    5.612126, 5.612363, 5.612297, 5.611853, 5.611874, 5.611944, 5.611911, 
    5.612008, 5.612032, 5.612054, 5.612079, 5.612082, 5.612097, 5.612072, 
    5.612097, 5.612005, 5.612046, 5.611937, 5.611963, 5.611951, 5.611938, 
    5.611979, 5.61202, 5.612023, 5.612037, 5.612074, 5.612009, 5.612219, 
    5.612088, 5.611896, 5.611934, 5.611941, 5.611926, 5.61203, 5.611992, 
    5.612097, 5.612069, 5.612115, 5.612092, 5.612089, 5.612059, 5.61204, 
    5.611993, 5.611957, 5.611928, 5.611935, 5.611967, 5.612023, 5.612082, 
    5.612069, 5.612112, 5.612001, 5.612047, 5.612028, 5.612076, 5.611975, 
    5.612057, 5.611954, 5.611963, 5.611991, 5.612049, 5.612064, 5.612078, 
    5.61207, 5.612025, 5.612019, 5.611991, 5.611982, 5.611961, 5.611943, 
    5.611959, 5.611976, 5.612026, 5.612073, 5.612123, 5.612136, 5.612192, 
    5.612145, 5.61222, 5.612154, 5.612269, 5.612064, 5.612154, 5.611993, 
    5.61201, 5.612041, 5.612114, 5.612076, 5.612121, 5.612019, 5.611967, 
    5.611955, 5.61193, 5.611956, 5.611953, 5.611978, 5.61197, 5.612028, 
    5.611997, 5.612088, 5.612121, 5.612215, 5.612271, 5.61233, 5.612356, 
    5.612364, 5.612367 ;

 URBAN_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 URBAN_HEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 VOCFLXT =
  6.476529e-15, 6.475328e-15, 6.475556e-15, 6.474602e-15, 6.475123e-15, 
    6.474504e-15, 6.476275e-15, 6.47529e-15, 6.475913e-15, 6.476407e-15, 
    6.472782e-15, 6.474556e-15, 6.47085e-15, 6.471993e-15, 6.469094e-15, 
    6.47104e-15, 6.468699e-15, 6.469128e-15, 6.467783e-15, 6.468166e-15, 
    6.466497e-15, 6.467606e-15, 6.465597e-15, 6.466749e-15, 6.466578e-15, 
    6.467646e-15, 6.474177e-15, 6.473009e-15, 6.474252e-15, 6.474084e-15, 
    6.474154e-15, 6.47512e-15, 6.475622e-15, 6.476605e-15, 6.476422e-15, 
    6.475691e-15, 6.474008e-15, 6.474564e-15, 6.47312e-15, 6.473152e-15, 
    6.471563e-15, 6.472279e-15, 6.469595e-15, 6.470353e-15, 6.46815e-15, 
    6.468706e-15, 6.46818e-15, 6.468337e-15, 6.468178e-15, 6.468993e-15, 
    6.468645e-15, 6.469355e-15, 6.47215e-15, 6.471334e-15, 6.473779e-15, 
    6.475287e-15, 6.476236e-15, 6.476927e-15, 6.476829e-15, 6.476648e-15, 
    6.475688e-15, 6.474767e-15, 6.474073e-15, 6.473613e-15, 6.473156e-15, 
    6.471836e-15, 6.471088e-15, 6.469453e-15, 6.469729e-15, 6.469247e-15, 
    6.468761e-15, 6.46797e-15, 6.468097e-15, 6.467754e-15, 6.469246e-15, 
    6.468261e-15, 6.46989e-15, 6.469447e-15, 6.473108e-15, 6.47441e-15, 
    6.47503e-15, 6.475515e-15, 6.476756e-15, 6.475903e-15, 6.476241e-15, 
    6.475422e-15, 6.474912e-15, 6.475161e-15, 6.4736e-15, 6.474209e-15, 
    6.471044e-15, 6.472405e-15, 6.468817e-15, 6.469671e-15, 6.468611e-15, 
    6.469147e-15, 6.468234e-15, 6.469056e-15, 6.46762e-15, 6.467316e-15, 
    6.467526e-15, 6.466698e-15, 6.469103e-15, 6.468188e-15, 6.475171e-15, 
    6.475132e-15, 6.474936e-15, 6.475798e-15, 6.475846e-15, 6.476614e-15, 
    6.475924e-15, 6.475636e-15, 6.474877e-15, 6.474442e-15, 6.474024e-15, 
    6.473105e-15, 6.472093e-15, 6.470658e-15, 6.469616e-15, 6.468923e-15, 
    6.469343e-15, 6.468973e-15, 6.469389e-15, 6.469582e-15, 6.467435e-15, 
    6.468646e-15, 6.466817e-15, 6.466915e-15, 6.467749e-15, 6.466904e-15, 
    6.475102e-15, 6.475335e-15, 6.47617e-15, 6.475516e-15, 6.476697e-15, 
    6.476045e-15, 6.475677e-15, 6.474213e-15, 6.473874e-15, 6.473583e-15, 
    6.472992e-15, 6.472243e-15, 6.470935e-15, 6.469786e-15, 6.468729e-15, 
    6.468805e-15, 6.468779e-15, 6.468551e-15, 6.469126e-15, 6.468456e-15, 
    6.468351e-15, 6.468637e-15, 6.466929e-15, 6.467415e-15, 6.466917e-15, 
    6.467233e-15, 6.475257e-15, 6.474862e-15, 6.475076e-15, 6.474677e-15, 
    6.474964e-15, 6.473707e-15, 6.47333e-15, 6.471551e-15, 6.472262e-15, 
    6.471109e-15, 6.472139e-15, 6.471961e-15, 6.471104e-15, 6.472078e-15, 
    6.469864e-15, 6.471393e-15, 6.468542e-15, 6.470096e-15, 6.468447e-15, 
    6.468734e-15, 6.468251e-15, 6.467827e-15, 6.46728e-15, 6.466294e-15, 
    6.466519e-15, 6.465683e-15, 6.474265e-15, 6.473759e-15, 6.47379e-15, 
    6.473251e-15, 6.472856e-15, 6.471983e-15, 6.470601e-15, 6.471116e-15, 
    6.470156e-15, 6.469967e-15, 6.471419e-15, 6.470541e-15, 6.47341e-15, 
    6.472961e-15, 6.473218e-15, 6.474233e-15, 6.471017e-15, 6.472674e-15, 
    6.469602e-15, 6.470495e-15, 6.467889e-15, 6.469198e-15, 6.466646e-15, 
    6.465595e-15, 6.464543e-15, 6.463391e-15, 6.473468e-15, 6.473813e-15, 
    6.473182e-15, 6.472338e-15, 6.471515e-15, 6.470444e-15, 6.470326e-15, 
    6.47013e-15, 6.469604e-15, 6.469169e-15, 6.470082e-15, 6.469059e-15, 
    6.472885e-15, 6.470867e-15, 6.473956e-15, 6.473044e-15, 6.472382e-15, 
    6.472658e-15, 6.471171e-15, 6.470826e-15, 6.469431e-15, 6.470144e-15, 
    6.465867e-15, 6.467757e-15, 6.462469e-15, 6.463951e-15, 6.473937e-15, 
    6.473462e-15, 6.471835e-15, 6.472607e-15, 6.470365e-15, 6.469819e-15, 
    6.469364e-15, 6.468808e-15, 6.468737e-15, 6.468405e-15, 6.46895e-15, 
    6.468421e-15, 6.470441e-15, 6.469535e-15, 6.472004e-15, 6.47141e-15, 
    6.471679e-15, 6.471983e-15, 6.471045e-15, 6.470071e-15, 6.470027e-15, 
    6.469718e-15, 6.468891e-15, 6.470355e-15, 6.465665e-15, 6.468596e-15, 
    6.472947e-15, 6.472067e-15, 6.471913e-15, 6.472259e-15, 6.469875e-15, 
    6.470741e-15, 6.46841e-15, 6.469034e-15, 6.468006e-15, 6.468518e-15, 
    6.468595e-15, 6.469249e-15, 6.469663e-15, 6.470706e-15, 6.471549e-15, 
    6.472205e-15, 6.472051e-15, 6.471329e-15, 6.470006e-15, 6.468741e-15, 
    6.469021e-15, 6.468084e-15, 6.470527e-15, 6.469513e-15, 6.469912e-15, 
    6.468868e-15, 6.471134e-15, 6.469273e-15, 6.471619e-15, 6.471408e-15, 
    6.470758e-15, 6.46946e-15, 6.469139e-15, 6.468838e-15, 6.469019e-15, 
    6.469967e-15, 6.470114e-15, 6.470768e-15, 6.47096e-15, 6.471453e-15, 
    6.471871e-15, 6.471495e-15, 6.471104e-15, 6.469957e-15, 6.46894e-15, 
    6.467825e-15, 6.467543e-15, 6.466299e-15, 6.467342e-15, 6.465653e-15, 
    6.467136e-15, 6.464548e-15, 6.469131e-15, 6.467134e-15, 6.470721e-15, 
    6.470328e-15, 6.469641e-15, 6.468024e-15, 6.468872e-15, 6.467869e-15, 
    6.470117e-15, 6.471315e-15, 6.471597e-15, 6.47217e-15, 6.471584e-15, 
    6.47163e-15, 6.471072e-15, 6.47125e-15, 6.469919e-15, 6.470633e-15, 
    6.468603e-15, 6.467871e-15, 6.465779e-15, 6.464514e-15, 6.463194e-15, 
    6.462624e-15, 6.462448e-15, 6.462376e-15 ;

 VOLR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WA =
  4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000 ;

 WASTEHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WF =
  7.115379, 7.142106, 7.136908, 7.158462, 7.146522, 7.160593, 7.120798, 
    7.143163, 7.128882, 7.11779, 7.199838, 7.159413, 7.242086, 7.216153, 
    7.281458, 7.238037, 7.290242, 7.280219, 7.310456, 7.301785, 7.340533, 
    7.314461, 7.360707, 7.334309, 7.338427, 7.3136, 7.167549, 7.19479, 
    7.165934, 7.169813, 7.168075, 7.146764, 7.135938, 7.113349, 7.117448, 
    7.134047, 7.171558, 7.158934, 7.190815, 7.190095, 7.225708, 7.209633, 
    7.269711, 7.2526, 7.302146, 7.289659, 7.301557, 7.29795, 7.301604, 
    7.283297, 7.291135, 7.275047, 7.212638, 7.230931, 7.176474, 7.143675, 
    7.121775, 7.106256, 7.108448, 7.112626, 7.134144, 7.154434, 7.169705, 
    7.179916, 7.189991, 7.220514, 7.236746, 7.273168, 7.266597, 7.277741, 
    7.288418, 7.306354, 7.303401, 7.311308, 7.277456, 7.299936, 7.262854, 
    7.27298, 7.192679, 7.162341, 7.14933, 7.137905, 7.110133, 7.1293, 
    7.121738, 7.139748, 7.151204, 7.145538, 7.180195, 7.166768, 7.237709, 
    7.207084, 7.287172, 7.267946, 7.291788, 7.279617, 7.300477, 7.281702, 
    7.314258, 7.321355, 7.316504, 7.335174, 7.280661, 7.301552, 7.145378, 
    7.146301, 7.15061, 7.131682, 7.130528, 7.113235, 7.128625, 7.135183, 
    7.151873, 7.161659, 7.170915, 7.191298, 7.214109, 7.246118, 7.269191, 
    7.284687, 7.275186, 7.283573, 7.274195, 7.269805, 7.318692, 7.291205, 
    7.332486, 7.330199, 7.311495, 7.330457, 7.14695, 7.141635, 7.123191, 
    7.137622, 7.111354, 7.126042, 7.134495, 7.167037, 7.174141, 7.180717, 
    7.193731, 7.210455, 7.239863, 7.265535, 7.289042, 7.287318, 7.287925, 
    7.293178, 7.280164, 7.295317, 7.297857, 7.291208, 7.329892, 7.318825, 
    7.33015, 7.322944, 7.143364, 7.152313, 7.147475, 7.156562, 7.150158, 
    7.178339, 7.186778, 7.226385, 7.210123, 7.236033, 7.212755, 7.216873, 
    7.236857, 7.214015, 7.264108, 7.230097, 7.293382, 7.25929, 7.295522, 
    7.28894, 7.299845, 7.309616, 7.321933, 7.344687, 7.339416, 7.358484, 
    7.165523, 7.176973, 7.175974, 7.187978, 7.196864, 7.216166, 7.247198, 
    7.235519, 7.256981, 7.261292, 7.228697, 7.248687, 7.184652, 7.194957, 
    7.188828, 7.16642, 7.238195, 7.201283, 7.269571, 7.249489, 7.308221, 
    7.278956, 7.336513, 7.361199, 7.384537, 7.411828, 7.183239, 7.175451, 
    7.18941, 7.20874, 7.226741, 7.250711, 7.253172, 7.257668, 7.269336, 
    7.279153, 7.259081, 7.281616, 7.197329, 7.241411, 7.172499, 7.193182, 
    7.207604, 7.201284, 7.234188, 7.241957, 7.273591, 7.25723, 7.355092, 
    7.311668, 7.432692, 7.398712, 7.172729, 7.183217, 7.2198, 7.202377, 
    7.252319, 7.264649, 7.274693, 7.287533, 7.288928, 7.296546, 7.284064, 
    7.296056, 7.250762, 7.270977, 7.215623, 7.229059, 7.222879, 7.216098, 
    7.237043, 7.259394, 7.259888, 7.267064, 7.287288, 7.252522, 7.360681, 
    7.29371, 7.194667, 7.214907, 7.217821, 7.20997, 7.263412, 7.244009, 
    7.296362, 7.282187, 7.305428, 7.293871, 7.292171, 7.277354, 7.268137, 
    7.244895, 7.226032, 7.21111, 7.214579, 7.230978, 7.260767, 7.289047, 
    7.282843, 7.30366, 7.248688, 7.271691, 7.262788, 7.286022, 7.235206, 
    7.278413, 7.224188, 7.228933, 7.243625, 7.273242, 7.279831, 7.286843, 
    7.282519, 7.261527, 7.2581, 7.243271, 7.239174, 7.227901, 7.218572, 
    7.227091, 7.236044, 7.261542, 7.284573, 7.309752, 7.315932, 7.345417, 
    7.321386, 7.361053, 7.327286, 7.38583, 7.280947, 7.326325, 7.244299, 
    7.253105, 7.269037, 7.305716, 7.285913, 7.309084, 7.257967, 7.231537, 
    7.22473, 7.212013, 7.225021, 7.223964, 7.236426, 7.23242, 7.262391, 
    7.246281, 7.292124, 7.308905, 7.356478, 7.385749, 7.415662, 7.428889, 
    7.43292, 7.434605 ;

 WIND =
  5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 5.566932, 
    5.566932, 5.566932 ;

 WOODC =
  0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 0.03074504, 
    0.03074504, 0.03074504 ;

 WOODC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOODC_LOSS =
  1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 1.94984e-11, 
    1.94984e-11, 1.94984e-11, 1.94984e-11 ;

 WOOD_HARVESTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOOD_HARVESTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WTGQ =
  0.0002000786, 0.0002000359, 0.000200044, 0.0002000104, 0.0002000287, 
    0.000200007, 0.0002000696, 0.0002000345, 0.0002000567, 0.0002000743, 
    0.0001999472, 0.0002000089, 0.0001998812, 0.0001999203, 0.0001998217, 
    0.0001998877, 0.0001998083, 0.0001998229, 0.0001997774, 0.0001997903, 
    0.0001997338, 0.0001997714, 0.0001997035, 0.0001997424, 0.0001997366, 
    0.0001997727, 0.0001999957, 0.000199955, 0.0001999983, 0.0001999924, 
    0.0001999949, 0.0002000286, 0.0002000462, 0.0002000815, 0.0002000749, 
    0.0002000487, 0.0001999898, 0.0002000092, 0.0001999591, 0.0001999602, 
    0.0001999056, 0.0001999302, 0.0001998387, 0.0001998644, 0.0001997898, 
    0.0001998086, 0.0001997908, 0.0001997961, 0.0001997907, 0.0001998183, 
    0.0001998065, 0.0001998306, 0.0001999257, 0.0001998978, 0.0001999818, 
    0.0002000344, 0.0002000682, 0.0002000931, 0.0002000895, 0.0002000829, 
    0.0002000486, 0.0002000163, 0.0001999921, 0.0001999761, 0.0001999604, 
    0.0001999148, 0.0001998894, 0.0001998339, 0.0001998433, 0.0001998269, 
    0.0001998104, 0.0001997837, 0.000199788, 0.0001997764, 0.0001998269, 
    0.0001997935, 0.0001998488, 0.0001998337, 0.0001999584, 0.0002000038, 
    0.0002000253, 0.0002000425, 0.0002000869, 0.0002000563, 0.0002000683, 
    0.0002000393, 0.0002000213, 0.0002000301, 0.0001999757, 0.0001999968, 
    0.0001998879, 0.0001999345, 0.0001998124, 0.0001998413, 0.0001998053, 
    0.0001998236, 0.0001997926, 0.0001998205, 0.0001997719, 0.0001997616, 
    0.0001997686, 0.0001997407, 0.0001998221, 0.000199791, 0.0002000305, 
    0.000200029, 0.0002000222, 0.0002000525, 0.0002000542, 0.0002000818, 
    0.000200057, 0.0002000468, 0.0002000201, 0.0002000049, 0.0001999904, 
    0.0001999586, 0.0001999237, 0.0001998748, 0.0001998394, 0.0001998159, 
    0.0001998302, 0.0001998176, 0.0001998318, 0.0001998383, 0.0001997656, 
    0.0001998065, 0.0001997447, 0.0001997481, 0.0001997762, 0.0001997477, 
    0.000200028, 0.0002000362, 0.0002000658, 0.0002000426, 0.0002000848, 
    0.0002000613, 0.0002000482, 0.0001999969, 0.0001999852, 0.0001999751, 
    0.0001999547, 0.0001999289, 0.0001998842, 0.0001998452, 0.0001998094, 
    0.000199812, 0.0001998111, 0.0001998033, 0.0001998228, 0.0001998001, 
    0.0001997965, 0.0001998063, 0.0001997485, 0.000199765, 0.0001997481, 
    0.0001997588, 0.0002000335, 0.0002000196, 0.0002000271, 0.0002000131, 
    0.0002000232, 0.0001999793, 0.0001999663, 0.0001999052, 0.0001999296, 
    0.0001998901, 0.0001999254, 0.0001999192, 0.0001998898, 0.0001999233, 
    0.0001998478, 0.0001998998, 0.000199803, 0.0001998556, 0.0001997998, 
    0.0001998096, 0.0001997932, 0.0001997788, 0.0001997604, 0.000199727, 
    0.0001997347, 0.0001997065, 0.0001999988, 0.0001999812, 0.0001999823, 
    0.0001999636, 0.00019995, 0.00019992, 0.0001998729, 0.0001998904, 
    0.0001998577, 0.0001998513, 0.0001999008, 0.0001998708, 0.0001999691, 
    0.0001999535, 0.0001999625, 0.0001999976, 0.000199887, 0.0001999437, 
    0.0001998389, 0.0001998693, 0.0001997809, 0.0001998252, 0.0001997389, 
    0.0001997034, 0.000199668, 0.0001996291, 0.0001999711, 0.0001999831, 
    0.0001999613, 0.0001999321, 0.000199904, 0.0001998675, 0.0001998635, 
    0.0001998568, 0.000199839, 0.0001998243, 0.0001998552, 0.0001998206, 
    0.0001999508, 0.0001998819, 0.000199988, 0.0001999564, 0.0001999337, 
    0.0001999432, 0.0001998923, 0.0001998806, 0.0001998331, 0.0001998573, 
    0.0001997126, 0.0001997764, 0.0001995981, 0.000199648, 0.0001999874, 
    0.0001999709, 0.0001999149, 0.0001999414, 0.0001998648, 0.0001998463, 
    0.0001998309, 0.000199812, 0.0001998096, 0.0001997984, 0.0001998169, 
    0.0001997989, 0.0001998674, 0.0001998367, 0.0001999207, 0.0001999004, 
    0.0001999096, 0.00019992, 0.000199888, 0.0001998548, 0.0001998534, 
    0.0001998429, 0.0001998146, 0.0001998645, 0.0001997056, 0.0001998047, 
    0.0001999531, 0.0001999228, 0.0001999176, 0.0001999295, 0.0001998482, 
    0.0001998776, 0.0001997986, 0.0001998197, 0.0001997849, 0.0001998022, 
    0.0001998048, 0.000199827, 0.000199841, 0.0001998764, 0.0001999051, 
    0.0001999277, 0.0001999224, 0.0001998976, 0.0001998526, 0.0001998097, 
    0.0001998192, 0.0001997875, 0.0001998704, 0.0001998359, 0.0001998495, 
    0.0001998141, 0.000199891, 0.0001998276, 0.0001999076, 0.0001999004, 
    0.0001998782, 0.000199834, 0.0001998233, 0.000199813, 0.0001998192, 
    0.0001998513, 0.0001998563, 0.0001998786, 0.0001998851, 0.0001999019, 
    0.0001999162, 0.0001999033, 0.00019989, 0.000199851, 0.0001998165, 
    0.0001997787, 0.0001997692, 0.0001997271, 0.0001997624, 0.0001997052, 
    0.0001997552, 0.000199668, 0.0001998229, 0.0001997553, 0.000199877, 
    0.0001998636, 0.0001998402, 0.0001997854, 0.0001998142, 0.0001997802, 
    0.0001998564, 0.0001998971, 0.0001999068, 0.0001999264, 0.0001999064, 
    0.000199908, 0.0001998889, 0.000199895, 0.0001998497, 0.000199874, 
    0.0001998051, 0.0001997803, 0.0001997097, 0.000199667, 0.0001996226, 
    0.0001996034, 0.0001995975, 0.000199595 ;

 W_SCALAR =
  0.6252279, 0.6268897, 0.6265668, 0.627906, 0.6271632, 0.62804, 0.6255649, 
    0.6269557, 0.6260679, 0.6253775, 0.6305014, 0.6279657, 0.6331295, 
    0.6315162, 0.6355648, 0.6328787, 0.6361057, 0.6354872, 0.6373473, 
    0.6368147, 0.6391912, 0.637593, 0.6404209, 0.6388096, 0.6390619, 
    0.6375403, 0.6284762, 0.6301861, 0.6283749, 0.6286188, 0.6285093, 
    0.6271786, 0.6265076, 0.6251007, 0.6253562, 0.6263894, 0.6287286, 
    0.6279349, 0.6299339, 0.6298888, 0.632111, 0.6311095, 0.6348386, 
    0.6337798, 0.6368369, 0.6360688, 0.6368009, 0.6365789, 0.6368037, 
    0.635677, 0.6361599, 0.635168, 0.6312972, 0.632436, 0.6290365, 0.6269884, 
    0.625626, 0.6246584, 0.6247953, 0.6250561, 0.6263955, 0.6276534, 
    0.6286113, 0.6292517, 0.6298823, 0.6317899, 0.632798, 0.6350527, 
    0.6346459, 0.6353348, 0.6359923, 0.6370957, 0.6369141, 0.6374001, 
    0.6353166, 0.6367017, 0.6344143, 0.6350403, 0.6300543, 0.628149, 
    0.6273388, 0.6266288, 0.6249005, 0.6260943, 0.6256238, 0.6267428, 
    0.6274533, 0.6271019, 0.6292692, 0.628427, 0.6328577, 0.6309511, 
    0.6359157, 0.6347294, 0.6361998, 0.6354497, 0.6367348, 0.6355783, 
    0.6375808, 0.6380165, 0.6377188, 0.6388618, 0.6355141, 0.6368009, 
    0.6270921, 0.6271494, 0.6274164, 0.6262425, 0.6261706, 0.6250937, 
    0.6260519, 0.6264598, 0.6274945, 0.6281062, 0.6286874, 0.6299645, 
    0.6313893, 0.633379, 0.6348064, 0.6357623, 0.6351762, 0.6356937, 
    0.6351152, 0.6348439, 0.6378533, 0.6361645, 0.6386974, 0.6385574, 
    0.6374117, 0.6385732, 0.6271897, 0.6268598, 0.625714, 0.6266108, 
    0.6249764, 0.6258916, 0.6264175, 0.6284448, 0.6288896, 0.6293021, 
    0.6301165, 0.6311608, 0.6329908, 0.6345809, 0.6360306, 0.6359244, 
    0.6359618, 0.6362855, 0.6354836, 0.6364171, 0.6365737, 0.6361642, 
    0.6385387, 0.6378608, 0.6385545, 0.6381131, 0.626967, 0.627522, 
    0.6272221, 0.6277859, 0.6273888, 0.629154, 0.6296828, 0.6321541, 
    0.6311403, 0.6327532, 0.6313041, 0.6315611, 0.6328061, 0.6313825, 
    0.6344934, 0.6323853, 0.6362981, 0.6341962, 0.6364297, 0.6360243, 
    0.6366953, 0.6372961, 0.6380513, 0.6394438, 0.6391215, 0.640285, 
    0.6283488, 0.6290679, 0.6290045, 0.6297566, 0.6303125, 0.6315166, 
    0.6334455, 0.6327204, 0.6340511, 0.6343181, 0.6322963, 0.6335381, 
    0.6295488, 0.6301943, 0.62981, 0.6284056, 0.6328877, 0.6305895, 0.63483, 
    0.6335874, 0.6372105, 0.6354101, 0.638944, 0.6404519, 0.6418688, 
    0.6435232, 0.6294601, 0.6289717, 0.629846, 0.6310548, 0.6321751, 
    0.6336632, 0.6338153, 0.6340939, 0.634815, 0.6354211, 0.634182, 0.635573, 
    0.6303442, 0.6330869, 0.6287871, 0.6300835, 0.6309835, 0.6305887, 
    0.6326375, 0.6331199, 0.6350786, 0.6340664, 0.64008, 0.6374231, 
    0.6447808, 0.6427293, 0.628801, 0.6294584, 0.6317437, 0.6306568, 
    0.6337624, 0.6345257, 0.6351458, 0.6359382, 0.6360236, 0.6364929, 
    0.6357239, 0.6364625, 0.6336663, 0.6349167, 0.6314825, 0.6323193, 
    0.6319344, 0.6315121, 0.6328149, 0.6342016, 0.634231, 0.6346754, 
    0.635927, 0.6337749, 0.6404229, 0.6363218, 0.6301748, 0.6314395, 
    0.6316199, 0.6311302, 0.6344492, 0.6332476, 0.6364814, 0.6356083, 
    0.6370386, 0.636328, 0.6362235, 0.6353102, 0.6347412, 0.6333028, 
    0.6321312, 0.6312012, 0.6314175, 0.6324388, 0.6342863, 0.6360315, 
    0.6356494, 0.6369299, 0.6335375, 0.6349612, 0.6344112, 0.6358448, 
    0.6327012, 0.6353792, 0.6320158, 0.632311, 0.6332238, 0.6350579, 
    0.635463, 0.6358957, 0.6356287, 0.6343331, 0.6341207, 0.6332015, 
    0.6329477, 0.6322467, 0.6316662, 0.6321967, 0.6327536, 0.6343336, 
    0.6357559, 0.6373047, 0.6376833, 0.6394903, 0.6380198, 0.6404457, 
    0.6383839, 0.6419505, 0.6355339, 0.6383228, 0.6332653, 0.6338111, 
    0.6347979, 0.6370578, 0.6358381, 0.6372644, 0.6341124, 0.6324741, 
    0.6320497, 0.6312578, 0.6320677, 0.6320019, 0.6327766, 0.6325276, 
    0.6343861, 0.6333881, 0.6362209, 0.6372531, 0.6401631, 0.6419437, 
    0.6437532, 0.6445512, 0.644794, 0.6448955,
  0.5466421, 0.5486842, 0.5482873, 0.5499333, 0.5490203, 0.5500979, 
    0.5470562, 0.5487653, 0.5476744, 0.5468259, 0.5531237, 0.5500066, 
    0.5563551, 0.5543713, 0.5593501, 0.5560466, 0.5600154, 0.5592547, 
    0.5615429, 0.5608876, 0.5638116, 0.5618452, 0.565325, 0.5633421, 
    0.5636525, 0.5617803, 0.5506341, 0.552736, 0.5505096, 0.5508094, 
    0.5506749, 0.5490392, 0.5482147, 0.5464858, 0.5467998, 0.5480694, 
    0.5509443, 0.5499687, 0.552426, 0.5523705, 0.5551025, 0.5538712, 
    0.558457, 0.5571547, 0.560915, 0.5599701, 0.5608706, 0.5605976, 
    0.5608742, 0.5594882, 0.5600822, 0.558862, 0.5541019, 0.5555023, 
    0.5513228, 0.5488056, 0.5471312, 0.5459424, 0.5461105, 0.546431, 
    0.5480768, 0.5496228, 0.5508001, 0.5515873, 0.5523625, 0.5547078, 
    0.5559474, 0.5587203, 0.55822, 0.5590673, 0.5598761, 0.5612334, 
    0.5610101, 0.5616078, 0.5590448, 0.5607487, 0.557935, 0.558705, 0.552574, 
    0.5502319, 0.5492362, 0.5483637, 0.5462398, 0.5477068, 0.5471286, 
    0.5485036, 0.549377, 0.5489451, 0.5516088, 0.5505736, 0.5560209, 
    0.5536765, 0.5597818, 0.5583227, 0.5601313, 0.5592086, 0.5607893, 
    0.5593668, 0.5618302, 0.5623662, 0.562, 0.5634063, 0.5592878, 0.5608708, 
    0.548933, 0.5490034, 0.5493315, 0.5478889, 0.5478005, 0.5464773, 
    0.5476547, 0.548156, 0.5494275, 0.5501794, 0.5508938, 0.5524635, 
    0.5542153, 0.5566618, 0.5584173, 0.5595931, 0.5588722, 0.5595087, 
    0.5587971, 0.5584635, 0.5621655, 0.5600878, 0.5632041, 0.5630318, 
    0.5616221, 0.5630512, 0.5490529, 0.5486475, 0.5472394, 0.5483415, 
    0.5463331, 0.5474576, 0.548104, 0.5505955, 0.5511423, 0.5516494, 
    0.5526503, 0.5539343, 0.5561845, 0.55814, 0.5599231, 0.5597925, 
    0.5598385, 0.5602367, 0.5592502, 0.5603986, 0.5605913, 0.5600874, 
    0.5630087, 0.5621746, 0.5630282, 0.5624851, 0.5487792, 0.5494613, 
    0.5490928, 0.5497857, 0.5492976, 0.5514672, 0.5521172, 0.5551556, 
    0.5539091, 0.5558923, 0.5541105, 0.5544264, 0.5559573, 0.5542068, 
    0.5580323, 0.5554399, 0.5602521, 0.5576669, 0.5604141, 0.5599154, 
    0.5607408, 0.5614799, 0.5624091, 0.5641225, 0.5637258, 0.5651577, 
    0.5504776, 0.5513614, 0.5512835, 0.5522079, 0.5528914, 0.5543717, 
    0.5567436, 0.555852, 0.5574883, 0.5578167, 0.5553305, 0.5568575, 
    0.5519527, 0.5527461, 0.5522736, 0.5505474, 0.5560577, 0.5532319, 
    0.5584463, 0.556918, 0.5613745, 0.5591598, 0.5635075, 0.5653632, 
    0.5671071, 0.5691437, 0.5518435, 0.5512431, 0.5523179, 0.553804, 
    0.5551814, 0.5570113, 0.5571983, 0.557541, 0.5584279, 0.5591734, 
    0.5576494, 0.5593603, 0.5529304, 0.5563027, 0.5510162, 0.5526099, 
    0.5537164, 0.5532309, 0.55575, 0.5563433, 0.5587521, 0.5575072, 
    0.5649055, 0.5616361, 0.5706921, 0.5681664, 0.5510334, 0.5518414, 
    0.554651, 0.5533147, 0.5571333, 0.5580721, 0.5588348, 0.5598095, 
    0.5599146, 0.5604918, 0.5595459, 0.5604544, 0.5570152, 0.5585529, 
    0.5543299, 0.5553587, 0.5548854, 0.5543662, 0.5559682, 0.5576735, 
    0.5577096, 0.5582561, 0.5597957, 0.5571488, 0.5653275, 0.5602815, 
    0.552722, 0.554277, 0.5544987, 0.5538967, 0.557978, 0.5565003, 0.5604777, 
    0.5594036, 0.5611631, 0.560289, 0.5601604, 0.559037, 0.5583372, 
    0.5565681, 0.5551274, 0.5539839, 0.5542499, 0.5555056, 0.5577776, 
    0.5599242, 0.5594543, 0.5610294, 0.5568568, 0.5586078, 0.5579312, 
    0.5596946, 0.5558283, 0.5591219, 0.5549856, 0.5553486, 0.5564709, 
    0.5587266, 0.5592249, 0.5597572, 0.5594288, 0.5578353, 0.557574, 
    0.5564436, 0.5561315, 0.5552695, 0.5545557, 0.555208, 0.5558928, 
    0.5578358, 0.5595852, 0.5614905, 0.5619563, 0.5641798, 0.5623703, 
    0.5653555, 0.5628183, 0.5672078, 0.5593122, 0.5627432, 0.5565219, 
    0.5571932, 0.5584068, 0.5611869, 0.5596863, 0.5614409, 0.5575637, 
    0.5555491, 0.5550272, 0.5540535, 0.5550494, 0.5549684, 0.555921, 
    0.5556149, 0.5579003, 0.556673, 0.5601572, 0.561427, 0.5650077, 
    0.5671993, 0.5694268, 0.5704094, 0.5707083, 0.5708333,
  0.5141742, 0.516424, 0.5159867, 0.5178004, 0.5167944, 0.5179818, 0.5146304, 
    0.5165133, 0.5153114, 0.5143767, 0.5213172, 0.5178813, 0.5248808, 
    0.5226929, 0.5281852, 0.5245405, 0.5289195, 0.5280799, 0.5306055, 
    0.5298822, 0.5331104, 0.5309392, 0.5347818, 0.5325919, 0.5329347, 
    0.5308676, 0.5185728, 0.5208897, 0.5184355, 0.518766, 0.5186177, 
    0.5168152, 0.5159066, 0.514002, 0.5143479, 0.5157466, 0.5189146, 
    0.5178395, 0.5205479, 0.5204868, 0.5234993, 0.5221415, 0.5271997, 
    0.5257629, 0.5299124, 0.5288695, 0.5298634, 0.5295621, 0.5298674, 
    0.5283377, 0.5289932, 0.5276467, 0.5223958, 0.5239401, 0.5193319, 
    0.5165578, 0.514713, 0.5134035, 0.5135887, 0.5139416, 0.5157548, 
    0.5174582, 0.5187557, 0.5196234, 0.520478, 0.523064, 0.5244311, 
    0.5274902, 0.5269382, 0.5278731, 0.5287657, 0.5302638, 0.5300173, 
    0.5306772, 0.5278483, 0.5297288, 0.5266237, 0.5274734, 0.5207111, 
    0.5181295, 0.5170323, 0.5160708, 0.5137311, 0.5153471, 0.5147101, 
    0.516225, 0.5171873, 0.5167114, 0.5196471, 0.5185062, 0.5245121, 
    0.5219267, 0.5286616, 0.5270515, 0.5290474, 0.528029, 0.5297737, 
    0.5282035, 0.5309227, 0.5315145, 0.53111, 0.5326628, 0.5281165, 
    0.5298635, 0.5166981, 0.5167757, 0.5171373, 0.5155477, 0.5154504, 
    0.5139926, 0.5152897, 0.515842, 0.517243, 0.5180716, 0.518859, 0.5205894, 
    0.5225208, 0.5252191, 0.5271559, 0.5284534, 0.5276578, 0.5283602, 
    0.527575, 0.5272069, 0.5312928, 0.5289993, 0.5324395, 0.5322493, 
    0.5306929, 0.5322707, 0.5168302, 0.5163835, 0.5148322, 0.5160463, 
    0.5138338, 0.5150726, 0.5157847, 0.5185302, 0.5191329, 0.5196919, 
    0.5207953, 0.522211, 0.5246926, 0.5268499, 0.5288176, 0.5286734, 
    0.5287242, 0.5291637, 0.528075, 0.5293424, 0.529555, 0.528999, 0.5322238, 
    0.5313029, 0.5322452, 0.5316457, 0.5165287, 0.5172803, 0.5168742, 
    0.5176378, 0.5170999, 0.5194911, 0.5202076, 0.5235578, 0.5221831, 
    0.5243703, 0.5224053, 0.5227537, 0.524442, 0.5225115, 0.5267311, 
    0.5238714, 0.5291808, 0.5263279, 0.5293595, 0.5288091, 0.5297201, 
    0.5305359, 0.5315617, 0.5334537, 0.5330157, 0.5345969, 0.5184003, 
    0.5193745, 0.5192885, 0.5203077, 0.5210611, 0.5226933, 0.5253093, 
    0.5243258, 0.526131, 0.5264933, 0.5237507, 0.525435, 0.5200261, 
    0.5209009, 0.52038, 0.5184772, 0.5245528, 0.5214365, 0.5271879, 
    0.5255018, 0.5304196, 0.5279752, 0.5327746, 0.534824, 0.5367505, 
    0.5390009, 0.5199059, 0.5192441, 0.5204288, 0.5220673, 0.5235863, 
    0.5256047, 0.525811, 0.526189, 0.5271676, 0.5279903, 0.5263087, 
    0.5281964, 0.5211041, 0.524823, 0.518994, 0.5207507, 0.5219707, 
    0.5214354, 0.5242134, 0.5248678, 0.5275254, 0.5261518, 0.5343184, 
    0.5307084, 0.5407125, 0.5379209, 0.5190129, 0.5199035, 0.5230013, 
    0.5215278, 0.5257393, 0.5267751, 0.5276166, 0.5286922, 0.5288082, 
    0.5294452, 0.5284013, 0.5294039, 0.525609, 0.5273055, 0.5226472, 
    0.5237818, 0.5232599, 0.5226873, 0.524454, 0.5263352, 0.5263751, 
    0.5269781, 0.5286769, 0.5257564, 0.5347845, 0.5292131, 0.5208744, 
    0.5225889, 0.5228334, 0.5221695, 0.5266712, 0.525041, 0.5294297, 
    0.5282443, 0.5301862, 0.5292214, 0.5290794, 0.5278397, 0.5270675, 
    0.5251158, 0.5235267, 0.5222657, 0.522559, 0.5239439, 0.5264502, 
    0.5288188, 0.5283002, 0.5300387, 0.5254341, 0.527366, 0.5266196, 
    0.5285654, 0.5242998, 0.5279334, 0.5233703, 0.5237706, 0.5250086, 
    0.5274972, 0.5280471, 0.5286345, 0.528272, 0.5265137, 0.5262254, 
    0.5249785, 0.5246342, 0.5236834, 0.5228962, 0.5236155, 0.5243708, 
    0.5265144, 0.5284447, 0.5305476, 0.5310619, 0.5335169, 0.5315189, 
    0.5348155, 0.5320136, 0.5368617, 0.5281434, 0.5319306, 0.5250648, 
    0.5258053, 0.5271443, 0.5302124, 0.5285562, 0.5304929, 0.5262141, 
    0.5239918, 0.5234162, 0.5223424, 0.5234407, 0.5233514, 0.524402, 
    0.5240644, 0.5265855, 0.5252315, 0.529076, 0.5304776, 0.5344313, 
    0.5368523, 0.5393139, 0.5404, 0.5407304, 0.5408686,
  0.507081, 0.5094715, 0.5090068, 0.5109347, 0.5098652, 0.5111276, 0.5075656, 
    0.5095665, 0.5082892, 0.507296, 0.5146751, 0.5110207, 0.5184683, 
    0.5161391, 0.5219885, 0.518106, 0.5227711, 0.5218763, 0.5245685, 
    0.5237973, 0.5272403, 0.5249244, 0.529024, 0.5266871, 0.5270529, 
    0.524848, 0.5117559, 0.5142202, 0.51161, 0.5119615, 0.5118037, 0.5098874, 
    0.5089217, 0.506898, 0.5072654, 0.5087516, 0.5121195, 0.5109762, 
    0.5138567, 0.5137916, 0.5169975, 0.5155522, 0.5209383, 0.5194078, 
    0.5238295, 0.5227178, 0.5237773, 0.523456, 0.5237815, 0.5221509, 
    0.5228496, 0.5214146, 0.5158229, 0.5174668, 0.5125632, 0.5096136, 
    0.5076534, 0.5062622, 0.5064589, 0.5068339, 0.5087603, 0.5105709, 
    0.5119505, 0.5128732, 0.5137823, 0.516534, 0.5179895, 0.5212479, 
    0.5206597, 0.5216559, 0.5226071, 0.5242043, 0.5239413, 0.524645, 
    0.5216295, 0.5236338, 0.5203248, 0.52123, 0.5140303, 0.5112846, 
    0.5101181, 0.5090961, 0.5066102, 0.5083271, 0.5076503, 0.5092601, 
    0.5102829, 0.509777, 0.5128984, 0.5116851, 0.5180758, 0.5153237, 
    0.5224962, 0.5207804, 0.5229074, 0.5218221, 0.5236816, 0.5220081, 
    0.5249068, 0.5255378, 0.5251066, 0.5267628, 0.5219153, 0.5237774, 
    0.5097629, 0.5098454, 0.5102297, 0.5085402, 0.5084368, 0.506888, 
    0.5082661, 0.5088529, 0.5103421, 0.511223, 0.5120603, 0.5139008, 
    0.5159559, 0.5188286, 0.5208917, 0.5222743, 0.5214265, 0.522175, 
    0.5213383, 0.520946, 0.5253015, 0.5228562, 0.5265246, 0.5263216, 
    0.5246617, 0.5263445, 0.5099033, 0.5094285, 0.50778, 0.5090701, 
    0.5067193, 0.5080354, 0.508792, 0.5117106, 0.5123515, 0.5129461, 
    0.5141199, 0.5156262, 0.5182679, 0.5205656, 0.5226625, 0.5225088, 
    0.5225629, 0.5230314, 0.5218711, 0.5232218, 0.5234486, 0.5228558, 
    0.5262945, 0.5253122, 0.5263174, 0.5256778, 0.5095828, 0.5103817, 
    0.50995, 0.5107618, 0.51019, 0.5127325, 0.5134947, 0.5170597, 0.5155966, 
    0.5179248, 0.515833, 0.5162038, 0.5180011, 0.515946, 0.5204391, 
    0.5173936, 0.5230495, 0.5200096, 0.52324, 0.5226534, 0.5236245, 
    0.5244943, 0.5255883, 0.5276066, 0.5271392, 0.5288267, 0.5115725, 
    0.5126085, 0.5125171, 0.5136011, 0.5144026, 0.5161396, 0.5189247, 
    0.5178775, 0.5197998, 0.5201857, 0.517265, 0.5190586, 0.5133016, 
    0.5142322, 0.513678, 0.5116543, 0.518119, 0.514802, 0.5209258, 0.5191297, 
    0.5243704, 0.5217647, 0.526882, 0.5290689, 0.5311258, 0.5335297, 
    0.5131736, 0.5124698, 0.5137299, 0.5154733, 0.5170901, 0.5192393, 
    0.5194591, 0.5198616, 0.5209042, 0.5217807, 0.5199891, 0.5220004, 
    0.5144483, 0.5184068, 0.5122038, 0.5140724, 0.5153704, 0.5148009, 
    0.5177577, 0.5184545, 0.5212854, 0.519822, 0.5285294, 0.5246783, 
    0.5353589, 0.5323759, 0.5122239, 0.5131711, 0.5164673, 0.5148991, 
    0.5193827, 0.5204859, 0.5213826, 0.5225288, 0.5226524, 0.5233315, 
    0.5222188, 0.5232875, 0.5192438, 0.5210511, 0.5160905, 0.5172982, 
    0.5167426, 0.5161331, 0.5180139, 0.5200174, 0.5200599, 0.5207022, 
    0.5225126, 0.5194008, 0.5290268, 0.523084, 0.514204, 0.5160284, 
    0.5162886, 0.515582, 0.5203753, 0.5186389, 0.5233149, 0.5220514, 
    0.5241215, 0.5230929, 0.5229416, 0.5216202, 0.5207976, 0.5187186, 
    0.5170266, 0.5156845, 0.5159966, 0.5174708, 0.5201398, 0.5226638, 
    0.522111, 0.5239642, 0.5190576, 0.5211156, 0.5203204, 0.5223936, 
    0.5178497, 0.5217201, 0.5168601, 0.5172863, 0.5186045, 0.5212553, 
    0.5218413, 0.5224674, 0.522081, 0.5202075, 0.5199004, 0.5185723, 
    0.5182058, 0.5171935, 0.5163555, 0.5171213, 0.5179254, 0.5202082, 
    0.522265, 0.5245068, 0.5250552, 0.5276741, 0.5255426, 0.5290599, 
    0.5260702, 0.5312445, 0.5219439, 0.5259817, 0.5186643, 0.5194529, 
    0.5208794, 0.5241494, 0.5223839, 0.5244485, 0.5198884, 0.5175217, 
    0.516909, 0.5157661, 0.5169351, 0.51684, 0.5179585, 0.517599, 0.520284, 
    0.5188419, 0.5229378, 0.5244321, 0.5286499, 0.5312346, 0.5338641, 
    0.5350249, 0.5353781, 0.5355257,
  0.5310283, 0.5334976, 0.5330174, 0.5350101, 0.5339045, 0.5352095, 
    0.5315287, 0.5335958, 0.532276, 0.5312504, 0.5388803, 0.535099, 0.542811, 
    0.5403967, 0.5464641, 0.5424354, 0.5472769, 0.5463476, 0.5491446, 
    0.5483431, 0.5519236, 0.5495147, 0.5537806, 0.551348, 0.5517285, 
    0.5494353, 0.5358595, 0.5384095, 0.5357085, 0.536072, 0.5359088, 
    0.5339274, 0.5329295, 0.5308394, 0.5312188, 0.5327538, 0.5362355, 
    0.5350531, 0.5380331, 0.5379658, 0.5412862, 0.5397888, 0.5453737, 
    0.5437855, 0.5483766, 0.5472215, 0.5483223, 0.5479885, 0.5483267, 
    0.5466328, 0.5473585, 0.5458682, 0.5400692, 0.5417727, 0.5366945, 
    0.5336445, 0.5316194, 0.5301831, 0.5303861, 0.5307732, 0.5327628, 
    0.534634, 0.5360606, 0.5370153, 0.5379561, 0.5408059, 0.5423146, 
    0.5456951, 0.5450845, 0.5461187, 0.5471066, 0.548766, 0.5484928, 
    0.5492241, 0.5460913, 0.5481732, 0.5447369, 0.5456765, 0.5382128, 
    0.535372, 0.5341659, 0.5331097, 0.5305422, 0.5323152, 0.5316162, 
    0.5332791, 0.5343363, 0.5338134, 0.5370414, 0.5357862, 0.542404, 
    0.5395521, 0.5469913, 0.5452098, 0.5474184, 0.5462912, 0.5482229, 
    0.5464844, 0.5494963, 0.5501525, 0.5497041, 0.5514268, 0.546388, 
    0.5483224, 0.5337988, 0.533884, 0.5342813, 0.5325354, 0.5324286, 
    0.5308291, 0.5322522, 0.5328584, 0.5343975, 0.5353082, 0.5361742, 
    0.5380787, 0.540207, 0.5431848, 0.5453253, 0.5467609, 0.5458805, 
    0.5466577, 0.5457889, 0.5453817, 0.5499067, 0.5473652, 0.5511789, 
    0.5509678, 0.5492415, 0.5509916, 0.5339439, 0.5334532, 0.5317501, 
    0.5330828, 0.5306549, 0.5320139, 0.5327955, 0.5358126, 0.5364755, 
    0.5370907, 0.5383056, 0.5398654, 0.5426033, 0.5449869, 0.547164, 
    0.5470045, 0.5470606, 0.5475472, 0.5463421, 0.5477451, 0.5479807, 
    0.5473648, 0.5509395, 0.5499179, 0.5509633, 0.550298, 0.5336127, 
    0.5344384, 0.5339922, 0.5348313, 0.5342402, 0.5368696, 0.5376584, 
    0.5413507, 0.5398347, 0.5422475, 0.5400797, 0.5404637, 0.5423266, 
    0.5401968, 0.5448556, 0.5416968, 0.5475661, 0.5444099, 0.5477641, 
    0.5471546, 0.5481636, 0.5490676, 0.550205, 0.5523049, 0.5518185, 
    0.5535751, 0.5356696, 0.5367413, 0.5366468, 0.5377685, 0.5385983, 
    0.5403972, 0.5432844, 0.5421984, 0.5441922, 0.5445926, 0.5415636, 
    0.5434232, 0.5374586, 0.5384218, 0.5378482, 0.5357543, 0.5424489, 
    0.5390118, 0.5453607, 0.543497, 0.5489387, 0.5462316, 0.5515508, 
    0.5538274, 0.5559705, 0.5584775, 0.5373262, 0.5365978, 0.5379019, 
    0.5397071, 0.5413823, 0.5436107, 0.5438387, 0.5442563, 0.5453383, 
    0.5462483, 0.5443886, 0.5464764, 0.5386456, 0.5427473, 0.5363227, 
    0.5382564, 0.5396006, 0.5390106, 0.5420743, 0.5427967, 0.545734, 
    0.5442152, 0.5532655, 0.5492588, 0.560387, 0.5572739, 0.5363435, 
    0.5373236, 0.5407369, 0.5391124, 0.5437594, 0.5449042, 0.5458349, 
    0.5470252, 0.5471537, 0.5478591, 0.5467032, 0.5478134, 0.5436154, 
    0.5454908, 0.5403464, 0.541598, 0.5410221, 0.5403906, 0.5423399, 
    0.5444179, 0.544462, 0.5451286, 0.5470083, 0.5437782, 0.5537835, 
    0.5476019, 0.5383926, 0.5402821, 0.5405517, 0.5398197, 0.5447894, 
    0.542988, 0.5478418, 0.5465294, 0.54868, 0.5476112, 0.547454, 0.5460817, 
    0.5452276, 0.5430706, 0.5413164, 0.5399258, 0.5402491, 0.5417768, 
    0.544545, 0.5471654, 0.5465913, 0.5485165, 0.5434223, 0.5455577, 
    0.5447323, 0.5468848, 0.5421696, 0.5461854, 0.5411439, 0.5415856, 
    0.5429522, 0.5457028, 0.5463111, 0.5469614, 0.5465601, 0.5446153, 
    0.5442966, 0.5429189, 0.5425388, 0.5414894, 0.540621, 0.5414145, 
    0.5422481, 0.5446159, 0.5467512, 0.5490805, 0.5496506, 0.5523751, 
    0.5501575, 0.553818, 0.5507062, 0.5560942, 0.5464178, 0.5506142, 
    0.5430143, 0.5438323, 0.5453125, 0.548709, 0.5468747, 0.5490199, 
    0.5442841, 0.5418296, 0.5411945, 0.5400104, 0.5412216, 0.541123, 
    0.5422824, 0.5419098, 0.5446946, 0.5431985, 0.5474501, 0.5490029, 
    0.553391, 0.5560839, 0.5588265, 0.5600382, 0.560407, 0.5605612,
  0.5352148, 0.5380582, 0.5375048, 0.5398021, 0.5385271, 0.5400322, 
    0.5357906, 0.5381713, 0.5366509, 0.5354704, 0.5442732, 0.5399046, 
    0.5488271, 0.5460284, 0.5530713, 0.5483913, 0.5540172, 0.5529357, 
    0.5561931, 0.5552589, 0.5594364, 0.5566245, 0.5616076, 0.558764, 
    0.5592085, 0.5565319, 0.5407822, 0.5437285, 0.5406079, 0.5410275, 
    0.5408392, 0.5385535, 0.5374035, 0.5349976, 0.535434, 0.5372011, 
    0.5412163, 0.5398516, 0.5432934, 0.5432155, 0.5470589, 0.5453244, 
    0.5518032, 0.5499581, 0.5552979, 0.5539527, 0.5552347, 0.5548458, 
    0.5552398, 0.5532675, 0.5541121, 0.5523781, 0.5456492, 0.5476228, 
    0.5417464, 0.5382274, 0.535895, 0.5342428, 0.5344762, 0.5349215, 
    0.5372114, 0.5393682, 0.5410145, 0.542117, 0.5432043, 0.5465024, 
    0.5482512, 0.5521768, 0.5514671, 0.5526695, 0.5538189, 0.5557517, 
    0.5554333, 0.5562858, 0.5526375, 0.5550609, 0.5510631, 0.5521552, 
    0.5435011, 0.5402196, 0.5388284, 0.5376112, 0.5346558, 0.536696, 
    0.5358914, 0.5378063, 0.5390249, 0.538422, 0.5421472, 0.5406976, 
    0.5483549, 0.5450505, 0.5536848, 0.5516127, 0.554182, 0.5528702, 
    0.5551189, 0.5530949, 0.5566031, 0.5573686, 0.5568454, 0.558856, 
    0.5529828, 0.5552348, 0.5384052, 0.5385035, 0.5389615, 0.5369496, 
    0.5368266, 0.5349857, 0.5366235, 0.5373217, 0.5390955, 0.5401461, 
    0.5411456, 0.5433461, 0.5458087, 0.5492607, 0.5517469, 0.5534166, 
    0.5523924, 0.5532966, 0.5522859, 0.5518125, 0.5570818, 0.5541201, 
    0.5585666, 0.5583201, 0.5563061, 0.5583479, 0.5385725, 0.5380069, 
    0.5360455, 0.5375802, 0.5347854, 0.5363491, 0.5372493, 0.5407281, 
    0.5414935, 0.5422041, 0.5436084, 0.5454132, 0.5485861, 0.5513536, 
    0.5538858, 0.5537, 0.5537654, 0.554332, 0.5529293, 0.5545623, 0.5548368, 
    0.5541196, 0.5582871, 0.5570949, 0.5583149, 0.5575384, 0.5381907, 
    0.5391427, 0.5386282, 0.5395958, 0.5389141, 0.5419488, 0.5428602, 
    0.5471337, 0.5453777, 0.5481734, 0.5456613, 0.5461061, 0.5482651, 
    0.5457968, 0.551201, 0.5475348, 0.554354, 0.5506831, 0.5545844, 
    0.5538749, 0.5550498, 0.5561033, 0.5574298, 0.5598819, 0.5593136, 
    0.5613672, 0.5405631, 0.5418006, 0.5416914, 0.5429875, 0.5439469, 
    0.546029, 0.5493764, 0.5481164, 0.5504304, 0.5508955, 0.5473804, 
    0.5495375, 0.5426292, 0.5437428, 0.5430796, 0.5406608, 0.5484069, 
    0.5444253, 0.5517881, 0.5496231, 0.555953, 0.5528008, 0.5590008, 
    0.5616624, 0.5641723, 0.5671139, 0.5424762, 0.5416348, 0.5431416, 
    0.5452299, 0.5471702, 0.5497551, 0.5500198, 0.5505049, 0.551762, 
    0.5528202, 0.5506585, 0.5530856, 0.5440016, 0.5487531, 0.541317, 
    0.5435515, 0.5451066, 0.5444239, 0.5479724, 0.5488104, 0.5522221, 
    0.5504571, 0.5610051, 0.5563262, 0.5693584, 0.5657008, 0.541341, 
    0.5424732, 0.5464224, 0.5445417, 0.5499278, 0.5512575, 0.5523394, 
    0.5537242, 0.5538737, 0.5546951, 0.5533494, 0.5546418, 0.5497606, 
    0.5519393, 0.5459701, 0.5474203, 0.5467528, 0.5460213, 0.5482805, 
    0.5506925, 0.5507438, 0.5515184, 0.5537045, 0.5499496, 0.5616111, 
    0.5543956, 0.543709, 0.5458956, 0.5462079, 0.5453603, 0.5511241, 
    0.5490324, 0.554675, 0.5531472, 0.5556515, 0.5544064, 0.5542234, 
    0.5526264, 0.5516334, 0.5491282, 0.5470939, 0.5454831, 0.5458574, 
    0.5476276, 0.5508401, 0.5538874, 0.5532192, 0.555461, 0.5495364, 
    0.5520171, 0.5510578, 0.5535609, 0.548083, 0.552747, 0.546894, 0.547406, 
    0.5489909, 0.5521858, 0.5528933, 0.5536499, 0.553183, 0.5509217, 
    0.5505516, 0.5489523, 0.5485112, 0.5472944, 0.5462881, 0.5472076, 
    0.548174, 0.5509226, 0.5534053, 0.5561183, 0.5567831, 0.5599639, 
    0.5573744, 0.5616514, 0.5580148, 0.5643173, 0.5530174, 0.5579073, 
    0.549063, 0.5500124, 0.5517321, 0.5556853, 0.5535491, 0.5560476, 
    0.550537, 0.5476888, 0.5469527, 0.545581, 0.546984, 0.5468699, 0.5482138, 
    0.5477818, 0.5510139, 0.5492766, 0.5542188, 0.5560278, 0.5611519, 
    0.5643051, 0.5675238, 0.5689481, 0.569382, 0.5695634,
  0.5840928, 0.5875039, 0.586839, 0.5896025, 0.5880677, 0.5898799, 0.5847825, 
    0.5876398, 0.585814, 0.5843988, 0.5950066, 0.5897262, 0.6005461, 
    0.5971375, 0.6057423, 0.6000144, 0.606905, 0.6055759, 0.6095858, 
    0.6084337, 0.6135982, 0.6101183, 0.6162958, 0.6127648, 0.6133156, 
    0.610004, 0.5907843, 0.5943465, 0.5905741, 0.5910804, 0.5908531, 
    0.5880995, 0.5867173, 0.5838327, 0.5843552, 0.5864743, 0.5913082, 
    0.5896623, 0.5938194, 0.5937251, 0.598391, 0.5962822, 0.6041864, 
    0.6019276, 0.6084818, 0.6068256, 0.6084039, 0.6079248, 0.6084102, 
    0.6059834, 0.6070218, 0.6048914, 0.5966766, 0.5990776, 0.5919484, 
    0.5877073, 0.5849076, 0.5829297, 0.5832089, 0.5837415, 0.5864867, 
    0.5890799, 0.5910646, 0.5923963, 0.5937116, 0.5977138, 0.5998436, 
    0.6046445, 0.6037745, 0.605249, 0.6066612, 0.6090413, 0.6086487, 
    0.6097001, 0.6052098, 0.6081898, 0.6032797, 0.6046181, 0.594071, 
    0.5901058, 0.5884302, 0.5869668, 0.5834236, 0.5858681, 0.5849032, 
    0.5872012, 0.5886666, 0.5879413, 0.5924327, 0.5906823, 0.59997, 
    0.5959496, 0.6064963, 0.6039529, 0.6071077, 0.6054955, 0.6082612, 
    0.6057714, 0.6100919, 0.6110377, 0.6103912, 0.6128787, 0.6056337, 
    0.608404, 0.5879211, 0.5880393, 0.5885903, 0.5861724, 0.5860248, 
    0.5838185, 0.5857811, 0.5866191, 0.5887516, 0.5900171, 0.5912228, 
    0.5938833, 0.5968704, 0.6010756, 0.6041175, 0.6061666, 0.6049091, 
    0.6060191, 0.6047784, 0.6041978, 0.6106831, 0.6070315, 0.6125202, 
    0.6122149, 0.6097252, 0.6122493, 0.5881223, 0.5874423, 0.585088, 
    0.5869296, 0.5835787, 0.585452, 0.5865321, 0.590719, 0.591643, 0.5925015, 
    0.5942009, 0.5963899, 0.600252, 0.6036355, 0.6067434, 0.606515, 
    0.6065954, 0.6072922, 0.6055681, 0.6075758, 0.6079137, 0.607031, 
    0.612174, 0.6106993, 0.6122084, 0.6112476, 0.5876632, 0.5888084, 
    0.5881893, 0.5893542, 0.5885333, 0.5921929, 0.593295, 0.598482, 
    0.5963468, 0.5997487, 0.5966913, 0.5972318, 0.5998605, 0.596856, 
    0.6034486, 0.5989705, 0.6073193, 0.6028146, 0.607603, 0.6067299, 
    0.6081761, 0.6094749, 0.6111133, 0.614151, 0.6134459, 0.6159966, 0.59052, 
    0.5920138, 0.5918819, 0.5934491, 0.5946111, 0.5971382, 0.6012169, 
    0.5996793, 0.6025052, 0.6030744, 0.5987824, 0.6014137, 0.5930157, 
    0.5943638, 0.5935606, 0.5906379, 0.6000335, 0.5951911, 0.6041679, 
    0.6015183, 0.6092895, 0.6054103, 0.6130582, 0.616364, 0.6194943, 
    0.6231793, 0.5928306, 0.5918136, 0.5936357, 0.5961673, 0.5985264, 
    0.6016796, 0.6020031, 0.6025964, 0.604136, 0.6054341, 0.6027843, 0.60576, 
    0.5946774, 0.6004558, 0.5914298, 0.5941321, 0.5960177, 0.5951895, 
    0.5995038, 0.6005259, 0.6047, 0.6025379, 0.6155463, 0.60975, 0.626003, 
    0.6214069, 0.5914588, 0.592827, 0.5976164, 0.5953322, 0.6018906, 
    0.6035177, 0.604844, 0.6065447, 0.6067286, 0.6077392, 0.6060841, 
    0.6076736, 0.6016863, 0.6043533, 0.5970665, 0.5988309, 0.5980184, 
    0.5971288, 0.5998793, 0.602826, 0.6028888, 0.6038374, 0.6065205, 
    0.6019173, 0.6163, 0.6073705, 0.5943229, 0.596976, 0.5973556, 0.5963256, 
    0.6033544, 0.6007968, 0.6077145, 0.6058357, 0.6089177, 0.6073838, 
    0.6071586, 0.6051962, 0.6039782, 0.6009138, 0.5984336, 0.5964748, 
    0.5969296, 0.5990835, 0.6030067, 0.6067454, 0.6059241, 0.6086828, 
    0.6014123, 0.6044487, 0.6032732, 0.6063439, 0.5996386, 0.6053442, 
    0.5981902, 0.5988135, 0.6007461, 0.6046556, 0.6055239, 0.6064534, 
    0.6058795, 0.6031066, 0.6026536, 0.6006989, 0.6001608, 0.5986777, 
    0.5974532, 0.598572, 0.5997495, 0.6031076, 0.6061528, 0.6094934, 
    0.6103141, 0.6142528, 0.6110448, 0.6163503, 0.6118369, 0.6196755, 
    0.6056762, 0.611704, 0.6008341, 0.6019941, 0.6040992, 0.6089593, 
    0.6063294, 0.6094062, 0.6026358, 0.5991581, 0.5982616, 0.5965938, 
    0.5982998, 0.5981608, 0.5997981, 0.5992714, 0.6032195, 0.601095, 
    0.6071531, 0.6093818, 0.6157289, 0.6196603, 0.6236942, 0.6254861, 
    0.6260327, 0.6262615,
  0.662225, 0.6677868, 0.6666974, 0.6712427, 0.6687127, 0.6717014, 0.6633441, 
    0.6680099, 0.665023, 0.6627212, 0.680266, 0.671447, 0.6897113, 0.683875, 
    0.6987641, 0.6887957, 0.7008164, 0.698471, 0.7055875, 0.7035305, 
    0.7128335, 0.706542, 0.7177785, 0.7113178, 0.712319, 0.7063369, 
    0.6732004, 0.6791539, 0.6728516, 0.6736922, 0.6733146, 0.6687649, 
    0.6664983, 0.6618037, 0.6626505, 0.6661009, 0.674071, 0.6713414, 
    0.6782679, 0.6781096, 0.6860121, 0.6824228, 0.6960331, 0.6920994, 
    0.703616, 0.700676, 0.7034774, 0.7026249, 0.7034885, 0.6991888, 
    0.7010232, 0.6972683, 0.6830918, 0.6871873, 0.6751373, 0.6681207, 
    0.6635474, 0.6603436, 0.6607946, 0.6616561, 0.6661212, 0.6703797, 
    0.673666, 0.6758847, 0.6780869, 0.6848563, 0.6885019, 0.6968353, 
    0.695313, 0.6978962, 0.7003852, 0.704614, 0.7039136, 0.7057922, 
    0.6978274, 0.7030962, 0.6944495, 0.6967888, 0.6786906, 0.6720753, 
    0.6693089, 0.6669066, 0.6611418, 0.6651112, 0.6635403, 0.6672907, 
    0.6696983, 0.668505, 0.6759456, 0.673031, 0.6887194, 0.6818594, 
    0.7000937, 0.6956248, 0.7011753, 0.6983294, 0.7032232, 0.6988151, 
    0.7064945, 0.7081947, 0.7070318, 0.7115247, 0.6985728, 0.7034776, 
    0.6684718, 0.6686661, 0.6695726, 0.6656078, 0.6653668, 0.6617806, 
    0.6649694, 0.6663377, 0.6698383, 0.6719286, 0.6739291, 0.6783752, 
    0.6834211, 0.6906249, 0.6959124, 0.6995118, 0.6972992, 0.6992517, 
    0.6970699, 0.696053, 0.7075566, 0.7010404, 0.7108741, 0.7103208, 
    0.7058372, 0.7103831, 0.6688025, 0.6676857, 0.6638407, 0.6668457, 
    0.6613926, 0.6644331, 0.6661955, 0.6730921, 0.6746283, 0.6760604, 
    0.6789089, 0.6826055, 0.6892046, 0.6950702, 0.7005305, 0.7001269, 
    0.700269, 0.7015022, 0.6984574, 0.7020051, 0.7026051, 0.7010394, 
    0.7102469, 0.7075857, 0.7103091, 0.7085731, 0.6680483, 0.6699319, 
    0.6689126, 0.6708323, 0.6694788, 0.6755452, 0.6773883, 0.6861677, 
    0.6825324, 0.6883389, 0.6831169, 0.6840355, 0.6885312, 0.6833965, 
    0.6947441, 0.6870037, 0.7015502, 0.6936396, 0.7020534, 0.7005067, 
    0.7030718, 0.7053891, 0.708331, 0.7138419, 0.7125561, 0.7172271, 
    0.6727619, 0.6752464, 0.6750264, 0.6776465, 0.6795993, 0.6838762, 
    0.690869, 0.6882196, 0.6931018, 0.694092, 0.6866816, 0.6912094, 
    0.6769204, 0.679183, 0.6778335, 0.6729574, 0.6888286, 0.6805772, 
    0.6960006, 0.6913904, 0.7050576, 0.6981798, 0.7118508, 0.7179043, 
    0.7237218, 0.7306814, 0.6766106, 0.6749126, 0.6779595, 0.6822281, 
    0.6862437, 0.6916696, 0.6922303, 0.6932602, 0.6959448, 0.6982216, 
    0.6935871, 0.6987951, 0.679711, 0.6895557, 0.6742734, 0.6787932, 
    0.6819746, 0.6805744, 0.6879182, 0.6896763, 0.6969326, 0.6931586, 
    0.7163985, 0.7058816, 0.7360994, 0.7273186, 0.6743217, 0.6766046, 
    0.6846904, 0.6808155, 0.6920352, 0.6948647, 0.697185, 0.7001794, 
    0.7005042, 0.7022953, 0.6993663, 0.7021788, 0.6916813, 0.6963251, 
    0.6837544, 0.6867647, 0.6853759, 0.6838603, 0.6885634, 0.6936595, 
    0.6937687, 0.6954227, 0.7001365, 0.6920815, 0.7177864, 0.701641, 
    0.6791142, 0.6836005, 0.6842462, 0.6824965, 0.6945798, 0.6901435, 
    0.7022514, 0.6989284, 0.7043933, 0.7016647, 0.7012655, 0.6978033, 
    0.6956689, 0.6903456, 0.6860849, 0.6827495, 0.6835217, 0.6871973, 
    0.693974, 0.700534, 0.6990843, 0.7039743, 0.6912071, 0.6964921, 
    0.6944382, 0.6998247, 0.6881497, 0.6980636, 0.6856692, 0.6867349, 
    0.6900561, 0.6968546, 0.6983795, 0.700018, 0.6990057, 0.694148, 
    0.6933596, 0.6899748, 0.6890475, 0.6865025, 0.6844124, 0.6863216, 
    0.6883402, 0.6941498, 0.6994875, 0.7054223, 0.7068934, 0.7140279, 
    0.7082076, 0.7178791, 0.709637, 0.7240613, 0.6986476, 0.7093968, 
    0.690208, 0.6922146, 0.6958805, 0.7044677, 0.6997991, 0.7052664, 
    0.6933287, 0.6873253, 0.6857911, 0.6829513, 0.6858563, 0.6856189, 
    0.6884237, 0.6875194, 0.6943446, 0.6906585, 0.7012556, 0.7052225, 
    0.7167342, 0.7240328, 0.7316638, 0.7351018, 0.7361567, 0.736599,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 XSMRPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 XSMRPOOL_RECOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZBOT =
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5 ;

 ZWT =
  8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882 ;

 ZWT_CH4_UNSAT =
  0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01157327, 0.01857286, 
    0.01857286, 0.01857286, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01952015, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01952015, 0.01952015, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01952015, 0.01952015, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01952015, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01952015, 0.01952015, 0.01952015, 0.01952015, 
    0.01857286, 0.01952015, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01157327, 0.01157327, 0.01157327, 0.01952015, 0.01952015, 
    0.01952015, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01952015, 0.01857286, 
    0.01952015, 0.01952015, 0.01857286, 0.01952015, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01157327, 0.01157327, 
    0.01952015, 0.01952015, 0.01857286, 0.01952015, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01157327, 0.01857286, 0.01952015, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01157327, 0.01857286, 0.01157327, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 0.01857286, 
    0.01857286, 0.01857286, 0.01857286, 0.01157327, 0.01157327, 0.01157327, 
    0.01157327, 0.01157327 ;

 ZWT_PERCH =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 o2_decomp_depth_unsat =
  3.415385e-11, 3.430415e-11, 3.427484e-11, 3.439615e-11, 3.432881e-11, 
    3.44082e-11, 3.418413e-11, 3.430988e-11, 3.422954e-11, 3.416707e-11, 
    3.463152e-11, 3.440128e-11, 3.487098e-11, 3.472383e-11, 3.509349e-11, 
    3.484798e-11, 3.5143e-11, 3.508631e-11, 3.525682e-11, 3.520789e-11, 
    3.542612e-11, 3.527928e-11, 3.553931e-11, 3.539098e-11, 3.541413e-11, 
    3.527426e-11, 3.444784e-11, 3.460311e-11, 3.443858e-11, 3.446072e-11, 
    3.445074e-11, 3.433005e-11, 3.426927e-11, 3.414204e-11, 3.416508e-11, 
    3.425849e-11, 3.447041e-11, 3.439837e-11, 3.457979e-11, 3.45757e-11, 
    3.477788e-11, 3.468667e-11, 3.502691e-11, 3.493008e-11, 3.520989e-11, 
    3.513942e-11, 3.520651e-11, 3.51861e-11, 3.520667e-11, 3.510341e-11, 
    3.514757e-11, 3.505674e-11, 3.470418e-11, 3.48079e-11, 3.449855e-11, 
    3.431278e-11, 3.418949e-11, 3.410211e-11, 3.411438e-11, 3.413794e-11, 
    3.425897e-11, 3.437283e-11, 3.445968e-11, 3.451776e-11, 3.457501e-11, 
    3.474858e-11, 3.484046e-11, 3.504641e-11, 3.500919e-11, 3.507216e-11, 
    3.513237e-11, 3.523348e-11, 3.521681e-11, 3.526133e-11, 3.50703e-11, 
    3.519722e-11, 3.498769e-11, 3.504496e-11, 3.459095e-11, 3.441795e-11, 
    3.434448e-11, 3.428015e-11, 3.412386e-11, 3.423175e-11, 3.418917e-11, 
    3.429033e-11, 3.435466e-11, 3.432278e-11, 3.45193e-11, 3.444281e-11, 
    3.484585e-11, 3.467212e-11, 3.512539e-11, 3.501675e-11, 3.515132e-11, 
    3.508262e-11, 3.520029e-11, 3.509432e-11, 3.527785e-11, 3.531787e-11, 
    3.529045e-11, 3.53955e-11, 3.508822e-11, 3.520615e-11, 3.43221e-11, 
    3.432729e-11, 3.435143e-11, 3.424509e-11, 3.423858e-11, 3.414119e-11, 
    3.422775e-11, 3.426465e-11, 3.43583e-11, 3.441369e-11, 3.446636e-11, 
    3.458236e-11, 3.471194e-11, 3.489331e-11, 3.502374e-11, 3.511119e-11, 
    3.505751e-11, 3.510483e-11, 3.505186e-11, 3.502698e-11, 3.530277e-11, 
    3.514784e-11, 3.538028e-11, 3.536741e-11, 3.526211e-11, 3.536876e-11, 
    3.433087e-11, 3.430094e-11, 3.419727e-11, 3.427833e-11, 3.413052e-11, 
    3.421323e-11, 3.426074e-11, 3.444436e-11, 3.448469e-11, 3.452215e-11, 
    3.45961e-11, 3.469106e-11, 3.485784e-11, 3.500303e-11, 3.513573e-11, 
    3.512594e-11, 3.512935e-11, 3.515896e-11, 3.508548e-11, 3.517095e-11, 
    3.518525e-11, 3.514773e-11, 3.536559e-11, 3.53033e-11, 3.536699e-11, 
    3.532638e-11, 3.431061e-11, 3.436082e-11, 3.433361e-11, 3.43847e-11, 
    3.434863e-11, 3.450873e-11, 3.455671e-11, 3.478158e-11, 3.468919e-11, 
    3.483619e-11, 3.470404e-11, 3.472744e-11, 3.484086e-11, 3.471108e-11, 
    3.499491e-11, 3.480237e-11, 3.516007e-11, 3.496762e-11, 3.517206e-11, 
    3.513485e-11, 3.519631e-11, 3.525143e-11, 3.53207e-11, 3.544874e-11, 
    3.5419e-11, 3.552613e-11, 3.443574e-11, 3.450094e-11, 3.449517e-11, 
    3.456343e-11, 3.461392e-11, 3.472352e-11, 3.489938e-11, 3.483315e-11, 
    3.49546e-11, 3.497899e-11, 3.479435e-11, 3.490766e-11, 3.454425e-11, 
    3.460285e-11, 3.456791e-11, 3.444034e-11, 3.484809e-11, 3.463864e-11, 
    3.502547e-11, 3.491184e-11, 3.524346e-11, 3.507844e-11, 3.540265e-11, 
    3.554147e-11, 3.567215e-11, 3.582498e-11, 3.453652e-11, 3.449211e-11, 
    3.457148e-11, 3.468143e-11, 3.478341e-11, 3.491921e-11, 3.493306e-11, 
    3.495845e-11, 3.502433e-11, 3.507981e-11, 3.496642e-11, 3.509361e-11, 
    3.461641e-11, 3.486627e-11, 3.447487e-11, 3.459263e-11, 3.467444e-11, 
    3.463852e-11, 3.482512e-11, 3.486908e-11, 3.504801e-11, 3.495548e-11, 
    3.550709e-11, 3.52628e-11, 3.594139e-11, 3.57515e-11, 3.447658e-11, 
    3.453621e-11, 3.474406e-11, 3.464512e-11, 3.492817e-11, 3.499792e-11, 
    3.505457e-11, 3.512713e-11, 3.513488e-11, 3.517789e-11, 3.510735e-11, 
    3.517504e-11, 3.49191e-11, 3.503339e-11, 3.471989e-11, 3.479608e-11, 
    3.476099e-11, 3.472246e-11, 3.484117e-11, 3.496779e-11, 3.497045e-11, 
    3.501099e-11, 3.512549e-11, 3.492865e-11, 3.553851e-11, 3.516155e-11, 
    3.460128e-11, 3.47163e-11, 3.473269e-11, 3.468811e-11, 3.499082e-11, 
    3.488107e-11, 3.517684e-11, 3.509678e-11, 3.522784e-11, 3.516269e-11, 
    3.515302e-11, 3.506938e-11, 3.501724e-11, 3.488581e-11, 3.477885e-11, 
    3.469415e-11, 3.471376e-11, 3.480683e-11, 3.497543e-11, 3.513514e-11, 
    3.51001e-11, 3.521742e-11, 3.490688e-11, 3.503701e-11, 3.498662e-11, 
    3.511783e-11, 3.483124e-11, 3.507591e-11, 3.476872e-11, 3.479557e-11, 
    3.487878e-11, 3.504639e-11, 3.508341e-11, 3.512304e-11, 3.509851e-11, 
    3.497997e-11, 3.496052e-11, 3.487652e-11, 3.48533e-11, 3.478938e-11, 
    3.473639e-11, 3.478474e-11, 3.483544e-11, 3.497973e-11, 3.510982e-11, 
    3.525177e-11, 3.528652e-11, 3.545254e-11, 3.531732e-11, 3.554043e-11, 
    3.535066e-11, 3.56792e-11, 3.508999e-11, 3.534583e-11, 3.488258e-11, 
    3.493237e-11, 3.502253e-11, 3.522951e-11, 3.511766e-11, 3.524843e-11, 
    3.495974e-11, 3.481011e-11, 3.477138e-11, 3.469925e-11, 3.477296e-11, 
    3.476696e-11, 3.483755e-11, 3.48148e-11, 3.498442e-11, 3.489328e-11, 
    3.51523e-11, 3.524696e-11, 3.551448e-11, 3.567864e-11, 3.584593e-11, 
    3.591978e-11, 3.594226e-11, 3.595163e-11,
  1.907756e-11, 1.922153e-11, 1.919351e-11, 1.930986e-11, 1.924529e-11, 
    1.932152e-11, 1.910672e-11, 1.922726e-11, 1.915028e-11, 1.909051e-11, 
    1.953639e-11, 1.931506e-11, 1.976728e-11, 1.962541e-11, 1.99825e-11, 
    1.974518e-11, 2.003047e-11, 1.997564e-11, 2.014085e-11, 2.009347e-11, 
    2.03053e-11, 2.016273e-11, 2.041543e-11, 2.027122e-11, 2.029376e-11, 
    2.015803e-11, 1.935953e-11, 1.950878e-11, 1.93507e-11, 1.937196e-11, 
    1.936242e-11, 1.924662e-11, 1.918836e-11, 1.906657e-11, 1.908866e-11, 
    1.917813e-11, 1.938152e-11, 1.931239e-11, 1.948679e-11, 1.948284e-11, 
    1.967766e-11, 1.958973e-11, 1.991821e-11, 1.982466e-11, 2.009545e-11, 
    2.002722e-11, 2.009224e-11, 2.007252e-11, 2.00925e-11, 1.999247e-11, 
    2.003531e-11, 1.994737e-11, 1.960619e-11, 1.970624e-11, 1.940838e-11, 
    1.923008e-11, 1.9112e-11, 1.902837e-11, 1.904018e-11, 1.906271e-11, 
    1.917865e-11, 1.92879e-11, 1.937131e-11, 1.942717e-11, 1.948228e-11, 
    1.964941e-11, 1.973808e-11, 1.993715e-11, 1.990117e-11, 1.996213e-11, 
    2.002044e-11, 2.011846e-11, 2.010232e-11, 2.014554e-11, 1.996053e-11, 
    2.008342e-11, 1.988069e-11, 1.993606e-11, 1.949725e-11, 1.933103e-11, 
    1.926052e-11, 1.91989e-11, 1.904927e-11, 1.915255e-11, 1.911181e-11, 
    1.920879e-11, 1.927051e-11, 1.923998e-11, 1.94287e-11, 1.935525e-11, 
    1.974334e-11, 1.957584e-11, 2.001363e-11, 1.990855e-11, 2.003885e-11, 
    1.997233e-11, 2.008636e-11, 1.998372e-11, 2.016164e-11, 2.020045e-11, 
    2.017393e-11, 2.02759e-11, 1.997803e-11, 2.009224e-11, 1.923912e-11, 
    1.92441e-11, 1.92673e-11, 1.916539e-11, 1.915917e-11, 1.906597e-11, 
    1.914889e-11, 1.918424e-11, 1.927409e-11, 1.932731e-11, 1.937795e-11, 
    1.948946e-11, 1.961427e-11, 1.978928e-11, 1.991536e-11, 2.000004e-11, 
    1.99481e-11, 1.999395e-11, 1.99427e-11, 1.991869e-11, 2.018591e-11, 
    2.00357e-11, 2.026122e-11, 2.024872e-11, 2.014657e-11, 2.025013e-11, 
    1.924759e-11, 1.921895e-11, 1.911962e-11, 1.919734e-11, 1.905583e-11, 
    1.913499e-11, 1.918056e-11, 1.935678e-11, 1.939558e-11, 1.943158e-11, 
    1.950275e-11, 1.959423e-11, 1.975507e-11, 1.989541e-11, 2.002383e-11, 
    2.001441e-11, 2.001773e-11, 2.004645e-11, 1.997533e-11, 2.005814e-11, 
    2.007205e-11, 2.003569e-11, 2.024705e-11, 2.018658e-11, 2.024846e-11, 
    2.020908e-11, 1.922826e-11, 1.927647e-11, 1.925042e-11, 1.929943e-11, 
    1.926489e-11, 1.941863e-11, 1.946481e-11, 1.968143e-11, 1.959243e-11, 
    1.973415e-11, 1.960681e-11, 1.962935e-11, 1.973877e-11, 1.961368e-11, 
    1.988766e-11, 1.970176e-11, 2.004757e-11, 1.986139e-11, 2.005926e-11, 
    2.002328e-11, 2.008287e-11, 2.013629e-11, 2.020357e-11, 2.032792e-11, 
    2.02991e-11, 2.040325e-11, 1.934844e-11, 1.941112e-11, 1.940561e-11, 
    1.947128e-11, 1.951991e-11, 1.962545e-11, 1.979516e-11, 1.973128e-11, 
    1.984861e-11, 1.987218e-11, 1.969396e-11, 1.980332e-11, 1.945312e-11, 
    1.950955e-11, 1.947595e-11, 1.935338e-11, 1.974599e-11, 1.954414e-11, 
    1.991744e-11, 1.980767e-11, 2.012867e-11, 1.996879e-11, 2.028324e-11, 
    2.041819e-11, 2.054549e-11, 2.06946e-11, 1.944537e-11, 1.940274e-11, 
    1.94791e-11, 1.958492e-11, 1.96833e-11, 1.981436e-11, 1.982779e-11, 
    1.985238e-11, 1.991613e-11, 1.996979e-11, 1.986016e-11, 1.998325e-11, 
    1.952263e-11, 1.976354e-11, 1.938663e-11, 1.949984e-11, 1.957868e-11, 
    1.954409e-11, 1.972398e-11, 1.976647e-11, 1.993944e-11, 1.984996e-11, 
    2.038485e-11, 2.014757e-11, 2.080839e-11, 2.062297e-11, 1.938785e-11, 
    1.944522e-11, 1.964538e-11, 1.955005e-11, 1.982312e-11, 1.989054e-11, 
    1.994541e-11, 2.001563e-11, 2.002322e-11, 2.006487e-11, 1.999663e-11, 
    2.006217e-11, 1.981464e-11, 1.992512e-11, 1.962247e-11, 1.969598e-11, 
    1.966215e-11, 1.962506e-11, 1.97396e-11, 1.986188e-11, 1.98645e-11, 
    1.990376e-11, 2.001456e-11, 1.982423e-11, 2.041554e-11, 2.004961e-11, 
    1.950786e-11, 1.961866e-11, 1.963451e-11, 1.959155e-11, 1.988377e-11, 
    1.977771e-11, 2.006386e-11, 1.998638e-11, 2.011338e-11, 2.005023e-11, 
    2.004095e-11, 1.995996e-11, 1.99096e-11, 1.978257e-11, 1.967943e-11, 
    1.959778e-11, 1.961676e-11, 1.970648e-11, 1.986937e-11, 2.00239e-11, 
    1.999001e-11, 2.010372e-11, 1.980327e-11, 1.992905e-11, 1.98804e-11, 
    2.000735e-11, 1.972958e-11, 1.996601e-11, 1.966931e-11, 1.969526e-11, 
    1.977561e-11, 1.993759e-11, 1.99735e-11, 2.001186e-11, 1.998819e-11, 
    1.987351e-11, 1.985475e-11, 1.977366e-11, 1.975129e-11, 1.968961e-11, 
    1.963859e-11, 1.96852e-11, 1.973419e-11, 1.987356e-11, 1.999946e-11, 
    2.013705e-11, 2.017077e-11, 2.033204e-11, 2.020072e-11, 2.041758e-11, 
    2.023315e-11, 2.055279e-11, 1.997975e-11, 2.022774e-11, 1.977927e-11, 
    1.982741e-11, 1.991459e-11, 2.011507e-11, 2.000675e-11, 2.013345e-11, 
    1.985401e-11, 1.970958e-11, 1.967228e-11, 1.960274e-11, 1.967387e-11, 
    1.966808e-11, 1.973622e-11, 1.971431e-11, 1.987819e-11, 1.979011e-11, 
    2.004071e-11, 2.013245e-11, 2.039232e-11, 2.055221e-11, 2.071542e-11, 
    2.078761e-11, 2.08096e-11, 2.081879e-11,
  1.784466e-11, 1.800237e-11, 1.797167e-11, 1.80992e-11, 1.802841e-11, 
    1.811199e-11, 1.787659e-11, 1.800864e-11, 1.79243e-11, 1.785884e-11, 
    1.834779e-11, 1.81049e-11, 1.860153e-11, 1.844557e-11, 1.88384e-11, 
    1.857722e-11, 1.889124e-11, 1.883084e-11, 1.901289e-11, 1.896066e-11, 
    1.919428e-11, 1.903701e-11, 1.931586e-11, 1.915668e-11, 1.918154e-11, 
    1.903183e-11, 1.815368e-11, 1.831747e-11, 1.814399e-11, 1.81673e-11, 
    1.815684e-11, 1.802987e-11, 1.796603e-11, 1.783264e-11, 1.785683e-11, 
    1.795481e-11, 1.817779e-11, 1.810197e-11, 1.829332e-11, 1.828899e-11, 
    1.850299e-11, 1.840637e-11, 1.876761e-11, 1.866464e-11, 1.896284e-11, 
    1.888766e-11, 1.89593e-11, 1.893757e-11, 1.895959e-11, 1.884938e-11, 
    1.889656e-11, 1.879971e-11, 1.842445e-11, 1.853441e-11, 1.820727e-11, 
    1.801174e-11, 1.788238e-11, 1.779081e-11, 1.780375e-11, 1.782841e-11, 
    1.795539e-11, 1.807512e-11, 1.816659e-11, 1.822789e-11, 1.828837e-11, 
    1.847194e-11, 1.856942e-11, 1.878846e-11, 1.874885e-11, 1.881597e-11, 
    1.888019e-11, 1.89882e-11, 1.897041e-11, 1.901806e-11, 1.88142e-11, 
    1.894958e-11, 1.872631e-11, 1.878727e-11, 1.830481e-11, 1.812242e-11, 
    1.804511e-11, 1.797757e-11, 1.781369e-11, 1.792679e-11, 1.788217e-11, 
    1.798841e-11, 1.805605e-11, 1.802259e-11, 1.822957e-11, 1.814898e-11, 
    1.857521e-11, 1.839111e-11, 1.887269e-11, 1.875698e-11, 1.890047e-11, 
    1.88272e-11, 1.895282e-11, 1.883974e-11, 1.903581e-11, 1.907861e-11, 
    1.904935e-11, 1.916184e-11, 1.883348e-11, 1.89593e-11, 1.802165e-11, 
    1.80271e-11, 1.805254e-11, 1.794086e-11, 1.793404e-11, 1.783198e-11, 
    1.792278e-11, 1.796151e-11, 1.805998e-11, 1.811833e-11, 1.817387e-11, 
    1.829625e-11, 1.843333e-11, 1.862573e-11, 1.876447e-11, 1.885771e-11, 
    1.880052e-11, 1.885101e-11, 1.879457e-11, 1.876814e-11, 1.906257e-11, 
    1.8897e-11, 1.914564e-11, 1.913185e-11, 1.901919e-11, 1.91334e-11, 
    1.803094e-11, 1.799954e-11, 1.789072e-11, 1.797586e-11, 1.782088e-11, 
    1.790756e-11, 1.795748e-11, 1.815066e-11, 1.819322e-11, 1.823272e-11, 
    1.831085e-11, 1.841131e-11, 1.858811e-11, 1.874251e-11, 1.888393e-11, 
    1.887355e-11, 1.88772e-11, 1.890885e-11, 1.88305e-11, 1.892173e-11, 
    1.893705e-11, 1.889699e-11, 1.913e-11, 1.906331e-11, 1.913156e-11, 
    1.908812e-11, 1.800974e-11, 1.806259e-11, 1.803403e-11, 1.808776e-11, 
    1.80499e-11, 1.821851e-11, 1.826919e-11, 1.850714e-11, 1.840933e-11, 
    1.856509e-11, 1.842513e-11, 1.84499e-11, 1.857018e-11, 1.843268e-11, 
    1.873398e-11, 1.852948e-11, 1.891008e-11, 1.870506e-11, 1.892296e-11, 
    1.888332e-11, 1.894897e-11, 1.900785e-11, 1.908204e-11, 1.921924e-11, 
    1.918743e-11, 1.930241e-11, 1.814151e-11, 1.821028e-11, 1.820422e-11, 
    1.82763e-11, 1.832968e-11, 1.844561e-11, 1.863219e-11, 1.856194e-11, 
    1.869099e-11, 1.871695e-11, 1.852091e-11, 1.864117e-11, 1.825637e-11, 
    1.831831e-11, 1.828142e-11, 1.814692e-11, 1.857811e-11, 1.835629e-11, 
    1.876677e-11, 1.864595e-11, 1.899945e-11, 1.88233e-11, 1.916993e-11, 
    1.931891e-11, 1.945956e-11, 1.962445e-11, 1.824786e-11, 1.820108e-11, 
    1.828488e-11, 1.840109e-11, 1.850919e-11, 1.865332e-11, 1.866809e-11, 
    1.869515e-11, 1.876532e-11, 1.882441e-11, 1.870371e-11, 1.883923e-11, 
    1.833268e-11, 1.859742e-11, 1.81834e-11, 1.830766e-11, 1.839423e-11, 
    1.835623e-11, 1.855392e-11, 1.860063e-11, 1.879099e-11, 1.869249e-11, 
    1.928209e-11, 1.90203e-11, 1.975039e-11, 1.954522e-11, 1.818474e-11, 
    1.82477e-11, 1.846751e-11, 1.836279e-11, 1.866295e-11, 1.873715e-11, 
    1.879756e-11, 1.887489e-11, 1.888325e-11, 1.892914e-11, 1.885396e-11, 
    1.892617e-11, 1.865362e-11, 1.877521e-11, 1.844234e-11, 1.852313e-11, 
    1.848594e-11, 1.844519e-11, 1.857109e-11, 1.87056e-11, 1.870849e-11, 
    1.875171e-11, 1.887371e-11, 1.866417e-11, 1.931598e-11, 1.891234e-11, 
    1.831645e-11, 1.843816e-11, 1.845558e-11, 1.840837e-11, 1.87297e-11, 
    1.861301e-11, 1.892802e-11, 1.884267e-11, 1.898261e-11, 1.891301e-11, 
    1.890278e-11, 1.881358e-11, 1.875813e-11, 1.861835e-11, 1.850494e-11, 
    1.841521e-11, 1.843606e-11, 1.853468e-11, 1.871384e-11, 1.8884e-11, 
    1.884667e-11, 1.897195e-11, 1.864112e-11, 1.877955e-11, 1.872599e-11, 
    1.886577e-11, 1.856007e-11, 1.882024e-11, 1.849381e-11, 1.852234e-11, 
    1.861069e-11, 1.878895e-11, 1.882849e-11, 1.887074e-11, 1.884466e-11, 
    1.87184e-11, 1.869775e-11, 1.860854e-11, 1.858394e-11, 1.851612e-11, 
    1.846005e-11, 1.851128e-11, 1.856514e-11, 1.871846e-11, 1.885708e-11, 
    1.900869e-11, 1.904588e-11, 1.922379e-11, 1.90789e-11, 1.931824e-11, 
    1.911467e-11, 1.946763e-11, 1.883537e-11, 1.910871e-11, 1.861472e-11, 
    1.866768e-11, 1.876362e-11, 1.898446e-11, 1.886511e-11, 1.900473e-11, 
    1.869695e-11, 1.853808e-11, 1.849708e-11, 1.842066e-11, 1.849882e-11, 
    1.849246e-11, 1.856737e-11, 1.854329e-11, 1.872356e-11, 1.862663e-11, 
    1.890253e-11, 1.900362e-11, 1.929034e-11, 1.946698e-11, 1.964748e-11, 
    1.972738e-11, 1.975172e-11, 1.97619e-11,
  1.830175e-11, 1.847542e-11, 1.84416e-11, 1.858212e-11, 1.850411e-11, 
    1.859621e-11, 1.833689e-11, 1.848233e-11, 1.838942e-11, 1.831735e-11, 
    1.88563e-11, 1.858841e-11, 1.91365e-11, 1.896423e-11, 1.939841e-11, 
    1.910965e-11, 1.945689e-11, 1.939005e-11, 1.959154e-11, 1.953371e-11, 
    1.979252e-11, 1.961825e-11, 1.992732e-11, 1.975083e-11, 1.977839e-11, 
    1.961252e-11, 1.864217e-11, 1.882285e-11, 1.863149e-11, 1.86572e-11, 
    1.864566e-11, 1.850572e-11, 1.843539e-11, 1.828851e-11, 1.831513e-11, 
    1.842303e-11, 1.866876e-11, 1.858517e-11, 1.879618e-11, 1.87914e-11, 
    1.902763e-11, 1.892095e-11, 1.93201e-11, 1.920625e-11, 1.953612e-11, 
    1.945291e-11, 1.953221e-11, 1.950815e-11, 1.953253e-11, 1.941055e-11, 
    1.946277e-11, 1.93556e-11, 1.89409e-11, 1.906234e-11, 1.870126e-11, 
    1.848575e-11, 1.834326e-11, 1.824247e-11, 1.825671e-11, 1.828385e-11, 
    1.842366e-11, 1.855557e-11, 1.86564e-11, 1.8724e-11, 1.879071e-11, 
    1.899336e-11, 1.910102e-11, 1.934316e-11, 1.929935e-11, 1.937359e-11, 
    1.944464e-11, 1.956421e-11, 1.95445e-11, 1.959727e-11, 1.937163e-11, 
    1.952145e-11, 1.927442e-11, 1.934184e-11, 1.880888e-11, 1.86077e-11, 
    1.852251e-11, 1.84481e-11, 1.826765e-11, 1.839217e-11, 1.834304e-11, 
    1.846003e-11, 1.853456e-11, 1.849768e-11, 1.872585e-11, 1.863698e-11, 
    1.910742e-11, 1.89041e-11, 1.943635e-11, 1.930834e-11, 1.946709e-11, 
    1.938601e-11, 1.952504e-11, 1.939989e-11, 1.961692e-11, 1.966434e-11, 
    1.963193e-11, 1.975655e-11, 1.939296e-11, 1.953221e-11, 1.849665e-11, 
    1.850266e-11, 1.853068e-11, 1.840766e-11, 1.840015e-11, 1.828778e-11, 
    1.838775e-11, 1.84304e-11, 1.853889e-11, 1.86032e-11, 1.866444e-11, 
    1.879941e-11, 1.895071e-11, 1.916324e-11, 1.931663e-11, 1.941977e-11, 
    1.935649e-11, 1.941236e-11, 1.934991e-11, 1.932068e-11, 1.964656e-11, 
    1.946326e-11, 1.97386e-11, 1.972332e-11, 1.959852e-11, 1.972504e-11, 
    1.850689e-11, 1.84723e-11, 1.835245e-11, 1.844621e-11, 1.827556e-11, 
    1.837099e-11, 1.842597e-11, 1.863884e-11, 1.868577e-11, 1.872933e-11, 
    1.881552e-11, 1.89264e-11, 1.912167e-11, 1.929234e-11, 1.944878e-11, 
    1.94373e-11, 1.944134e-11, 1.947636e-11, 1.938966e-11, 1.949061e-11, 
    1.950758e-11, 1.946323e-11, 1.972127e-11, 1.964738e-11, 1.972299e-11, 
    1.967487e-11, 1.848354e-11, 1.854177e-11, 1.851029e-11, 1.856951e-11, 
    1.852778e-11, 1.871367e-11, 1.876957e-11, 1.903222e-11, 1.892421e-11, 
    1.909624e-11, 1.894165e-11, 1.8969e-11, 1.910187e-11, 1.894999e-11, 
    1.928291e-11, 1.90569e-11, 1.947772e-11, 1.925094e-11, 1.949198e-11, 
    1.94481e-11, 1.952077e-11, 1.958597e-11, 1.966814e-11, 1.982018e-11, 
    1.978492e-11, 1.991239e-11, 1.862875e-11, 1.870458e-11, 1.86979e-11, 
    1.87774e-11, 1.88363e-11, 1.896427e-11, 1.917038e-11, 1.909275e-11, 
    1.923538e-11, 1.926407e-11, 1.904743e-11, 1.918031e-11, 1.875541e-11, 
    1.882376e-11, 1.878305e-11, 1.863473e-11, 1.911062e-11, 1.886568e-11, 
    1.931917e-11, 1.918559e-11, 1.957667e-11, 1.938171e-11, 1.976552e-11, 
    1.99307e-11, 2.008675e-11, 2.026986e-11, 1.874603e-11, 1.869443e-11, 
    1.878686e-11, 1.891512e-11, 1.903448e-11, 1.919373e-11, 1.921006e-11, 
    1.923997e-11, 1.931756e-11, 1.938292e-11, 1.924944e-11, 1.939932e-11, 
    1.883963e-11, 1.913196e-11, 1.867494e-11, 1.881201e-11, 1.890754e-11, 
    1.88656e-11, 1.908388e-11, 1.91355e-11, 1.934596e-11, 1.923703e-11, 
    1.988988e-11, 1.959976e-11, 2.04098e-11, 2.018185e-11, 1.867642e-11, 
    1.874585e-11, 1.898846e-11, 1.887284e-11, 1.920438e-11, 1.928641e-11, 
    1.935322e-11, 1.943878e-11, 1.944803e-11, 1.949882e-11, 1.941562e-11, 
    1.949553e-11, 1.919407e-11, 1.932851e-11, 1.896065e-11, 1.904987e-11, 
    1.90088e-11, 1.89638e-11, 1.910285e-11, 1.925154e-11, 1.925472e-11, 
    1.930251e-11, 1.943751e-11, 1.920573e-11, 1.992748e-11, 1.948025e-11, 
    1.88217e-11, 1.895605e-11, 1.897527e-11, 1.892315e-11, 1.927818e-11, 
    1.914918e-11, 1.949758e-11, 1.940312e-11, 1.955801e-11, 1.948097e-11, 
    1.946965e-11, 1.937094e-11, 1.930961e-11, 1.915508e-11, 1.902978e-11, 
    1.89307e-11, 1.895372e-11, 1.906263e-11, 1.926065e-11, 1.944887e-11, 
    1.940756e-11, 1.954622e-11, 1.918025e-11, 1.93333e-11, 1.927408e-11, 
    1.942869e-11, 1.909069e-11, 1.937834e-11, 1.901749e-11, 1.9049e-11, 
    1.914662e-11, 1.934371e-11, 1.938744e-11, 1.943419e-11, 1.940533e-11, 
    1.926569e-11, 1.924285e-11, 1.914424e-11, 1.911706e-11, 1.904213e-11, 
    1.898021e-11, 1.903679e-11, 1.909629e-11, 1.926574e-11, 1.941907e-11, 
    1.95869e-11, 1.962807e-11, 1.982524e-11, 1.966467e-11, 1.992998e-11, 
    1.970432e-11, 2.009572e-11, 1.939507e-11, 1.969769e-11, 1.915107e-11, 
    1.92096e-11, 1.931569e-11, 1.956008e-11, 1.942796e-11, 1.958251e-11, 
    1.924196e-11, 1.90664e-11, 1.90211e-11, 1.893672e-11, 1.902303e-11, 
    1.9016e-11, 1.909875e-11, 1.907214e-11, 1.927138e-11, 1.916423e-11, 
    1.946937e-11, 1.958129e-11, 1.989901e-11, 2.0095e-11, 2.029543e-11, 
    2.038421e-11, 2.041127e-11, 2.042259e-11,
  1.973899e-11, 1.992296e-11, 1.988711e-11, 2.003606e-11, 1.995335e-11, 
    2.0051e-11, 1.97762e-11, 1.993028e-11, 1.983184e-11, 1.97555e-11, 
    2.032694e-11, 2.004272e-11, 2.062455e-11, 2.044151e-11, 2.09031e-11, 
    2.059602e-11, 2.096533e-11, 2.089419e-11, 2.11087e-11, 2.104712e-11, 
    2.132291e-11, 2.113716e-11, 2.146667e-11, 2.127846e-11, 2.130784e-11, 
    2.113105e-11, 2.009972e-11, 2.029144e-11, 2.008839e-11, 2.011566e-11, 
    2.010342e-11, 1.995506e-11, 1.988055e-11, 1.972496e-11, 1.975315e-11, 
    1.986744e-11, 2.012793e-11, 2.003928e-11, 2.02631e-11, 2.025803e-11, 
    2.050885e-11, 2.039554e-11, 2.081977e-11, 2.069868e-11, 2.104969e-11, 
    2.096109e-11, 2.104552e-11, 2.10199e-11, 2.104586e-11, 2.091601e-11, 
    2.097159e-11, 2.085754e-11, 2.041674e-11, 2.054573e-11, 2.01624e-11, 
    1.993392e-11, 1.978295e-11, 1.967622e-11, 1.969129e-11, 1.972004e-11, 
    1.986811e-11, 2.000791e-11, 2.011481e-11, 2.018651e-11, 2.02573e-11, 
    2.047246e-11, 2.058684e-11, 2.084431e-11, 2.07977e-11, 2.087669e-11, 
    2.095229e-11, 2.10796e-11, 2.105861e-11, 2.111481e-11, 2.087459e-11, 
    2.103407e-11, 2.077117e-11, 2.084289e-11, 2.027661e-11, 2.006317e-11, 
    1.997288e-11, 1.9894e-11, 1.970288e-11, 1.983476e-11, 1.978271e-11, 
    1.990665e-11, 1.998563e-11, 1.994654e-11, 2.018847e-11, 2.009422e-11, 
    2.059364e-11, 2.037766e-11, 2.094347e-11, 2.080726e-11, 2.097619e-11, 
    2.088989e-11, 2.103789e-11, 2.090466e-11, 2.113575e-11, 2.118627e-11, 
    2.115174e-11, 2.128454e-11, 2.089729e-11, 2.104553e-11, 1.994545e-11, 
    1.995182e-11, 1.998152e-11, 1.985117e-11, 1.984321e-11, 1.972419e-11, 
    1.983006e-11, 1.987525e-11, 1.999021e-11, 2.00584e-11, 2.012333e-11, 
    2.026653e-11, 2.042715e-11, 2.065297e-11, 2.081607e-11, 2.092582e-11, 
    2.085848e-11, 2.091793e-11, 2.085148e-11, 2.082038e-11, 2.116733e-11, 
    2.097211e-11, 2.126541e-11, 2.124912e-11, 2.111615e-11, 2.125095e-11, 
    1.99563e-11, 1.991964e-11, 1.979268e-11, 1.9892e-11, 1.971125e-11, 
    1.981231e-11, 1.987056e-11, 2.00962e-11, 2.014596e-11, 2.019217e-11, 
    2.028362e-11, 2.040133e-11, 2.060878e-11, 2.079024e-11, 2.095669e-11, 
    2.094447e-11, 2.094877e-11, 2.098606e-11, 2.089378e-11, 2.100123e-11, 
    2.10193e-11, 2.097208e-11, 2.124694e-11, 2.11682e-11, 2.124877e-11, 
    2.119748e-11, 1.993155e-11, 1.999327e-11, 1.995991e-11, 2.002268e-11, 
    1.997845e-11, 2.017556e-11, 2.023488e-11, 2.051374e-11, 2.039901e-11, 
    2.058176e-11, 2.041753e-11, 2.044658e-11, 2.058775e-11, 2.042638e-11, 
    2.078022e-11, 2.053997e-11, 2.098751e-11, 2.074623e-11, 2.100268e-11, 
    2.095597e-11, 2.103334e-11, 2.110278e-11, 2.119031e-11, 2.135239e-11, 
    2.131479e-11, 2.145074e-11, 2.008549e-11, 2.016592e-11, 2.015882e-11, 
    2.024317e-11, 2.030568e-11, 2.044155e-11, 2.066055e-11, 2.057803e-11, 
    2.072965e-11, 2.076017e-11, 2.052988e-11, 2.067111e-11, 2.021985e-11, 
    2.029238e-11, 2.024917e-11, 2.009183e-11, 2.059704e-11, 2.033687e-11, 
    2.081878e-11, 2.067672e-11, 2.109287e-11, 2.088532e-11, 2.129411e-11, 
    2.14703e-11, 2.163684e-11, 2.183246e-11, 2.020989e-11, 2.015514e-11, 
    2.025321e-11, 2.038936e-11, 2.051613e-11, 2.068537e-11, 2.070273e-11, 
    2.073454e-11, 2.081707e-11, 2.08866e-11, 2.074461e-11, 2.090405e-11, 
    2.030924e-11, 2.061971e-11, 2.013448e-11, 2.027991e-11, 2.038132e-11, 
    2.033679e-11, 2.056861e-11, 2.062348e-11, 2.084728e-11, 2.073141e-11, 
    2.142674e-11, 2.111747e-11, 2.198207e-11, 2.173843e-11, 2.013604e-11, 
    2.020969e-11, 2.046724e-11, 2.034447e-11, 2.069669e-11, 2.078393e-11, 
    2.0855e-11, 2.094606e-11, 2.09559e-11, 2.100997e-11, 2.09214e-11, 
    2.100647e-11, 2.068573e-11, 2.082871e-11, 2.04377e-11, 2.053248e-11, 
    2.048884e-11, 2.044105e-11, 2.058877e-11, 2.074685e-11, 2.075022e-11, 
    2.080106e-11, 2.094474e-11, 2.069813e-11, 2.146688e-11, 2.099023e-11, 
    2.029018e-11, 2.043283e-11, 2.045323e-11, 2.039788e-11, 2.077517e-11, 
    2.063801e-11, 2.100865e-11, 2.09081e-11, 2.107299e-11, 2.099096e-11, 
    2.097891e-11, 2.087386e-11, 2.080861e-11, 2.064429e-11, 2.051114e-11, 
    2.04059e-11, 2.043034e-11, 2.054604e-11, 2.075654e-11, 2.09568e-11, 
    2.091283e-11, 2.106043e-11, 2.067104e-11, 2.083382e-11, 2.077082e-11, 
    2.093531e-11, 2.057585e-11, 2.088177e-11, 2.049807e-11, 2.053155e-11, 
    2.063529e-11, 2.08449e-11, 2.089141e-11, 2.094117e-11, 2.091045e-11, 
    2.076189e-11, 2.073761e-11, 2.063276e-11, 2.060388e-11, 2.052426e-11, 
    2.045848e-11, 2.051858e-11, 2.05818e-11, 2.076195e-11, 2.092508e-11, 
    2.110377e-11, 2.114763e-11, 2.135781e-11, 2.118664e-11, 2.146955e-11, 
    2.122892e-11, 2.164645e-11, 2.089955e-11, 2.122183e-11, 2.064002e-11, 
    2.070224e-11, 2.081509e-11, 2.107521e-11, 2.093453e-11, 2.10991e-11, 
    2.073665e-11, 2.055005e-11, 2.050191e-11, 2.041229e-11, 2.050396e-11, 
    2.049649e-11, 2.058441e-11, 2.055613e-11, 2.076795e-11, 2.065401e-11, 
    2.097861e-11, 2.10978e-11, 2.143648e-11, 2.164566e-11, 2.185978e-11, 
    2.195471e-11, 2.198365e-11, 2.199575e-11,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
