netcdf ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-1.clm2.h0.0001-12-02-00000 {
dimensions:
	lndgrid = 338 ;
	gridcell = 338 ;
	landunit = 1352 ;
	column = 5408 ;
	pft = 10816 ;
	levgrnd = 15 ;
	levurb = 5 ;
	levlak = 10 ;
	numrad = 2 ;
	levsno = 5 ;
	ltype = 9 ;
	natpft = 17 ;
	string_length = 8 ;
	levdcmp = 15 ;
	hist_interval = 2 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float levgrnd(levgrnd) ;
		levgrnd:long_name = "coordinate soil levels" ;
		levgrnd:units = "m" ;
	float levlak(levlak) ;
		levlak:long_name = "coordinate lake levels" ;
		levlak:units = "m" ;
	float levdcmp(levdcmp) ;
		levdcmp:long_name = "coordinate soil levels" ;
		levdcmp:units = "m" ;
	float time(time) ;
		time:long_name = "time" ;
		time:units = "days since 0001-12-01 00:00:00" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bounds" ;
	int mcdate(time) ;
		mcdate:long_name = "current date (YYYYMMDD)" ;
	int mcsec(time) ;
		mcsec:long_name = "current seconds of current date" ;
		mcsec:units = "s" ;
	int mdcur(time) ;
		mdcur:long_name = "current day (from base day)" ;
	int mscur(time) ;
		mscur:long_name = "current seconds of current day" ;
	int nstep(time) ;
		nstep:long_name = "time step" ;
	double time_bounds(time, hist_interval) ;
		time_bounds:long_name = "history time interval endpoints" ;
	char date_written(time, string_length) ;
	char time_written(time, string_length) ;
	float lon(lndgrid) ;
		lon:long_name = "coordinate longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = 1.e+36f ;
		lon:missing_value = 1.e+36f ;
	float lat(lndgrid) ;
		lat:long_name = "coordinate latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = 1.e+36f ;
		lat:missing_value = 1.e+36f ;
	float area(lndgrid) ;
		area:long_name = "grid cell areas" ;
		area:units = "km^2" ;
		area:_FillValue = 1.e+36f ;
		area:missing_value = 1.e+36f ;
	float topo(lndgrid) ;
		topo:long_name = "grid cell topography" ;
		topo:units = "m" ;
		topo:_FillValue = 1.e+36f ;
		topo:missing_value = 1.e+36f ;
	float landfrac(lndgrid) ;
		landfrac:long_name = "land fraction" ;
		landfrac:_FillValue = 1.e+36f ;
		landfrac:missing_value = 1.e+36f ;
	int landmask(lndgrid) ;
		landmask:long_name = "land/ocean mask (0.=ocean and 1.=land)" ;
		landmask:_FillValue = -9999 ;
		landmask:missing_value = -9999 ;
	int pftmask(lndgrid) ;
		pftmask:long_name = "pft real/fake mask (0.=fake and 1.=real)" ;
		pftmask:_FillValue = -9999 ;
		pftmask:missing_value = -9999 ;
	float ACTUAL_IMMOB(time, lndgrid) ;
		ACTUAL_IMMOB:long_name = "actual N immobilization" ;
		ACTUAL_IMMOB:units = "gN/m^2/s" ;
		ACTUAL_IMMOB:cell_methods = "time: mean" ;
		ACTUAL_IMMOB:_FillValue = 1.e+36f ;
		ACTUAL_IMMOB:missing_value = 1.e+36f ;
	float AGNPP(time, lndgrid) ;
		AGNPP:long_name = "aboveground NPP" ;
		AGNPP:units = "gC/m^2/s" ;
		AGNPP:cell_methods = "time: mean" ;
		AGNPP:_FillValue = 1.e+36f ;
		AGNPP:missing_value = 1.e+36f ;
	float ALT(time, lndgrid) ;
		ALT:long_name = "current active layer thickness" ;
		ALT:units = "m" ;
		ALT:cell_methods = "time: mean" ;
		ALT:_FillValue = 1.e+36f ;
		ALT:missing_value = 1.e+36f ;
	float ALTMAX(time, lndgrid) ;
		ALTMAX:long_name = "maximum annual active layer thickness" ;
		ALTMAX:units = "m" ;
		ALTMAX:cell_methods = "time: mean" ;
		ALTMAX:_FillValue = 1.e+36f ;
		ALTMAX:missing_value = 1.e+36f ;
	float ALTMAX_LASTYEAR(time, lndgrid) ;
		ALTMAX_LASTYEAR:long_name = "maximum prior year active layer thickness" ;
		ALTMAX_LASTYEAR:units = "m" ;
		ALTMAX_LASTYEAR:cell_methods = "time: mean" ;
		ALTMAX_LASTYEAR:_FillValue = 1.e+36f ;
		ALTMAX_LASTYEAR:missing_value = 1.e+36f ;
	float AR(time, lndgrid) ;
		AR:long_name = "autotrophic respiration (MR + GR)" ;
		AR:units = "gC/m^2/s" ;
		AR:cell_methods = "time: mean" ;
		AR:_FillValue = 1.e+36f ;
		AR:missing_value = 1.e+36f ;
	float BAF_CROP(time, lndgrid) ;
		BAF_CROP:long_name = "fractional area burned for crop" ;
		BAF_CROP:units = "proportion/sec" ;
		BAF_CROP:cell_methods = "time: mean" ;
		BAF_CROP:_FillValue = 1.e+36f ;
		BAF_CROP:missing_value = 1.e+36f ;
	float BAF_PEATF(time, lndgrid) ;
		BAF_PEATF:long_name = "fractional area burned in peatland" ;
		BAF_PEATF:units = "proportion/sec" ;
		BAF_PEATF:cell_methods = "time: mean" ;
		BAF_PEATF:_FillValue = 1.e+36f ;
		BAF_PEATF:missing_value = 1.e+36f ;
	float BCDEP(time, lndgrid) ;
		BCDEP:long_name = "total BC deposition (dry+wet) from atmosphere" ;
		BCDEP:units = "kg/m^2/s" ;
		BCDEP:cell_methods = "time: mean" ;
		BCDEP:_FillValue = 1.e+36f ;
		BCDEP:missing_value = 1.e+36f ;
	float BGNPP(time, lndgrid) ;
		BGNPP:long_name = "belowground NPP" ;
		BGNPP:units = "gC/m^2/s" ;
		BGNPP:cell_methods = "time: mean" ;
		BGNPP:_FillValue = 1.e+36f ;
		BGNPP:missing_value = 1.e+36f ;
	float BTRAN(time, lndgrid) ;
		BTRAN:long_name = "transpiration beta factor" ;
		BTRAN:units = "unitless" ;
		BTRAN:cell_methods = "time: mean" ;
		BTRAN:_FillValue = 1.e+36f ;
		BTRAN:missing_value = 1.e+36f ;
	float BUILDHEAT(time, lndgrid) ;
		BUILDHEAT:long_name = "heat flux from urban building interior to walls and roof" ;
		BUILDHEAT:units = "W/m^2" ;
		BUILDHEAT:cell_methods = "time: mean" ;
		BUILDHEAT:_FillValue = 1.e+36f ;
		BUILDHEAT:missing_value = 1.e+36f ;
	float CH4PROD(time, lndgrid) ;
		CH4PROD:long_name = "Gridcell total production of CH4" ;
		CH4PROD:units = "gC/m2/s" ;
		CH4PROD:cell_methods = "time: mean" ;
		CH4PROD:_FillValue = 1.e+36f ;
		CH4PROD:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_SAT(time, lndgrid) ;
		CH4_SURF_AERE_SAT:long_name = "aerenchyma surface CH4 flux for inundated area; (+ to atm)" ;
		CH4_SURF_AERE_SAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_SAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_UNSAT(time, lndgrid) ;
		CH4_SURF_AERE_UNSAT:long_name = "aerenchyma surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_AERE_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_SAT(time, lndgrid) ;
		CH4_SURF_DIFF_SAT:long_name = "diffusive surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_DIFF_SAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_SAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_UNSAT(time, lndgrid) ;
		CH4_SURF_DIFF_UNSAT:long_name = "diffusive surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_DIFF_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_SAT(time, lndgrid) ;
		CH4_SURF_EBUL_SAT:long_name = "ebullition surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_EBUL_SAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_SAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_UNSAT(time, lndgrid) ;
		CH4_SURF_EBUL_UNSAT:long_name = "ebullition surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_EBUL_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_UNSAT:missing_value = 1.e+36f ;
	float COL_CTRUNC(time, lndgrid) ;
		COL_CTRUNC:long_name = "column-level sink for C truncation" ;
		COL_CTRUNC:units = "gC/m^2" ;
		COL_CTRUNC:cell_methods = "time: mean" ;
		COL_CTRUNC:_FillValue = 1.e+36f ;
		COL_CTRUNC:missing_value = 1.e+36f ;
	float COL_FIRE_CLOSS(time, lndgrid) ;
		COL_FIRE_CLOSS:long_name = "total column-level fire C loss for non-peat fires outside land-type converted region" ;
		COL_FIRE_CLOSS:units = "gC/m^2/s" ;
		COL_FIRE_CLOSS:cell_methods = "time: mean" ;
		COL_FIRE_CLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_CLOSS:missing_value = 1.e+36f ;
	float COL_FIRE_NLOSS(time, lndgrid) ;
		COL_FIRE_NLOSS:long_name = "total column-level fire N loss" ;
		COL_FIRE_NLOSS:units = "gN/m^2/s" ;
		COL_FIRE_NLOSS:cell_methods = "time: mean" ;
		COL_FIRE_NLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_NLOSS:missing_value = 1.e+36f ;
	float COL_NTRUNC(time, lndgrid) ;
		COL_NTRUNC:long_name = "column-level sink for N truncation" ;
		COL_NTRUNC:units = "gN/m^2" ;
		COL_NTRUNC:cell_methods = "time: mean" ;
		COL_NTRUNC:_FillValue = 1.e+36f ;
		COL_NTRUNC:missing_value = 1.e+36f ;
	float CONC_CH4_SAT(time, levgrnd, lndgrid) ;
		CONC_CH4_SAT:long_name = "CH4 soil Concentration for inundated / lake area" ;
		CONC_CH4_SAT:units = "mol/m3" ;
		CONC_CH4_SAT:cell_methods = "time: mean" ;
		CONC_CH4_SAT:_FillValue = 1.e+36f ;
		CONC_CH4_SAT:missing_value = 1.e+36f ;
	float CONC_CH4_UNSAT(time, levgrnd, lndgrid) ;
		CONC_CH4_UNSAT:long_name = "CH4 soil Concentration for non-inundated area" ;
		CONC_CH4_UNSAT:units = "mol/m3" ;
		CONC_CH4_UNSAT:cell_methods = "time: mean" ;
		CONC_CH4_UNSAT:_FillValue = 1.e+36f ;
		CONC_CH4_UNSAT:missing_value = 1.e+36f ;
	float CONC_O2_SAT(time, levgrnd, lndgrid) ;
		CONC_O2_SAT:long_name = "O2 soil Concentration for inundated / lake area" ;
		CONC_O2_SAT:units = "mol/m3" ;
		CONC_O2_SAT:cell_methods = "time: mean" ;
		CONC_O2_SAT:_FillValue = 1.e+36f ;
		CONC_O2_SAT:missing_value = 1.e+36f ;
	float CONC_O2_UNSAT(time, levgrnd, lndgrid) ;
		CONC_O2_UNSAT:long_name = "O2 soil Concentration for non-inundated area" ;
		CONC_O2_UNSAT:units = "mol/m3" ;
		CONC_O2_UNSAT:cell_methods = "time: mean" ;
		CONC_O2_UNSAT:_FillValue = 1.e+36f ;
		CONC_O2_UNSAT:missing_value = 1.e+36f ;
	float CPOOL(time, lndgrid) ;
		CPOOL:long_name = "temporary photosynthate C pool" ;
		CPOOL:units = "gC/m^2" ;
		CPOOL:cell_methods = "time: mean" ;
		CPOOL:_FillValue = 1.e+36f ;
		CPOOL:missing_value = 1.e+36f ;
	float CWDC(time, lndgrid) ;
		CWDC:long_name = "CWD C" ;
		CWDC:units = "gC/m^2" ;
		CWDC:cell_methods = "time: mean" ;
		CWDC:_FillValue = 1.e+36f ;
		CWDC:missing_value = 1.e+36f ;
	float CWDC_HR(time, lndgrid) ;
		CWDC_HR:long_name = "coarse woody debris C heterotrophic respiration" ;
		CWDC_HR:units = "gC/m^2/s" ;
		CWDC_HR:cell_methods = "time: mean" ;
		CWDC_HR:_FillValue = 1.e+36f ;
		CWDC_HR:missing_value = 1.e+36f ;
	float CWDC_LOSS(time, lndgrid) ;
		CWDC_LOSS:long_name = "coarse woody debris C loss" ;
		CWDC_LOSS:units = "gC/m^2/s" ;
		CWDC_LOSS:cell_methods = "time: mean" ;
		CWDC_LOSS:_FillValue = 1.e+36f ;
		CWDC_LOSS:missing_value = 1.e+36f ;
	float CWDC_TO_LITR2C(time, lndgrid) ;
		CWDC_TO_LITR2C:long_name = "decomp. of coarse woody debris C to litter 2 C" ;
		CWDC_TO_LITR2C:units = "gC/m^2/s" ;
		CWDC_TO_LITR2C:cell_methods = "time: mean" ;
		CWDC_TO_LITR2C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR2C:missing_value = 1.e+36f ;
	float CWDC_TO_LITR3C(time, lndgrid) ;
		CWDC_TO_LITR3C:long_name = "decomp. of coarse woody debris C to litter 3 C" ;
		CWDC_TO_LITR3C:units = "gC/m^2/s" ;
		CWDC_TO_LITR3C:cell_methods = "time: mean" ;
		CWDC_TO_LITR3C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR3C:missing_value = 1.e+36f ;
	float CWDC_vr(time, levdcmp, lndgrid) ;
		CWDC_vr:long_name = "CWD C (vertically resolved)" ;
		CWDC_vr:units = "gC/m^3" ;
		CWDC_vr:cell_methods = "time: mean" ;
		CWDC_vr:_FillValue = 1.e+36f ;
		CWDC_vr:missing_value = 1.e+36f ;
	float CWDN(time, lndgrid) ;
		CWDN:long_name = "CWD N" ;
		CWDN:units = "gN/m^2" ;
		CWDN:cell_methods = "time: mean" ;
		CWDN:_FillValue = 1.e+36f ;
		CWDN:missing_value = 1.e+36f ;
	float CWDN_TO_LITR2N(time, lndgrid) ;
		CWDN_TO_LITR2N:long_name = "decomp. of coarse woody debris N to litter 2 N" ;
		CWDN_TO_LITR2N:units = "gN/m^2" ;
		CWDN_TO_LITR2N:cell_methods = "time: mean" ;
		CWDN_TO_LITR2N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR2N:missing_value = 1.e+36f ;
	float CWDN_TO_LITR3N(time, lndgrid) ;
		CWDN_TO_LITR3N:long_name = "decomp. of coarse woody debris N to litter 3 N" ;
		CWDN_TO_LITR3N:units = "gN/m^2" ;
		CWDN_TO_LITR3N:cell_methods = "time: mean" ;
		CWDN_TO_LITR3N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR3N:missing_value = 1.e+36f ;
	float CWDN_vr(time, levdcmp, lndgrid) ;
		CWDN_vr:long_name = "CWD N (vertically resolved)" ;
		CWDN_vr:units = "gN/m^3" ;
		CWDN_vr:cell_methods = "time: mean" ;
		CWDN_vr:_FillValue = 1.e+36f ;
		CWDN_vr:missing_value = 1.e+36f ;
	float DEADCROOTC(time, lndgrid) ;
		DEADCROOTC:long_name = "dead coarse root C" ;
		DEADCROOTC:units = "gC/m^2" ;
		DEADCROOTC:cell_methods = "time: mean" ;
		DEADCROOTC:_FillValue = 1.e+36f ;
		DEADCROOTC:missing_value = 1.e+36f ;
	float DEADCROOTN(time, lndgrid) ;
		DEADCROOTN:long_name = "dead coarse root N" ;
		DEADCROOTN:units = "gN/m^2" ;
		DEADCROOTN:cell_methods = "time: mean" ;
		DEADCROOTN:_FillValue = 1.e+36f ;
		DEADCROOTN:missing_value = 1.e+36f ;
	float DEADSTEMC(time, lndgrid) ;
		DEADSTEMC:long_name = "dead stem C" ;
		DEADSTEMC:units = "gC/m^2" ;
		DEADSTEMC:cell_methods = "time: mean" ;
		DEADSTEMC:_FillValue = 1.e+36f ;
		DEADSTEMC:missing_value = 1.e+36f ;
	float DEADSTEMN(time, lndgrid) ;
		DEADSTEMN:long_name = "dead stem N" ;
		DEADSTEMN:units = "gN/m^2" ;
		DEADSTEMN:cell_methods = "time: mean" ;
		DEADSTEMN:_FillValue = 1.e+36f ;
		DEADSTEMN:missing_value = 1.e+36f ;
	float DENIT(time, lndgrid) ;
		DENIT:long_name = "total rate of denitrification" ;
		DENIT:units = "gN/m^2/s" ;
		DENIT:cell_methods = "time: mean" ;
		DENIT:_FillValue = 1.e+36f ;
		DENIT:missing_value = 1.e+36f ;
	float DISPVEGC(time, lndgrid) ;
		DISPVEGC:long_name = "displayed veg carbon, excluding storage and cpool" ;
		DISPVEGC:units = "gC/m^2" ;
		DISPVEGC:cell_methods = "time: mean" ;
		DISPVEGC:_FillValue = 1.e+36f ;
		DISPVEGC:missing_value = 1.e+36f ;
	float DISPVEGN(time, lndgrid) ;
		DISPVEGN:long_name = "displayed vegetation nitrogen" ;
		DISPVEGN:units = "gN/m^2" ;
		DISPVEGN:cell_methods = "time: mean" ;
		DISPVEGN:_FillValue = 1.e+36f ;
		DISPVEGN:missing_value = 1.e+36f ;
	float DSTDEP(time, lndgrid) ;
		DSTDEP:long_name = "total dust deposition (dry+wet) from atmosphere" ;
		DSTDEP:units = "kg/m^2/s" ;
		DSTDEP:cell_methods = "time: mean" ;
		DSTDEP:_FillValue = 1.e+36f ;
		DSTDEP:missing_value = 1.e+36f ;
	float DSTFLXT(time, lndgrid) ;
		DSTFLXT:long_name = "total surface dust emission" ;
		DSTFLXT:units = "kg/m2/s" ;
		DSTFLXT:cell_methods = "time: mean" ;
		DSTFLXT:_FillValue = 1.e+36f ;
		DSTFLXT:missing_value = 1.e+36f ;
	float DWT_CLOSS(time, lndgrid) ;
		DWT_CLOSS:long_name = "total carbon loss from land cover conversion" ;
		DWT_CLOSS:units = "gC/m^2/s" ;
		DWT_CLOSS:cell_methods = "time: mean" ;
		DWT_CLOSS:_FillValue = 1.e+36f ;
		DWT_CLOSS:missing_value = 1.e+36f ;
	float DWT_CONV_CFLUX(time, lndgrid) ;
		DWT_CONV_CFLUX:long_name = "conversion C flux (immediate loss to atm)" ;
		DWT_CONV_CFLUX:units = "gC/m^2/s" ;
		DWT_CONV_CFLUX:cell_methods = "time: mean" ;
		DWT_CONV_CFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_CFLUX:missing_value = 1.e+36f ;
	float DWT_CONV_NFLUX(time, lndgrid) ;
		DWT_CONV_NFLUX:long_name = "conversion N flux (immediate loss to atm)" ;
		DWT_CONV_NFLUX:units = "gN/m^2/s" ;
		DWT_CONV_NFLUX:cell_methods = "time: mean" ;
		DWT_CONV_NFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_NFLUX:missing_value = 1.e+36f ;
	float DWT_NLOSS(time, lndgrid) ;
		DWT_NLOSS:long_name = "total nitrogen loss from landcover conversion" ;
		DWT_NLOSS:units = "gN/m^2/s" ;
		DWT_NLOSS:cell_methods = "time: mean" ;
		DWT_NLOSS:_FillValue = 1.e+36f ;
		DWT_NLOSS:missing_value = 1.e+36f ;
	float DWT_PROD100C_GAIN(time, lndgrid) ;
		DWT_PROD100C_GAIN:long_name = "landcover change-driven addition to 100-yr wood product pool" ;
		DWT_PROD100C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD100C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD100N_GAIN(time, lndgrid) ;
		DWT_PROD100N_GAIN:long_name = "addition to 100-yr wood product pool" ;
		DWT_PROD100N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD100N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100N_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10C_GAIN(time, lndgrid) ;
		DWT_PROD10C_GAIN:long_name = "landcover change-driven addition to 10-yr wood product pool" ;
		DWT_PROD10C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD10C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10N_GAIN(time, lndgrid) ;
		DWT_PROD10N_GAIN:long_name = "addition to 10-yr wood product pool" ;
		DWT_PROD10N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD10N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10N_GAIN:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDC_TO_DEADSTEM:long_name = "seed source to patch-level deadstem" ;
		DWT_SEEDC_TO_DEADSTEM:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_LEAF(time, lndgrid) ;
		DWT_SEEDC_TO_LEAF:long_name = "seed source to patch-level leaf" ;
		DWT_SEEDC_TO_LEAF:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_LEAF:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDN_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDN_TO_DEADSTEM:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_LEAF(time, lndgrid) ;
		DWT_SEEDN_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDN_TO_LEAF:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_LEAF:missing_value = 1.e+36f ;
	float EFLX_DYNBAL(time, lndgrid) ;
		EFLX_DYNBAL:long_name = "dynamic land cover change conversion energy flux" ;
		EFLX_DYNBAL:units = "W/m^2" ;
		EFLX_DYNBAL:cell_methods = "time: mean" ;
		EFLX_DYNBAL:_FillValue = 1.e+36f ;
		EFLX_DYNBAL:missing_value = 1.e+36f ;
	float EFLX_GRND_LAKE(time, lndgrid) ;
		EFLX_GRND_LAKE:long_name = "net heat flux into lake/snow surface, excluding light transmission" ;
		EFLX_GRND_LAKE:units = "W/m^2" ;
		EFLX_GRND_LAKE:cell_methods = "time: mean" ;
		EFLX_GRND_LAKE:_FillValue = 1.e+36f ;
		EFLX_GRND_LAKE:missing_value = 1.e+36f ;
	float EFLX_LH_TOT(time, lndgrid) ;
		EFLX_LH_TOT:long_name = "total latent heat flux [+ to atm]" ;
		EFLX_LH_TOT:units = "W/m^2" ;
		EFLX_LH_TOT:cell_methods = "time: mean" ;
		EFLX_LH_TOT:_FillValue = 1.e+36f ;
		EFLX_LH_TOT:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_R(time, lndgrid) ;
		EFLX_LH_TOT_R:long_name = "Rural total evaporation" ;
		EFLX_LH_TOT_R:units = "W/m^2" ;
		EFLX_LH_TOT_R:cell_methods = "time: mean" ;
		EFLX_LH_TOT_R:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_R:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_U(time, lndgrid) ;
		EFLX_LH_TOT_U:long_name = "Urban total evaporation" ;
		EFLX_LH_TOT_U:units = "W/m^2" ;
		EFLX_LH_TOT_U:cell_methods = "time: mean" ;
		EFLX_LH_TOT_U:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_U:missing_value = 1.e+36f ;
	float ELAI(time, lndgrid) ;
		ELAI:long_name = "exposed one-sided leaf area index" ;
		ELAI:units = "m^2/m^2" ;
		ELAI:cell_methods = "time: mean" ;
		ELAI:_FillValue = 1.e+36f ;
		ELAI:missing_value = 1.e+36f ;
	float ER(time, lndgrid) ;
		ER:long_name = "total ecosystem respiration, autotrophic + heterotrophic" ;
		ER:units = "gC/m^2/s" ;
		ER:cell_methods = "time: mean" ;
		ER:_FillValue = 1.e+36f ;
		ER:missing_value = 1.e+36f ;
	float ERRH2O(time, lndgrid) ;
		ERRH2O:long_name = "total water conservation error" ;
		ERRH2O:units = "mm" ;
		ERRH2O:cell_methods = "time: mean" ;
		ERRH2O:_FillValue = 1.e+36f ;
		ERRH2O:missing_value = 1.e+36f ;
	float ERRH2OSNO(time, lndgrid) ;
		ERRH2OSNO:long_name = "imbalance in snow depth (liquid water)" ;
		ERRH2OSNO:units = "mm" ;
		ERRH2OSNO:cell_methods = "time: mean" ;
		ERRH2OSNO:_FillValue = 1.e+36f ;
		ERRH2OSNO:missing_value = 1.e+36f ;
	float ERRSEB(time, lndgrid) ;
		ERRSEB:long_name = "surface energy conservation error" ;
		ERRSEB:units = "W/m^2" ;
		ERRSEB:cell_methods = "time: mean" ;
		ERRSEB:_FillValue = 1.e+36f ;
		ERRSEB:missing_value = 1.e+36f ;
	float ERRSOI(time, lndgrid) ;
		ERRSOI:long_name = "soil/lake energy conservation error" ;
		ERRSOI:units = "W/m^2" ;
		ERRSOI:cell_methods = "time: mean" ;
		ERRSOI:_FillValue = 1.e+36f ;
		ERRSOI:missing_value = 1.e+36f ;
	float ERRSOL(time, lndgrid) ;
		ERRSOL:long_name = "solar radiation conservation error" ;
		ERRSOL:units = "W/m^2" ;
		ERRSOL:cell_methods = "time: mean" ;
		ERRSOL:_FillValue = 1.e+36f ;
		ERRSOL:missing_value = 1.e+36f ;
	float ESAI(time, lndgrid) ;
		ESAI:long_name = "exposed one-sided stem area index" ;
		ESAI:units = "m^2/m^2" ;
		ESAI:cell_methods = "time: mean" ;
		ESAI:_FillValue = 1.e+36f ;
		ESAI:missing_value = 1.e+36f ;
	float FAREA_BURNED(time, lndgrid) ;
		FAREA_BURNED:long_name = "timestep fractional area burned" ;
		FAREA_BURNED:units = "proportion" ;
		FAREA_BURNED:cell_methods = "time: mean" ;
		FAREA_BURNED:_FillValue = 1.e+36f ;
		FAREA_BURNED:missing_value = 1.e+36f ;
	float FCEV(time, lndgrid) ;
		FCEV:long_name = "canopy evaporation" ;
		FCEV:units = "W/m^2" ;
		FCEV:cell_methods = "time: mean" ;
		FCEV:_FillValue = 1.e+36f ;
		FCEV:missing_value = 1.e+36f ;
	float FCH4(time, lndgrid) ;
		FCH4:long_name = "Gridcell surface CH4 flux to atmosphere (+ to atm)" ;
		FCH4:units = "kgC/m2/s" ;
		FCH4:cell_methods = "time: mean" ;
		FCH4:_FillValue = 1.e+36f ;
		FCH4:missing_value = 1.e+36f ;
	float FCH4TOCO2(time, lndgrid) ;
		FCH4TOCO2:long_name = "Gridcell oxidation of CH4 to CO2" ;
		FCH4TOCO2:units = "gC/m2/s" ;
		FCH4TOCO2:cell_methods = "time: mean" ;
		FCH4TOCO2:_FillValue = 1.e+36f ;
		FCH4TOCO2:missing_value = 1.e+36f ;
	float FCH4_DFSAT(time, lndgrid) ;
		FCH4_DFSAT:long_name = "CH4 additional flux due to changing fsat, vegetated landunits only" ;
		FCH4_DFSAT:units = "kgC/m2/s" ;
		FCH4_DFSAT:cell_methods = "time: mean" ;
		FCH4_DFSAT:_FillValue = 1.e+36f ;
		FCH4_DFSAT:missing_value = 1.e+36f ;
	float FCOV(time, lndgrid) ;
		FCOV:long_name = "fractional impermeable area" ;
		FCOV:units = "unitless" ;
		FCOV:cell_methods = "time: mean" ;
		FCOV:_FillValue = 1.e+36f ;
		FCOV:missing_value = 1.e+36f ;
	float FCTR(time, lndgrid) ;
		FCTR:long_name = "canopy transpiration" ;
		FCTR:units = "W/m^2" ;
		FCTR:cell_methods = "time: mean" ;
		FCTR:_FillValue = 1.e+36f ;
		FCTR:missing_value = 1.e+36f ;
	float FGEV(time, lndgrid) ;
		FGEV:long_name = "ground evaporation" ;
		FGEV:units = "W/m^2" ;
		FGEV:cell_methods = "time: mean" ;
		FGEV:_FillValue = 1.e+36f ;
		FGEV:missing_value = 1.e+36f ;
	float FGR(time, lndgrid) ;
		FGR:long_name = "heat flux into soil/snow including snow melt and lake / snow light transmission" ;
		FGR:units = "W/m^2" ;
		FGR:cell_methods = "time: mean" ;
		FGR:_FillValue = 1.e+36f ;
		FGR:missing_value = 1.e+36f ;
	float FGR12(time, lndgrid) ;
		FGR12:long_name = "heat flux between soil layers 1 and 2" ;
		FGR12:units = "W/m^2" ;
		FGR12:cell_methods = "time: mean" ;
		FGR12:_FillValue = 1.e+36f ;
		FGR12:missing_value = 1.e+36f ;
	float FGR_R(time, lndgrid) ;
		FGR_R:long_name = "Rural heat flux into soil/snow including snow melt and snow light transmission" ;
		FGR_R:units = "W/m^2" ;
		FGR_R:cell_methods = "time: mean" ;
		FGR_R:_FillValue = 1.e+36f ;
		FGR_R:missing_value = 1.e+36f ;
	float FGR_U(time, lndgrid) ;
		FGR_U:long_name = "Urban heat flux into soil/snow including snow melt" ;
		FGR_U:units = "W/m^2" ;
		FGR_U:cell_methods = "time: mean" ;
		FGR_U:_FillValue = 1.e+36f ;
		FGR_U:missing_value = 1.e+36f ;
	float FH2OSFC(time, lndgrid) ;
		FH2OSFC:long_name = "fraction of ground covered by surface water" ;
		FH2OSFC:units = "unitless" ;
		FH2OSFC:cell_methods = "time: mean" ;
		FH2OSFC:_FillValue = 1.e+36f ;
		FH2OSFC:missing_value = 1.e+36f ;
	float FINUNDATED(time, lndgrid) ;
		FINUNDATED:long_name = "fractional inundated area of vegetated columns" ;
		FINUNDATED:units = "unitless" ;
		FINUNDATED:cell_methods = "time: mean" ;
		FINUNDATED:_FillValue = 1.e+36f ;
		FINUNDATED:missing_value = 1.e+36f ;
	float FINUNDATED_LAG(time, lndgrid) ;
		FINUNDATED_LAG:long_name = "time-lagged inundated fraction of vegetated columns" ;
		FINUNDATED_LAG:units = "unitless" ;
		FINUNDATED_LAG:cell_methods = "time: mean" ;
		FINUNDATED_LAG:_FillValue = 1.e+36f ;
		FINUNDATED_LAG:missing_value = 1.e+36f ;
	float FIRA(time, lndgrid) ;
		FIRA:long_name = "net infrared (longwave) radiation" ;
		FIRA:units = "W/m^2" ;
		FIRA:cell_methods = "time: mean" ;
		FIRA:_FillValue = 1.e+36f ;
		FIRA:missing_value = 1.e+36f ;
	float FIRA_R(time, lndgrid) ;
		FIRA_R:long_name = "Rural net infrared (longwave) radiation" ;
		FIRA_R:units = "W/m^2" ;
		FIRA_R:cell_methods = "time: mean" ;
		FIRA_R:_FillValue = 1.e+36f ;
		FIRA_R:missing_value = 1.e+36f ;
	float FIRA_U(time, lndgrid) ;
		FIRA_U:long_name = "Urban net infrared (longwave) radiation" ;
		FIRA_U:units = "W/m^2" ;
		FIRA_U:cell_methods = "time: mean" ;
		FIRA_U:_FillValue = 1.e+36f ;
		FIRA_U:missing_value = 1.e+36f ;
	float FIRE(time, lndgrid) ;
		FIRE:long_name = "emitted infrared (longwave) radiation" ;
		FIRE:units = "W/m^2" ;
		FIRE:cell_methods = "time: mean" ;
		FIRE:_FillValue = 1.e+36f ;
		FIRE:missing_value = 1.e+36f ;
	float FIRE_R(time, lndgrid) ;
		FIRE_R:long_name = "Rural emitted infrared (longwave) radiation" ;
		FIRE_R:units = "W/m^2" ;
		FIRE_R:cell_methods = "time: mean" ;
		FIRE_R:_FillValue = 1.e+36f ;
		FIRE_R:missing_value = 1.e+36f ;
	float FIRE_U(time, lndgrid) ;
		FIRE_U:long_name = "Urban emitted infrared (longwave) radiation" ;
		FIRE_U:units = "W/m^2" ;
		FIRE_U:cell_methods = "time: mean" ;
		FIRE_U:_FillValue = 1.e+36f ;
		FIRE_U:missing_value = 1.e+36f ;
	float FLDS(time, lndgrid) ;
		FLDS:long_name = "atmospheric longwave radiation" ;
		FLDS:units = "W/m^2" ;
		FLDS:cell_methods = "time: mean" ;
		FLDS:_FillValue = 1.e+36f ;
		FLDS:missing_value = 1.e+36f ;
	float FPG(time, lndgrid) ;
		FPG:long_name = "fraction of potential gpp" ;
		FPG:units = "proportion" ;
		FPG:cell_methods = "time: mean" ;
		FPG:_FillValue = 1.e+36f ;
		FPG:missing_value = 1.e+36f ;
	float FPI(time, lndgrid) ;
		FPI:long_name = "fraction of potential immobilization" ;
		FPI:units = "proportion" ;
		FPI:cell_methods = "time: mean" ;
		FPI:_FillValue = 1.e+36f ;
		FPI:missing_value = 1.e+36f ;
	float FPI_vr(time, levdcmp, lndgrid) ;
		FPI_vr:long_name = "fraction of potential immobilization" ;
		FPI_vr:units = "proportion" ;
		FPI_vr:cell_methods = "time: mean" ;
		FPI_vr:_FillValue = 1.e+36f ;
		FPI_vr:missing_value = 1.e+36f ;
	float FPSN(time, lndgrid) ;
		FPSN:long_name = "photosynthesis" ;
		FPSN:units = "umol/m2s" ;
		FPSN:cell_methods = "time: mean" ;
		FPSN:_FillValue = 1.e+36f ;
		FPSN:missing_value = 1.e+36f ;
	float FPSN_WC(time, lndgrid) ;
		FPSN_WC:long_name = "Rubisco-limited photosynthesis" ;
		FPSN_WC:units = "umol/m2s" ;
		FPSN_WC:cell_methods = "time: mean" ;
		FPSN_WC:_FillValue = 1.e+36f ;
		FPSN_WC:missing_value = 1.e+36f ;
	float FPSN_WJ(time, lndgrid) ;
		FPSN_WJ:long_name = "RuBP-limited photosynthesis" ;
		FPSN_WJ:units = "umol/m2s" ;
		FPSN_WJ:cell_methods = "time: mean" ;
		FPSN_WJ:_FillValue = 1.e+36f ;
		FPSN_WJ:missing_value = 1.e+36f ;
	float FPSN_WP(time, lndgrid) ;
		FPSN_WP:long_name = "Product-limited photosynthesis" ;
		FPSN_WP:units = "umol/m2s" ;
		FPSN_WP:cell_methods = "time: mean" ;
		FPSN_WP:_FillValue = 1.e+36f ;
		FPSN_WP:missing_value = 1.e+36f ;
	float FROOTC(time, lndgrid) ;
		FROOTC:long_name = "fine root C" ;
		FROOTC:units = "gC/m^2" ;
		FROOTC:cell_methods = "time: mean" ;
		FROOTC:_FillValue = 1.e+36f ;
		FROOTC:missing_value = 1.e+36f ;
	float FROOTC_ALLOC(time, lndgrid) ;
		FROOTC_ALLOC:long_name = "fine root C allocation" ;
		FROOTC_ALLOC:units = "gC/m^2/s" ;
		FROOTC_ALLOC:cell_methods = "time: mean" ;
		FROOTC_ALLOC:_FillValue = 1.e+36f ;
		FROOTC_ALLOC:missing_value = 1.e+36f ;
	float FROOTC_LOSS(time, lndgrid) ;
		FROOTC_LOSS:long_name = "fine root C loss" ;
		FROOTC_LOSS:units = "gC/m^2/s" ;
		FROOTC_LOSS:cell_methods = "time: mean" ;
		FROOTC_LOSS:_FillValue = 1.e+36f ;
		FROOTC_LOSS:missing_value = 1.e+36f ;
	float FROOTN(time, lndgrid) ;
		FROOTN:long_name = "fine root N" ;
		FROOTN:units = "gN/m^2" ;
		FROOTN:cell_methods = "time: mean" ;
		FROOTN:_FillValue = 1.e+36f ;
		FROOTN:missing_value = 1.e+36f ;
	float FROST_TABLE(time, lndgrid) ;
		FROST_TABLE:long_name = "frost table depth (vegetated landunits only)" ;
		FROST_TABLE:units = "m" ;
		FROST_TABLE:cell_methods = "time: mean" ;
		FROST_TABLE:_FillValue = 1.e+36f ;
		FROST_TABLE:missing_value = 1.e+36f ;
	float FSA(time, lndgrid) ;
		FSA:long_name = "absorbed solar radiation" ;
		FSA:units = "W/m^2" ;
		FSA:cell_methods = "time: mean" ;
		FSA:_FillValue = 1.e+36f ;
		FSA:missing_value = 1.e+36f ;
	float FSAT(time, lndgrid) ;
		FSAT:long_name = "fractional area with water table at surface" ;
		FSAT:units = "unitless" ;
		FSAT:cell_methods = "time: mean" ;
		FSAT:_FillValue = 1.e+36f ;
		FSAT:missing_value = 1.e+36f ;
	float FSA_R(time, lndgrid) ;
		FSA_R:long_name = "Rural absorbed solar radiation" ;
		FSA_R:units = "W/m^2" ;
		FSA_R:cell_methods = "time: mean" ;
		FSA_R:_FillValue = 1.e+36f ;
		FSA_R:missing_value = 1.e+36f ;
	float FSA_U(time, lndgrid) ;
		FSA_U:long_name = "Urban absorbed solar radiation" ;
		FSA_U:units = "W/m^2" ;
		FSA_U:cell_methods = "time: mean" ;
		FSA_U:_FillValue = 1.e+36f ;
		FSA_U:missing_value = 1.e+36f ;
	float FSDS(time, lndgrid) ;
		FSDS:long_name = "atmospheric incident solar radiation" ;
		FSDS:units = "W/m^2" ;
		FSDS:cell_methods = "time: mean" ;
		FSDS:_FillValue = 1.e+36f ;
		FSDS:missing_value = 1.e+36f ;
	float FSDSND(time, lndgrid) ;
		FSDSND:long_name = "direct nir incident solar radiation" ;
		FSDSND:units = "W/m^2" ;
		FSDSND:cell_methods = "time: mean" ;
		FSDSND:_FillValue = 1.e+36f ;
		FSDSND:missing_value = 1.e+36f ;
	float FSDSNDLN(time, lndgrid) ;
		FSDSNDLN:long_name = "direct nir incident solar radiation at local noon" ;
		FSDSNDLN:units = "W/m^2" ;
		FSDSNDLN:cell_methods = "time: mean" ;
		FSDSNDLN:_FillValue = 1.e+36f ;
		FSDSNDLN:missing_value = 1.e+36f ;
	float FSDSNI(time, lndgrid) ;
		FSDSNI:long_name = "diffuse nir incident solar radiation" ;
		FSDSNI:units = "W/m^2" ;
		FSDSNI:cell_methods = "time: mean" ;
		FSDSNI:_FillValue = 1.e+36f ;
		FSDSNI:missing_value = 1.e+36f ;
	float FSDSVD(time, lndgrid) ;
		FSDSVD:long_name = "direct vis incident solar radiation" ;
		FSDSVD:units = "W/m^2" ;
		FSDSVD:cell_methods = "time: mean" ;
		FSDSVD:_FillValue = 1.e+36f ;
		FSDSVD:missing_value = 1.e+36f ;
	float FSDSVDLN(time, lndgrid) ;
		FSDSVDLN:long_name = "direct vis incident solar radiation at local noon" ;
		FSDSVDLN:units = "W/m^2" ;
		FSDSVDLN:cell_methods = "time: mean" ;
		FSDSVDLN:_FillValue = 1.e+36f ;
		FSDSVDLN:missing_value = 1.e+36f ;
	float FSDSVI(time, lndgrid) ;
		FSDSVI:long_name = "diffuse vis incident solar radiation" ;
		FSDSVI:units = "W/m^2" ;
		FSDSVI:cell_methods = "time: mean" ;
		FSDSVI:_FillValue = 1.e+36f ;
		FSDSVI:missing_value = 1.e+36f ;
	float FSDSVILN(time, lndgrid) ;
		FSDSVILN:long_name = "diffuse vis incident solar radiation at local noon" ;
		FSDSVILN:units = "W/m^2" ;
		FSDSVILN:cell_methods = "time: mean" ;
		FSDSVILN:_FillValue = 1.e+36f ;
		FSDSVILN:missing_value = 1.e+36f ;
	float FSH(time, lndgrid) ;
		FSH:long_name = "sensible heat" ;
		FSH:units = "W/m^2" ;
		FSH:cell_methods = "time: mean" ;
		FSH:_FillValue = 1.e+36f ;
		FSH:missing_value = 1.e+36f ;
	float FSH_G(time, lndgrid) ;
		FSH_G:long_name = "sensible heat from ground" ;
		FSH_G:units = "W/m^2" ;
		FSH_G:cell_methods = "time: mean" ;
		FSH_G:_FillValue = 1.e+36f ;
		FSH_G:missing_value = 1.e+36f ;
	float FSH_NODYNLNDUSE(time, lndgrid) ;
		FSH_NODYNLNDUSE:long_name = "sensible heat not including correction for land use change" ;
		FSH_NODYNLNDUSE:units = "W/m^2" ;
		FSH_NODYNLNDUSE:cell_methods = "time: mean" ;
		FSH_NODYNLNDUSE:_FillValue = 1.e+36f ;
		FSH_NODYNLNDUSE:missing_value = 1.e+36f ;
	float FSH_R(time, lndgrid) ;
		FSH_R:long_name = "Rural sensible heat" ;
		FSH_R:units = "W/m^2" ;
		FSH_R:cell_methods = "time: mean" ;
		FSH_R:_FillValue = 1.e+36f ;
		FSH_R:missing_value = 1.e+36f ;
	float FSH_U(time, lndgrid) ;
		FSH_U:long_name = "Urban sensible heat" ;
		FSH_U:units = "W/m^2" ;
		FSH_U:cell_methods = "time: mean" ;
		FSH_U:_FillValue = 1.e+36f ;
		FSH_U:missing_value = 1.e+36f ;
	float FSH_V(time, lndgrid) ;
		FSH_V:long_name = "sensible heat from veg" ;
		FSH_V:units = "W/m^2" ;
		FSH_V:cell_methods = "time: mean" ;
		FSH_V:_FillValue = 1.e+36f ;
		FSH_V:missing_value = 1.e+36f ;
	float FSM(time, lndgrid) ;
		FSM:long_name = "snow melt heat flux" ;
		FSM:units = "W/m^2" ;
		FSM:cell_methods = "time: mean" ;
		FSM:_FillValue = 1.e+36f ;
		FSM:missing_value = 1.e+36f ;
	float FSM_R(time, lndgrid) ;
		FSM_R:long_name = "Rural snow melt heat flux" ;
		FSM_R:units = "W/m^2" ;
		FSM_R:cell_methods = "time: mean" ;
		FSM_R:_FillValue = 1.e+36f ;
		FSM_R:missing_value = 1.e+36f ;
	float FSM_U(time, lndgrid) ;
		FSM_U:long_name = "Urban snow melt heat flux" ;
		FSM_U:units = "W/m^2" ;
		FSM_U:cell_methods = "time: mean" ;
		FSM_U:_FillValue = 1.e+36f ;
		FSM_U:missing_value = 1.e+36f ;
	float FSNO(time, lndgrid) ;
		FSNO:long_name = "fraction of ground covered by snow" ;
		FSNO:units = "unitless" ;
		FSNO:cell_methods = "time: mean" ;
		FSNO:_FillValue = 1.e+36f ;
		FSNO:missing_value = 1.e+36f ;
	float FSNO_EFF(time, lndgrid) ;
		FSNO_EFF:long_name = "effective fraction of ground covered by snow" ;
		FSNO_EFF:units = "unitless" ;
		FSNO_EFF:cell_methods = "time: mean" ;
		FSNO_EFF:_FillValue = 1.e+36f ;
		FSNO_EFF:missing_value = 1.e+36f ;
	float FSR(time, lndgrid) ;
		FSR:long_name = "reflected solar radiation" ;
		FSR:units = "W/m^2" ;
		FSR:cell_methods = "time: mean" ;
		FSR:_FillValue = 1.e+36f ;
		FSR:missing_value = 1.e+36f ;
	float FSRND(time, lndgrid) ;
		FSRND:long_name = "direct nir reflected solar radiation" ;
		FSRND:units = "W/m^2" ;
		FSRND:cell_methods = "time: mean" ;
		FSRND:_FillValue = 1.e+36f ;
		FSRND:missing_value = 1.e+36f ;
	float FSRNDLN(time, lndgrid) ;
		FSRNDLN:long_name = "direct nir reflected solar radiation at local noon" ;
		FSRNDLN:units = "W/m^2" ;
		FSRNDLN:cell_methods = "time: mean" ;
		FSRNDLN:_FillValue = 1.e+36f ;
		FSRNDLN:missing_value = 1.e+36f ;
	float FSRNI(time, lndgrid) ;
		FSRNI:long_name = "diffuse nir reflected solar radiation" ;
		FSRNI:units = "W/m^2" ;
		FSRNI:cell_methods = "time: mean" ;
		FSRNI:_FillValue = 1.e+36f ;
		FSRNI:missing_value = 1.e+36f ;
	float FSRVD(time, lndgrid) ;
		FSRVD:long_name = "direct vis reflected solar radiation" ;
		FSRVD:units = "W/m^2" ;
		FSRVD:cell_methods = "time: mean" ;
		FSRVD:_FillValue = 1.e+36f ;
		FSRVD:missing_value = 1.e+36f ;
	float FSRVDLN(time, lndgrid) ;
		FSRVDLN:long_name = "direct vis reflected solar radiation at local noon" ;
		FSRVDLN:units = "W/m^2" ;
		FSRVDLN:cell_methods = "time: mean" ;
		FSRVDLN:_FillValue = 1.e+36f ;
		FSRVDLN:missing_value = 1.e+36f ;
	float FSRVI(time, lndgrid) ;
		FSRVI:long_name = "diffuse vis reflected solar radiation" ;
		FSRVI:units = "W/m^2" ;
		FSRVI:cell_methods = "time: mean" ;
		FSRVI:_FillValue = 1.e+36f ;
		FSRVI:missing_value = 1.e+36f ;
	float FUELC(time, lndgrid) ;
		FUELC:long_name = "fuel load" ;
		FUELC:units = "gC/m^2" ;
		FUELC:cell_methods = "time: mean" ;
		FUELC:_FillValue = 1.e+36f ;
		FUELC:missing_value = 1.e+36f ;
	float F_DENIT(time, lndgrid) ;
		F_DENIT:long_name = "denitrification flux" ;
		F_DENIT:units = "gN/m^2/s" ;
		F_DENIT:cell_methods = "time: mean" ;
		F_DENIT:_FillValue = 1.e+36f ;
		F_DENIT:missing_value = 1.e+36f ;
	float F_DENIT_vr(time, levdcmp, lndgrid) ;
		F_DENIT_vr:long_name = "denitrification flux" ;
		F_DENIT_vr:units = "gN/m^3/s" ;
		F_DENIT_vr:cell_methods = "time: mean" ;
		F_DENIT_vr:_FillValue = 1.e+36f ;
		F_DENIT_vr:missing_value = 1.e+36f ;
	float F_N2O_DENIT(time, lndgrid) ;
		F_N2O_DENIT:long_name = "denitrification N2O flux" ;
		F_N2O_DENIT:units = "gN/m^2/s" ;
		F_N2O_DENIT:cell_methods = "time: mean" ;
		F_N2O_DENIT:_FillValue = 1.e+36f ;
		F_N2O_DENIT:missing_value = 1.e+36f ;
	float F_N2O_NIT(time, lndgrid) ;
		F_N2O_NIT:long_name = "nitrification N2O flux" ;
		F_N2O_NIT:units = "gN/m^2/s" ;
		F_N2O_NIT:cell_methods = "time: mean" ;
		F_N2O_NIT:_FillValue = 1.e+36f ;
		F_N2O_NIT:missing_value = 1.e+36f ;
	float F_NIT(time, lndgrid) ;
		F_NIT:long_name = "nitrification flux" ;
		F_NIT:units = "gN/m^2/s" ;
		F_NIT:cell_methods = "time: mean" ;
		F_NIT:_FillValue = 1.e+36f ;
		F_NIT:missing_value = 1.e+36f ;
	float F_NIT_vr(time, levdcmp, lndgrid) ;
		F_NIT_vr:long_name = "nitrification flux" ;
		F_NIT_vr:units = "gN/m^3/s" ;
		F_NIT_vr:cell_methods = "time: mean" ;
		F_NIT_vr:_FillValue = 1.e+36f ;
		F_NIT_vr:missing_value = 1.e+36f ;
	float GC_HEAT1(time, lndgrid) ;
		GC_HEAT1:long_name = "initial gridcell total heat content" ;
		GC_HEAT1:units = "J/m^2" ;
		GC_HEAT1:cell_methods = "time: mean" ;
		GC_HEAT1:_FillValue = 1.e+36f ;
		GC_HEAT1:missing_value = 1.e+36f ;
	float GC_ICE1(time, lndgrid) ;
		GC_ICE1:long_name = "initial gridcell total ice content" ;
		GC_ICE1:units = "mm" ;
		GC_ICE1:cell_methods = "time: mean" ;
		GC_ICE1:_FillValue = 1.e+36f ;
		GC_ICE1:missing_value = 1.e+36f ;
	float GC_LIQ1(time, lndgrid) ;
		GC_LIQ1:long_name = "initial gridcell total liq content" ;
		GC_LIQ1:units = "mm" ;
		GC_LIQ1:cell_methods = "time: mean" ;
		GC_LIQ1:_FillValue = 1.e+36f ;
		GC_LIQ1:missing_value = 1.e+36f ;
	float GPP(time, lndgrid) ;
		GPP:long_name = "gross primary production" ;
		GPP:units = "gC/m^2/s" ;
		GPP:cell_methods = "time: mean" ;
		GPP:_FillValue = 1.e+36f ;
		GPP:missing_value = 1.e+36f ;
	float GR(time, lndgrid) ;
		GR:long_name = "total growth respiration" ;
		GR:units = "gC/m^2/s" ;
		GR:cell_methods = "time: mean" ;
		GR:_FillValue = 1.e+36f ;
		GR:missing_value = 1.e+36f ;
	float GROSS_NMIN(time, lndgrid) ;
		GROSS_NMIN:long_name = "gross rate of N mineralization" ;
		GROSS_NMIN:units = "gN/m^2/s" ;
		GROSS_NMIN:cell_methods = "time: mean" ;
		GROSS_NMIN:_FillValue = 1.e+36f ;
		GROSS_NMIN:missing_value = 1.e+36f ;
	float H2OCAN(time, lndgrid) ;
		H2OCAN:long_name = "intercepted water" ;
		H2OCAN:units = "mm" ;
		H2OCAN:cell_methods = "time: mean" ;
		H2OCAN:_FillValue = 1.e+36f ;
		H2OCAN:missing_value = 1.e+36f ;
	float H2OSFC(time, lndgrid) ;
		H2OSFC:long_name = "surface water depth" ;
		H2OSFC:units = "mm" ;
		H2OSFC:cell_methods = "time: mean" ;
		H2OSFC:_FillValue = 1.e+36f ;
		H2OSFC:missing_value = 1.e+36f ;
	float H2OSNO(time, lndgrid) ;
		H2OSNO:long_name = "snow depth (liquid water)" ;
		H2OSNO:units = "mm" ;
		H2OSNO:cell_methods = "time: mean" ;
		H2OSNO:_FillValue = 1.e+36f ;
		H2OSNO:missing_value = 1.e+36f ;
	float H2OSNO_TOP(time, lndgrid) ;
		H2OSNO_TOP:long_name = "mass of snow in top snow layer" ;
		H2OSNO_TOP:units = "kg/m2" ;
		H2OSNO_TOP:cell_methods = "time: mean" ;
		H2OSNO_TOP:_FillValue = 1.e+36f ;
		H2OSNO_TOP:missing_value = 1.e+36f ;
	float H2OSOI(time, levgrnd, lndgrid) ;
		H2OSOI:long_name = "volumetric soil water (vegetated landunits only)" ;
		H2OSOI:units = "mm3/mm3" ;
		H2OSOI:cell_methods = "time: mean" ;
		H2OSOI:_FillValue = 1.e+36f ;
		H2OSOI:missing_value = 1.e+36f ;
	float HC(time, lndgrid) ;
		HC:long_name = "heat content of soil/snow/lake" ;
		HC:units = "MJ/m2" ;
		HC:cell_methods = "time: mean" ;
		HC:_FillValue = 1.e+36f ;
		HC:missing_value = 1.e+36f ;
	float HCSOI(time, lndgrid) ;
		HCSOI:long_name = "soil heat content" ;
		HCSOI:units = "MJ/m2" ;
		HCSOI:cell_methods = "time: mean" ;
		HCSOI:_FillValue = 1.e+36f ;
		HCSOI:missing_value = 1.e+36f ;
	float HEAT_FROM_AC(time, lndgrid) ;
		HEAT_FROM_AC:long_name = "sensible heat flux put into canyon due to heat removed from air conditioning" ;
		HEAT_FROM_AC:units = "W/m^2" ;
		HEAT_FROM_AC:cell_methods = "time: mean" ;
		HEAT_FROM_AC:_FillValue = 1.e+36f ;
		HEAT_FROM_AC:missing_value = 1.e+36f ;
	float HR(time, lndgrid) ;
		HR:long_name = "total heterotrophic respiration" ;
		HR:units = "gC/m^2/s" ;
		HR:cell_methods = "time: mean" ;
		HR:_FillValue = 1.e+36f ;
		HR:missing_value = 1.e+36f ;
	float HR_vr(time, levdcmp, lndgrid) ;
		HR_vr:long_name = "total vertically resolved heterotrophic respiration" ;
		HR_vr:units = "gC/m^3/s" ;
		HR_vr:cell_methods = "time: mean" ;
		HR_vr:_FillValue = 1.e+36f ;
		HR_vr:missing_value = 1.e+36f ;
	float HTOP(time, lndgrid) ;
		HTOP:long_name = "canopy top" ;
		HTOP:units = "m" ;
		HTOP:cell_methods = "time: mean" ;
		HTOP:_FillValue = 1.e+36f ;
		HTOP:missing_value = 1.e+36f ;
	float INT_SNOW(time, lndgrid) ;
		INT_SNOW:long_name = "accumulated swe (vegetated landunits only)" ;
		INT_SNOW:units = "mm" ;
		INT_SNOW:cell_methods = "time: mean" ;
		INT_SNOW:_FillValue = 1.e+36f ;
		INT_SNOW:missing_value = 1.e+36f ;
	float LAISHA(time, lndgrid) ;
		LAISHA:long_name = "shaded projected leaf area index" ;
		LAISHA:units = "none" ;
		LAISHA:cell_methods = "time: mean" ;
		LAISHA:_FillValue = 1.e+36f ;
		LAISHA:missing_value = 1.e+36f ;
	float LAISUN(time, lndgrid) ;
		LAISUN:long_name = "sunlit projected leaf area index" ;
		LAISUN:units = "none" ;
		LAISUN:cell_methods = "time: mean" ;
		LAISUN:_FillValue = 1.e+36f ;
		LAISUN:missing_value = 1.e+36f ;
	float LAKEICEFRAC(time, levlak, lndgrid) ;
		LAKEICEFRAC:long_name = "lake layer ice mass fraction" ;
		LAKEICEFRAC:units = "unitless" ;
		LAKEICEFRAC:cell_methods = "time: mean" ;
		LAKEICEFRAC:_FillValue = 1.e+36f ;
		LAKEICEFRAC:missing_value = 1.e+36f ;
	float LAKEICETHICK(time, lndgrid) ;
		LAKEICETHICK:long_name = "thickness of lake ice (including physical expansion on freezing)" ;
		LAKEICETHICK:units = "m" ;
		LAKEICETHICK:cell_methods = "time: mean" ;
		LAKEICETHICK:_FillValue = 1.e+36f ;
		LAKEICETHICK:missing_value = 1.e+36f ;
	float LAND_UPTAKE(time, lndgrid) ;
		LAND_UPTAKE:long_name = "NEE minus LAND_USE_FLUX, negative for update" ;
		LAND_UPTAKE:units = "gC/m^2/s" ;
		LAND_UPTAKE:cell_methods = "time: mean" ;
		LAND_UPTAKE:_FillValue = 1.e+36f ;
		LAND_UPTAKE:missing_value = 1.e+36f ;
	float LAND_USE_FLUX(time, lndgrid) ;
		LAND_USE_FLUX:long_name = "total C emitted from land cover conversion and wood product pools" ;
		LAND_USE_FLUX:units = "gC/m^2/s" ;
		LAND_USE_FLUX:cell_methods = "time: mean" ;
		LAND_USE_FLUX:_FillValue = 1.e+36f ;
		LAND_USE_FLUX:missing_value = 1.e+36f ;
	float LEAFC(time, lndgrid) ;
		LEAFC:long_name = "leaf C" ;
		LEAFC:units = "gC/m^2" ;
		LEAFC:cell_methods = "time: mean" ;
		LEAFC:_FillValue = 1.e+36f ;
		LEAFC:missing_value = 1.e+36f ;
	float LEAFC_ALLOC(time, lndgrid) ;
		LEAFC_ALLOC:long_name = "leaf C allocation" ;
		LEAFC_ALLOC:units = "gC/m^2/s" ;
		LEAFC_ALLOC:cell_methods = "time: mean" ;
		LEAFC_ALLOC:_FillValue = 1.e+36f ;
		LEAFC_ALLOC:missing_value = 1.e+36f ;
	float LEAFC_LOSS(time, lndgrid) ;
		LEAFC_LOSS:long_name = "leaf C loss" ;
		LEAFC_LOSS:units = "gC/m^2/s" ;
		LEAFC_LOSS:cell_methods = "time: mean" ;
		LEAFC_LOSS:_FillValue = 1.e+36f ;
		LEAFC_LOSS:missing_value = 1.e+36f ;
	float LEAFN(time, lndgrid) ;
		LEAFN:long_name = "leaf N" ;
		LEAFN:units = "gN/m^2" ;
		LEAFN:cell_methods = "time: mean" ;
		LEAFN:_FillValue = 1.e+36f ;
		LEAFN:missing_value = 1.e+36f ;
	float LEAF_MR(time, lndgrid) ;
		LEAF_MR:long_name = "leaf maintenance respiration" ;
		LEAF_MR:units = "gC/m^2/s" ;
		LEAF_MR:cell_methods = "time: mean" ;
		LEAF_MR:_FillValue = 1.e+36f ;
		LEAF_MR:missing_value = 1.e+36f ;
	float LFC2(time, lndgrid) ;
		LFC2:long_name = "conversion area fraction of BET and BDT that burned" ;
		LFC2:units = "per sec" ;
		LFC2:cell_methods = "time: mean" ;
		LFC2:_FillValue = 1.e+36f ;
		LFC2:missing_value = 1.e+36f ;
	float LF_CONV_CFLUX(time, lndgrid) ;
		LF_CONV_CFLUX:long_name = "conversion carbon due to BET and BDT area decreasing" ;
		LF_CONV_CFLUX:units = "gC/m^2/s" ;
		LF_CONV_CFLUX:cell_methods = "time: mean" ;
		LF_CONV_CFLUX:_FillValue = 1.e+36f ;
		LF_CONV_CFLUX:missing_value = 1.e+36f ;
	float LITFALL(time, lndgrid) ;
		LITFALL:long_name = "litterfall (leaves and fine roots)" ;
		LITFALL:units = "gC/m^2/s" ;
		LITFALL:cell_methods = "time: mean" ;
		LITFALL:_FillValue = 1.e+36f ;
		LITFALL:missing_value = 1.e+36f ;
	float LITHR(time, lndgrid) ;
		LITHR:long_name = "litter heterotrophic respiration" ;
		LITHR:units = "gC/m^2/s" ;
		LITHR:cell_methods = "time: mean" ;
		LITHR:_FillValue = 1.e+36f ;
		LITHR:missing_value = 1.e+36f ;
	float LITR1C(time, lndgrid) ;
		LITR1C:long_name = "LITR1 C" ;
		LITR1C:units = "gC/m^2" ;
		LITR1C:cell_methods = "time: mean" ;
		LITR1C:_FillValue = 1.e+36f ;
		LITR1C:missing_value = 1.e+36f ;
	float LITR1C_TO_SOIL1C(time, lndgrid) ;
		LITR1C_TO_SOIL1C:long_name = "decomp. of litter 1 C to soil 1 C" ;
		LITR1C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR1C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR1C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR1C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR1C_vr(time, levdcmp, lndgrid) ;
		LITR1C_vr:long_name = "LITR1 C (vertically resolved)" ;
		LITR1C_vr:units = "gC/m^3" ;
		LITR1C_vr:cell_methods = "time: mean" ;
		LITR1C_vr:_FillValue = 1.e+36f ;
		LITR1C_vr:missing_value = 1.e+36f ;
	float LITR1N(time, lndgrid) ;
		LITR1N:long_name = "LITR1 N" ;
		LITR1N:units = "gN/m^2" ;
		LITR1N:cell_methods = "time: mean" ;
		LITR1N:_FillValue = 1.e+36f ;
		LITR1N:missing_value = 1.e+36f ;
	float LITR1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR1N_TNDNCY_VERT_TRANS:long_name = "litter 1 N tendency due to vertical transport" ;
		LITR1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR1N_TO_SOIL1N(time, lndgrid) ;
		LITR1N_TO_SOIL1N:long_name = "decomp. of litter 1 N to soil 1 N" ;
		LITR1N_TO_SOIL1N:units = "gN/m^2" ;
		LITR1N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR1N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR1N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR1N_vr(time, levdcmp, lndgrid) ;
		LITR1N_vr:long_name = "LITR1 N (vertically resolved)" ;
		LITR1N_vr:units = "gN/m^3" ;
		LITR1N_vr:cell_methods = "time: mean" ;
		LITR1N_vr:_FillValue = 1.e+36f ;
		LITR1N_vr:missing_value = 1.e+36f ;
	float LITR1_HR(time, lndgrid) ;
		LITR1_HR:long_name = "Het. Resp. from litter 1" ;
		LITR1_HR:units = "gC/m^2/s" ;
		LITR1_HR:cell_methods = "time: mean" ;
		LITR1_HR:_FillValue = 1.e+36f ;
		LITR1_HR:missing_value = 1.e+36f ;
	float LITR2C(time, lndgrid) ;
		LITR2C:long_name = "LITR2 C" ;
		LITR2C:units = "gC/m^2" ;
		LITR2C:cell_methods = "time: mean" ;
		LITR2C:_FillValue = 1.e+36f ;
		LITR2C:missing_value = 1.e+36f ;
	float LITR2C_TO_SOIL1C(time, lndgrid) ;
		LITR2C_TO_SOIL1C:long_name = "decomp. of litter 2 C to soil 1 C" ;
		LITR2C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR2C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR2C_vr(time, levdcmp, lndgrid) ;
		LITR2C_vr:long_name = "LITR2 C (vertically resolved)" ;
		LITR2C_vr:units = "gC/m^3" ;
		LITR2C_vr:cell_methods = "time: mean" ;
		LITR2C_vr:_FillValue = 1.e+36f ;
		LITR2C_vr:missing_value = 1.e+36f ;
	float LITR2N(time, lndgrid) ;
		LITR2N:long_name = "LITR2 N" ;
		LITR2N:units = "gN/m^2" ;
		LITR2N:cell_methods = "time: mean" ;
		LITR2N:_FillValue = 1.e+36f ;
		LITR2N:missing_value = 1.e+36f ;
	float LITR2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR2N_TNDNCY_VERT_TRANS:long_name = "litter 2 N tendency due to vertical transport" ;
		LITR2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR2N_TO_SOIL1N(time, lndgrid) ;
		LITR2N_TO_SOIL1N:long_name = "decomp. of litter 2 N to soil 1 N" ;
		LITR2N_TO_SOIL1N:units = "gN/m^2" ;
		LITR2N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR2N_vr(time, levdcmp, lndgrid) ;
		LITR2N_vr:long_name = "LITR2 N (vertically resolved)" ;
		LITR2N_vr:units = "gN/m^3" ;
		LITR2N_vr:cell_methods = "time: mean" ;
		LITR2N_vr:_FillValue = 1.e+36f ;
		LITR2N_vr:missing_value = 1.e+36f ;
	float LITR2_HR(time, lndgrid) ;
		LITR2_HR:long_name = "Het. Resp. from litter 2" ;
		LITR2_HR:units = "gC/m^2/s" ;
		LITR2_HR:cell_methods = "time: mean" ;
		LITR2_HR:_FillValue = 1.e+36f ;
		LITR2_HR:missing_value = 1.e+36f ;
	float LITR3C(time, lndgrid) ;
		LITR3C:long_name = "LITR3 C" ;
		LITR3C:units = "gC/m^2" ;
		LITR3C:cell_methods = "time: mean" ;
		LITR3C:_FillValue = 1.e+36f ;
		LITR3C:missing_value = 1.e+36f ;
	float LITR3C_TO_SOIL2C(time, lndgrid) ;
		LITR3C_TO_SOIL2C:long_name = "decomp. of litter 3 C to soil 2 C" ;
		LITR3C_TO_SOIL2C:units = "gC/m^2/s" ;
		LITR3C_TO_SOIL2C:cell_methods = "time: mean" ;
		LITR3C_TO_SOIL2C:_FillValue = 1.e+36f ;
		LITR3C_TO_SOIL2C:missing_value = 1.e+36f ;
	float LITR3C_vr(time, levdcmp, lndgrid) ;
		LITR3C_vr:long_name = "LITR3 C (vertically resolved)" ;
		LITR3C_vr:units = "gC/m^3" ;
		LITR3C_vr:cell_methods = "time: mean" ;
		LITR3C_vr:_FillValue = 1.e+36f ;
		LITR3C_vr:missing_value = 1.e+36f ;
	float LITR3N(time, lndgrid) ;
		LITR3N:long_name = "LITR3 N" ;
		LITR3N:units = "gN/m^2" ;
		LITR3N:cell_methods = "time: mean" ;
		LITR3N:_FillValue = 1.e+36f ;
		LITR3N:missing_value = 1.e+36f ;
	float LITR3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR3N_TNDNCY_VERT_TRANS:long_name = "litter 3 N tendency due to vertical transport" ;
		LITR3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR3N_TO_SOIL2N(time, lndgrid) ;
		LITR3N_TO_SOIL2N:long_name = "decomp. of litter 3 N to soil 2 N" ;
		LITR3N_TO_SOIL2N:units = "gN/m^2" ;
		LITR3N_TO_SOIL2N:cell_methods = "time: mean" ;
		LITR3N_TO_SOIL2N:_FillValue = 1.e+36f ;
		LITR3N_TO_SOIL2N:missing_value = 1.e+36f ;
	float LITR3N_vr(time, levdcmp, lndgrid) ;
		LITR3N_vr:long_name = "LITR3 N (vertically resolved)" ;
		LITR3N_vr:units = "gN/m^3" ;
		LITR3N_vr:cell_methods = "time: mean" ;
		LITR3N_vr:_FillValue = 1.e+36f ;
		LITR3N_vr:missing_value = 1.e+36f ;
	float LITR3_HR(time, lndgrid) ;
		LITR3_HR:long_name = "Het. Resp. from litter 3" ;
		LITR3_HR:units = "gC/m^2/s" ;
		LITR3_HR:cell_methods = "time: mean" ;
		LITR3_HR:_FillValue = 1.e+36f ;
		LITR3_HR:missing_value = 1.e+36f ;
	float LITTERC(time, lndgrid) ;
		LITTERC:long_name = "litter C" ;
		LITTERC:units = "gC/m^2" ;
		LITTERC:cell_methods = "time: mean" ;
		LITTERC:_FillValue = 1.e+36f ;
		LITTERC:missing_value = 1.e+36f ;
	float LITTERC_HR(time, lndgrid) ;
		LITTERC_HR:long_name = "litter C heterotrophic respiration" ;
		LITTERC_HR:units = "gC/m^2/s" ;
		LITTERC_HR:cell_methods = "time: mean" ;
		LITTERC_HR:_FillValue = 1.e+36f ;
		LITTERC_HR:missing_value = 1.e+36f ;
	float LITTERC_LOSS(time, lndgrid) ;
		LITTERC_LOSS:long_name = "litter C loss" ;
		LITTERC_LOSS:units = "gC/m^2/s" ;
		LITTERC_LOSS:cell_methods = "time: mean" ;
		LITTERC_LOSS:_FillValue = 1.e+36f ;
		LITTERC_LOSS:missing_value = 1.e+36f ;
	float LIVECROOTC(time, lndgrid) ;
		LIVECROOTC:long_name = "live coarse root C" ;
		LIVECROOTC:units = "gC/m^2" ;
		LIVECROOTC:cell_methods = "time: mean" ;
		LIVECROOTC:_FillValue = 1.e+36f ;
		LIVECROOTC:missing_value = 1.e+36f ;
	float LIVECROOTN(time, lndgrid) ;
		LIVECROOTN:long_name = "live coarse root N" ;
		LIVECROOTN:units = "gN/m^2" ;
		LIVECROOTN:cell_methods = "time: mean" ;
		LIVECROOTN:_FillValue = 1.e+36f ;
		LIVECROOTN:missing_value = 1.e+36f ;
	float LIVESTEMC(time, lndgrid) ;
		LIVESTEMC:long_name = "live stem C" ;
		LIVESTEMC:units = "gC/m^2" ;
		LIVESTEMC:cell_methods = "time: mean" ;
		LIVESTEMC:_FillValue = 1.e+36f ;
		LIVESTEMC:missing_value = 1.e+36f ;
	float LIVESTEMN(time, lndgrid) ;
		LIVESTEMN:long_name = "live stem N" ;
		LIVESTEMN:units = "gN/m^2" ;
		LIVESTEMN:cell_methods = "time: mean" ;
		LIVESTEMN:_FillValue = 1.e+36f ;
		LIVESTEMN:missing_value = 1.e+36f ;
	float MEG_acetaldehyde(time, lndgrid) ;
		MEG_acetaldehyde:long_name = "MEGAN flux" ;
		MEG_acetaldehyde:units = "kg/m2/sec" ;
		MEG_acetaldehyde:cell_methods = "time: mean" ;
		MEG_acetaldehyde:_FillValue = 1.e+36f ;
		MEG_acetaldehyde:missing_value = 1.e+36f ;
	float MEG_acetic_acid(time, lndgrid) ;
		MEG_acetic_acid:long_name = "MEGAN flux" ;
		MEG_acetic_acid:units = "kg/m2/sec" ;
		MEG_acetic_acid:cell_methods = "time: mean" ;
		MEG_acetic_acid:_FillValue = 1.e+36f ;
		MEG_acetic_acid:missing_value = 1.e+36f ;
	float MEG_acetone(time, lndgrid) ;
		MEG_acetone:long_name = "MEGAN flux" ;
		MEG_acetone:units = "kg/m2/sec" ;
		MEG_acetone:cell_methods = "time: mean" ;
		MEG_acetone:_FillValue = 1.e+36f ;
		MEG_acetone:missing_value = 1.e+36f ;
	float MEG_carene_3(time, lndgrid) ;
		MEG_carene_3:long_name = "MEGAN flux" ;
		MEG_carene_3:units = "kg/m2/sec" ;
		MEG_carene_3:cell_methods = "time: mean" ;
		MEG_carene_3:_FillValue = 1.e+36f ;
		MEG_carene_3:missing_value = 1.e+36f ;
	float MEG_ethanol(time, lndgrid) ;
		MEG_ethanol:long_name = "MEGAN flux" ;
		MEG_ethanol:units = "kg/m2/sec" ;
		MEG_ethanol:cell_methods = "time: mean" ;
		MEG_ethanol:_FillValue = 1.e+36f ;
		MEG_ethanol:missing_value = 1.e+36f ;
	float MEG_formaldehyde(time, lndgrid) ;
		MEG_formaldehyde:long_name = "MEGAN flux" ;
		MEG_formaldehyde:units = "kg/m2/sec" ;
		MEG_formaldehyde:cell_methods = "time: mean" ;
		MEG_formaldehyde:_FillValue = 1.e+36f ;
		MEG_formaldehyde:missing_value = 1.e+36f ;
	float MEG_isoprene(time, lndgrid) ;
		MEG_isoprene:long_name = "MEGAN flux" ;
		MEG_isoprene:units = "kg/m2/sec" ;
		MEG_isoprene:cell_methods = "time: mean" ;
		MEG_isoprene:_FillValue = 1.e+36f ;
		MEG_isoprene:missing_value = 1.e+36f ;
	float MEG_methanol(time, lndgrid) ;
		MEG_methanol:long_name = "MEGAN flux" ;
		MEG_methanol:units = "kg/m2/sec" ;
		MEG_methanol:cell_methods = "time: mean" ;
		MEG_methanol:_FillValue = 1.e+36f ;
		MEG_methanol:missing_value = 1.e+36f ;
	float MEG_pinene_a(time, lndgrid) ;
		MEG_pinene_a:long_name = "MEGAN flux" ;
		MEG_pinene_a:units = "kg/m2/sec" ;
		MEG_pinene_a:cell_methods = "time: mean" ;
		MEG_pinene_a:_FillValue = 1.e+36f ;
		MEG_pinene_a:missing_value = 1.e+36f ;
	float MEG_thujene_a(time, lndgrid) ;
		MEG_thujene_a:long_name = "MEGAN flux" ;
		MEG_thujene_a:units = "kg/m2/sec" ;
		MEG_thujene_a:cell_methods = "time: mean" ;
		MEG_thujene_a:_FillValue = 1.e+36f ;
		MEG_thujene_a:missing_value = 1.e+36f ;
	float MR(time, lndgrid) ;
		MR:long_name = "maintenance respiration" ;
		MR:units = "gC/m^2/s" ;
		MR:cell_methods = "time: mean" ;
		MR:_FillValue = 1.e+36f ;
		MR:missing_value = 1.e+36f ;
	float M_LITR1C_TO_LEACHING(time, lndgrid) ;
		M_LITR1C_TO_LEACHING:long_name = "litter 1 C leaching loss" ;
		M_LITR1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR2C_TO_LEACHING(time, lndgrid) ;
		M_LITR2C_TO_LEACHING:long_name = "litter 2 C leaching loss" ;
		M_LITR2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR3C_TO_LEACHING(time, lndgrid) ;
		M_LITR3C_TO_LEACHING:long_name = "litter 3 C leaching loss" ;
		M_LITR3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR3C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL1C_TO_LEACHING(time, lndgrid) ;
		M_SOIL1C_TO_LEACHING:long_name = "soil 1 C leaching loss" ;
		M_SOIL1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL2C_TO_LEACHING(time, lndgrid) ;
		M_SOIL2C_TO_LEACHING:long_name = "soil 2 C leaching loss" ;
		M_SOIL2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL3C_TO_LEACHING(time, lndgrid) ;
		M_SOIL3C_TO_LEACHING:long_name = "soil 3 C leaching loss" ;
		M_SOIL3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL3C_TO_LEACHING:missing_value = 1.e+36f ;
	float NBP(time, lndgrid) ;
		NBP:long_name = "net biome production, includes fire, landuse, and harvest flux, positive for sink" ;
		NBP:units = "gC/m^2/s" ;
		NBP:cell_methods = "time: mean" ;
		NBP:_FillValue = 1.e+36f ;
		NBP:missing_value = 1.e+36f ;
	float NDEPLOY(time, lndgrid) ;
		NDEPLOY:long_name = "total N deployed in new growth" ;
		NDEPLOY:units = "gN/m^2/s" ;
		NDEPLOY:cell_methods = "time: mean" ;
		NDEPLOY:_FillValue = 1.e+36f ;
		NDEPLOY:missing_value = 1.e+36f ;
	float NDEP_TO_SMINN(time, lndgrid) ;
		NDEP_TO_SMINN:long_name = "atmospheric N deposition to soil mineral N" ;
		NDEP_TO_SMINN:units = "gN/m^2/s" ;
		NDEP_TO_SMINN:cell_methods = "time: mean" ;
		NDEP_TO_SMINN:_FillValue = 1.e+36f ;
		NDEP_TO_SMINN:missing_value = 1.e+36f ;
	float NEE(time, lndgrid) ;
		NEE:long_name = "net ecosystem exchange of carbon, includes fire, landuse, harvest, and hrv_xsmrpool flux, positive for source" ;
		NEE:units = "gC/m^2/s" ;
		NEE:cell_methods = "time: mean" ;
		NEE:_FillValue = 1.e+36f ;
		NEE:missing_value = 1.e+36f ;
	float NEM(time, lndgrid) ;
		NEM:long_name = "Gridcell net adjustment to NEE passed to atm. for methane production" ;
		NEM:units = "gC/m2/s" ;
		NEM:cell_methods = "time: mean" ;
		NEM:_FillValue = 1.e+36f ;
		NEM:missing_value = 1.e+36f ;
	float NEP(time, lndgrid) ;
		NEP:long_name = "net ecosystem production, excludes fire, landuse, and harvest flux, positive for sink" ;
		NEP:units = "gC/m^2/s" ;
		NEP:cell_methods = "time: mean" ;
		NEP:_FillValue = 1.e+36f ;
		NEP:missing_value = 1.e+36f ;
	float NET_NMIN(time, lndgrid) ;
		NET_NMIN:long_name = "net rate of N mineralization" ;
		NET_NMIN:units = "gN/m^2/s" ;
		NET_NMIN:cell_methods = "time: mean" ;
		NET_NMIN:_FillValue = 1.e+36f ;
		NET_NMIN:missing_value = 1.e+36f ;
	float NFIRE(time, lndgrid) ;
		NFIRE:long_name = "fire counts valid only in Reg.C" ;
		NFIRE:units = "counts/km2/sec" ;
		NFIRE:cell_methods = "time: mean" ;
		NFIRE:_FillValue = 1.e+36f ;
		NFIRE:missing_value = 1.e+36f ;
	float NFIX_TO_SMINN(time, lndgrid) ;
		NFIX_TO_SMINN:long_name = "symbiotic/asymbiotic N fixation to soil mineral N" ;
		NFIX_TO_SMINN:units = "gN/m^2/s" ;
		NFIX_TO_SMINN:cell_methods = "time: mean" ;
		NFIX_TO_SMINN:_FillValue = 1.e+36f ;
		NFIX_TO_SMINN:missing_value = 1.e+36f ;
	float NPP(time, lndgrid) ;
		NPP:long_name = "net primary production" ;
		NPP:units = "gC/m^2/s" ;
		NPP:cell_methods = "time: mean" ;
		NPP:_FillValue = 1.e+36f ;
		NPP:missing_value = 1.e+36f ;
	float OCDEP(time, lndgrid) ;
		OCDEP:long_name = "total OC deposition (dry+wet) from atmosphere" ;
		OCDEP:units = "kg/m^2/s" ;
		OCDEP:cell_methods = "time: mean" ;
		OCDEP:_FillValue = 1.e+36f ;
		OCDEP:missing_value = 1.e+36f ;
	float O_SCALAR(time, levdcmp, lndgrid) ;
		O_SCALAR:long_name = "fraction by which decomposition is reduced due to anoxia" ;
		O_SCALAR:units = "unitless" ;
		O_SCALAR:cell_methods = "time: mean" ;
		O_SCALAR:_FillValue = 1.e+36f ;
		O_SCALAR:missing_value = 1.e+36f ;
	float PARVEGLN(time, lndgrid) ;
		PARVEGLN:long_name = "absorbed par by vegetation at local noon" ;
		PARVEGLN:units = "W/m^2" ;
		PARVEGLN:cell_methods = "time: mean" ;
		PARVEGLN:_FillValue = 1.e+36f ;
		PARVEGLN:missing_value = 1.e+36f ;
	float PBOT(time, lndgrid) ;
		PBOT:long_name = "atmospheric pressure" ;
		PBOT:units = "Pa" ;
		PBOT:cell_methods = "time: mean" ;
		PBOT:_FillValue = 1.e+36f ;
		PBOT:missing_value = 1.e+36f ;
	float PCH4(time, lndgrid) ;
		PCH4:long_name = "atmospheric partial pressure of CH4" ;
		PCH4:units = "Pa" ;
		PCH4:cell_methods = "time: mean" ;
		PCH4:_FillValue = 1.e+36f ;
		PCH4:missing_value = 1.e+36f ;
	float PCO2(time, lndgrid) ;
		PCO2:long_name = "atmospheric partial pressure of CO2" ;
		PCO2:units = "Pa" ;
		PCO2:cell_methods = "time: mean" ;
		PCO2:_FillValue = 1.e+36f ;
		PCO2:missing_value = 1.e+36f ;
	float PCT_LANDUNIT(time, ltype, lndgrid) ;
		PCT_LANDUNIT:long_name = "% of each landunit on grid cell" ;
		PCT_LANDUNIT:units = "%" ;
		PCT_LANDUNIT:cell_methods = "time: mean" ;
		PCT_LANDUNIT:_FillValue = 1.e+36f ;
		PCT_LANDUNIT:missing_value = 1.e+36f ;
	float PCT_NAT_PFT(time, natpft, lndgrid) ;
		PCT_NAT_PFT:long_name = "% of each PFT on the natural vegetation (i.e., soil) landunit" ;
		PCT_NAT_PFT:units = "%" ;
		PCT_NAT_PFT:cell_methods = "time: mean" ;
		PCT_NAT_PFT:_FillValue = 1.e+36f ;
		PCT_NAT_PFT:missing_value = 1.e+36f ;
	float PFT_CTRUNC(time, lndgrid) ;
		PFT_CTRUNC:long_name = "patch-level sink for C truncation" ;
		PFT_CTRUNC:units = "gC/m^2" ;
		PFT_CTRUNC:cell_methods = "time: mean" ;
		PFT_CTRUNC:_FillValue = 1.e+36f ;
		PFT_CTRUNC:missing_value = 1.e+36f ;
	float PFT_FIRE_CLOSS(time, lndgrid) ;
		PFT_FIRE_CLOSS:long_name = "total patch-level fire C loss for non-peat fires outside land-type converted region" ;
		PFT_FIRE_CLOSS:units = "gC/m^2/s" ;
		PFT_FIRE_CLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_CLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_CLOSS:missing_value = 1.e+36f ;
	float PFT_FIRE_NLOSS(time, lndgrid) ;
		PFT_FIRE_NLOSS:long_name = "total pft-level fire N loss" ;
		PFT_FIRE_NLOSS:units = "gN/m^2/s" ;
		PFT_FIRE_NLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_NLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_NLOSS:missing_value = 1.e+36f ;
	float PFT_NTRUNC(time, lndgrid) ;
		PFT_NTRUNC:long_name = "pft-level sink for N truncation" ;
		PFT_NTRUNC:units = "gN/m^2" ;
		PFT_NTRUNC:cell_methods = "time: mean" ;
		PFT_NTRUNC:_FillValue = 1.e+36f ;
		PFT_NTRUNC:missing_value = 1.e+36f ;
	float PLANT_NDEMAND(time, lndgrid) ;
		PLANT_NDEMAND:long_name = "N flux required to support initial GPP" ;
		PLANT_NDEMAND:units = "gN/m^2/s" ;
		PLANT_NDEMAND:cell_methods = "time: mean" ;
		PLANT_NDEMAND:_FillValue = 1.e+36f ;
		PLANT_NDEMAND:missing_value = 1.e+36f ;
	float POTENTIAL_IMMOB(time, lndgrid) ;
		POTENTIAL_IMMOB:long_name = "potential N immobilization" ;
		POTENTIAL_IMMOB:units = "gN/m^2/s" ;
		POTENTIAL_IMMOB:cell_methods = "time: mean" ;
		POTENTIAL_IMMOB:_FillValue = 1.e+36f ;
		POTENTIAL_IMMOB:missing_value = 1.e+36f ;
	float POT_F_DENIT(time, lndgrid) ;
		POT_F_DENIT:long_name = "potential denitrification flux" ;
		POT_F_DENIT:units = "gN/m^2/s" ;
		POT_F_DENIT:cell_methods = "time: mean" ;
		POT_F_DENIT:_FillValue = 1.e+36f ;
		POT_F_DENIT:missing_value = 1.e+36f ;
	float POT_F_NIT(time, lndgrid) ;
		POT_F_NIT:long_name = "potential nitrification flux" ;
		POT_F_NIT:units = "gN/m^2/s" ;
		POT_F_NIT:cell_methods = "time: mean" ;
		POT_F_NIT:_FillValue = 1.e+36f ;
		POT_F_NIT:missing_value = 1.e+36f ;
	float PROD100C(time, lndgrid) ;
		PROD100C:long_name = "100-yr wood product C" ;
		PROD100C:units = "gC/m^2" ;
		PROD100C:cell_methods = "time: mean" ;
		PROD100C:_FillValue = 1.e+36f ;
		PROD100C:missing_value = 1.e+36f ;
	float PROD100C_LOSS(time, lndgrid) ;
		PROD100C_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100C_LOSS:units = "gC/m^2/s" ;
		PROD100C_LOSS:cell_methods = "time: mean" ;
		PROD100C_LOSS:_FillValue = 1.e+36f ;
		PROD100C_LOSS:missing_value = 1.e+36f ;
	float PROD100N(time, lndgrid) ;
		PROD100N:long_name = "100-yr wood product N" ;
		PROD100N:units = "gN/m^2" ;
		PROD100N:cell_methods = "time: mean" ;
		PROD100N:_FillValue = 1.e+36f ;
		PROD100N:missing_value = 1.e+36f ;
	float PROD100N_LOSS(time, lndgrid) ;
		PROD100N_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100N_LOSS:units = "gN/m^2/s" ;
		PROD100N_LOSS:cell_methods = "time: mean" ;
		PROD100N_LOSS:_FillValue = 1.e+36f ;
		PROD100N_LOSS:missing_value = 1.e+36f ;
	float PROD10C(time, lndgrid) ;
		PROD10C:long_name = "10-yr wood product C" ;
		PROD10C:units = "gC/m^2" ;
		PROD10C:cell_methods = "time: mean" ;
		PROD10C:_FillValue = 1.e+36f ;
		PROD10C:missing_value = 1.e+36f ;
	float PROD10C_LOSS(time, lndgrid) ;
		PROD10C_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10C_LOSS:units = "gC/m^2/s" ;
		PROD10C_LOSS:cell_methods = "time: mean" ;
		PROD10C_LOSS:_FillValue = 1.e+36f ;
		PROD10C_LOSS:missing_value = 1.e+36f ;
	float PROD10N(time, lndgrid) ;
		PROD10N:long_name = "10-yr wood product N" ;
		PROD10N:units = "gN/m^2" ;
		PROD10N:cell_methods = "time: mean" ;
		PROD10N:_FillValue = 1.e+36f ;
		PROD10N:missing_value = 1.e+36f ;
	float PROD10N_LOSS(time, lndgrid) ;
		PROD10N_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10N_LOSS:units = "gN/m^2/s" ;
		PROD10N_LOSS:cell_methods = "time: mean" ;
		PROD10N_LOSS:_FillValue = 1.e+36f ;
		PROD10N_LOSS:missing_value = 1.e+36f ;
	float PRODUCT_CLOSS(time, lndgrid) ;
		PRODUCT_CLOSS:long_name = "total carbon loss from wood product pools" ;
		PRODUCT_CLOSS:units = "gC/m^2/s" ;
		PRODUCT_CLOSS:cell_methods = "time: mean" ;
		PRODUCT_CLOSS:_FillValue = 1.e+36f ;
		PRODUCT_CLOSS:missing_value = 1.e+36f ;
	float PRODUCT_NLOSS(time, lndgrid) ;
		PRODUCT_NLOSS:long_name = "total N loss from wood product pools" ;
		PRODUCT_NLOSS:units = "gN/m^2/s" ;
		PRODUCT_NLOSS:cell_methods = "time: mean" ;
		PRODUCT_NLOSS:_FillValue = 1.e+36f ;
		PRODUCT_NLOSS:missing_value = 1.e+36f ;
	float PSNSHA(time, lndgrid) ;
		PSNSHA:long_name = "shaded leaf photosynthesis" ;
		PSNSHA:units = "umolCO2/m^2/s" ;
		PSNSHA:cell_methods = "time: mean" ;
		PSNSHA:_FillValue = 1.e+36f ;
		PSNSHA:missing_value = 1.e+36f ;
	float PSNSHADE_TO_CPOOL(time, lndgrid) ;
		PSNSHADE_TO_CPOOL:long_name = "C fixation from shaded canopy" ;
		PSNSHADE_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSHADE_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSHADE_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSHADE_TO_CPOOL:missing_value = 1.e+36f ;
	float PSNSUN(time, lndgrid) ;
		PSNSUN:long_name = "sunlit leaf photosynthesis" ;
		PSNSUN:units = "umolCO2/m^2/s" ;
		PSNSUN:cell_methods = "time: mean" ;
		PSNSUN:_FillValue = 1.e+36f ;
		PSNSUN:missing_value = 1.e+36f ;
	float PSNSUN_TO_CPOOL(time, lndgrid) ;
		PSNSUN_TO_CPOOL:long_name = "C fixation from sunlit canopy" ;
		PSNSUN_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSUN_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSUN_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSUN_TO_CPOOL:missing_value = 1.e+36f ;
	float Q2M(time, lndgrid) ;
		Q2M:long_name = "2m specific humidity" ;
		Q2M:units = "kg/kg" ;
		Q2M:cell_methods = "time: mean" ;
		Q2M:_FillValue = 1.e+36f ;
		Q2M:missing_value = 1.e+36f ;
	float QBOT(time, lndgrid) ;
		QBOT:long_name = "atmospheric specific humidity" ;
		QBOT:units = "kg/kg" ;
		QBOT:cell_methods = "time: mean" ;
		QBOT:_FillValue = 1.e+36f ;
		QBOT:missing_value = 1.e+36f ;
	float QCHARGE(time, lndgrid) ;
		QCHARGE:long_name = "aquifer recharge rate (vegetated landunits only)" ;
		QCHARGE:units = "mm/s" ;
		QCHARGE:cell_methods = "time: mean" ;
		QCHARGE:_FillValue = 1.e+36f ;
		QCHARGE:missing_value = 1.e+36f ;
	float QDRAI(time, lndgrid) ;
		QDRAI:long_name = "sub-surface drainage" ;
		QDRAI:units = "mm/s" ;
		QDRAI:cell_methods = "time: mean" ;
		QDRAI:_FillValue = 1.e+36f ;
		QDRAI:missing_value = 1.e+36f ;
	float QDRAI_PERCH(time, lndgrid) ;
		QDRAI_PERCH:long_name = "perched wt drainage" ;
		QDRAI_PERCH:units = "mm/s" ;
		QDRAI_PERCH:cell_methods = "time: mean" ;
		QDRAI_PERCH:_FillValue = 1.e+36f ;
		QDRAI_PERCH:missing_value = 1.e+36f ;
	float QDRAI_XS(time, lndgrid) ;
		QDRAI_XS:long_name = "saturation excess drainage" ;
		QDRAI_XS:units = "mm/s" ;
		QDRAI_XS:cell_methods = "time: mean" ;
		QDRAI_XS:_FillValue = 1.e+36f ;
		QDRAI_XS:missing_value = 1.e+36f ;
	float QDRIP(time, lndgrid) ;
		QDRIP:long_name = "throughfall" ;
		QDRIP:units = "mm/s" ;
		QDRIP:cell_methods = "time: mean" ;
		QDRIP:_FillValue = 1.e+36f ;
		QDRIP:missing_value = 1.e+36f ;
	float QFLOOD(time, lndgrid) ;
		QFLOOD:long_name = "runoff from river flooding" ;
		QFLOOD:units = "mm/s" ;
		QFLOOD:cell_methods = "time: mean" ;
		QFLOOD:_FillValue = 1.e+36f ;
		QFLOOD:missing_value = 1.e+36f ;
	float QFLX_ICE_DYNBAL(time, lndgrid) ;
		QFLX_ICE_DYNBAL:long_name = "ice dynamic land cover change conversion runoff flux" ;
		QFLX_ICE_DYNBAL:units = "mm/s" ;
		QFLX_ICE_DYNBAL:cell_methods = "time: mean" ;
		QFLX_ICE_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_ICE_DYNBAL:missing_value = 1.e+36f ;
	float QFLX_LIQ_DYNBAL(time, lndgrid) ;
		QFLX_LIQ_DYNBAL:long_name = "liq dynamic land cover change conversion runoff flux" ;
		QFLX_LIQ_DYNBAL:units = "mm/s" ;
		QFLX_LIQ_DYNBAL:cell_methods = "time: mean" ;
		QFLX_LIQ_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_LIQ_DYNBAL:missing_value = 1.e+36f ;
	float QH2OSFC(time, lndgrid) ;
		QH2OSFC:long_name = "surface water runoff" ;
		QH2OSFC:units = "mm/s" ;
		QH2OSFC:cell_methods = "time: mean" ;
		QH2OSFC:_FillValue = 1.e+36f ;
		QH2OSFC:missing_value = 1.e+36f ;
	float QINFL(time, lndgrid) ;
		QINFL:long_name = "infiltration" ;
		QINFL:units = "mm/s" ;
		QINFL:cell_methods = "time: mean" ;
		QINFL:_FillValue = 1.e+36f ;
		QINFL:missing_value = 1.e+36f ;
	float QINTR(time, lndgrid) ;
		QINTR:long_name = "interception" ;
		QINTR:units = "mm/s" ;
		QINTR:cell_methods = "time: mean" ;
		QINTR:_FillValue = 1.e+36f ;
		QINTR:missing_value = 1.e+36f ;
	float QIRRIG(time, lndgrid) ;
		QIRRIG:long_name = "water added through irrigation" ;
		QIRRIG:units = "mm/s" ;
		QIRRIG:cell_methods = "time: mean" ;
		QIRRIG:_FillValue = 1.e+36f ;
		QIRRIG:missing_value = 1.e+36f ;
	float QOVER(time, lndgrid) ;
		QOVER:long_name = "surface runoff" ;
		QOVER:units = "mm/s" ;
		QOVER:cell_methods = "time: mean" ;
		QOVER:_FillValue = 1.e+36f ;
		QOVER:missing_value = 1.e+36f ;
	float QOVER_LAG(time, lndgrid) ;
		QOVER_LAG:long_name = "time-lagged surface runoff for soil columns" ;
		QOVER_LAG:units = "mm/s" ;
		QOVER_LAG:cell_methods = "time: mean" ;
		QOVER_LAG:_FillValue = 1.e+36f ;
		QOVER_LAG:missing_value = 1.e+36f ;
	float QRGWL(time, lndgrid) ;
		QRGWL:long_name = "surface runoff at glaciers (liquid only), wetlands, lakes" ;
		QRGWL:units = "mm/s" ;
		QRGWL:cell_methods = "time: mean" ;
		QRGWL:_FillValue = 1.e+36f ;
		QRGWL:missing_value = 1.e+36f ;
	float QRUNOFF(time, lndgrid) ;
		QRUNOFF:long_name = "total liquid runoff (does not include QSNWCPICE)" ;
		QRUNOFF:units = "mm/s" ;
		QRUNOFF:cell_methods = "time: mean" ;
		QRUNOFF:_FillValue = 1.e+36f ;
		QRUNOFF:missing_value = 1.e+36f ;
	float QRUNOFF_NODYNLNDUSE(time, lndgrid) ;
		QRUNOFF_NODYNLNDUSE:long_name = "total liquid runoff (does not include QSNWCPICE) not including correction for land use change" ;
		QRUNOFF_NODYNLNDUSE:units = "mm/s" ;
		QRUNOFF_NODYNLNDUSE:cell_methods = "time: mean" ;
		QRUNOFF_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QRUNOFF_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QRUNOFF_R(time, lndgrid) ;
		QRUNOFF_R:long_name = "Rural total runoff" ;
		QRUNOFF_R:units = "mm/s" ;
		QRUNOFF_R:cell_methods = "time: mean" ;
		QRUNOFF_R:_FillValue = 1.e+36f ;
		QRUNOFF_R:missing_value = 1.e+36f ;
	float QRUNOFF_U(time, lndgrid) ;
		QRUNOFF_U:long_name = "Urban total runoff" ;
		QRUNOFF_U:units = "mm/s" ;
		QRUNOFF_U:cell_methods = "time: mean" ;
		QRUNOFF_U:_FillValue = 1.e+36f ;
		QRUNOFF_U:missing_value = 1.e+36f ;
	float QSNOMELT(time, lndgrid) ;
		QSNOMELT:long_name = "snow melt" ;
		QSNOMELT:units = "mm/s" ;
		QSNOMELT:cell_methods = "time: mean" ;
		QSNOMELT:_FillValue = 1.e+36f ;
		QSNOMELT:missing_value = 1.e+36f ;
	float QSNWCPICE(time, lndgrid) ;
		QSNWCPICE:long_name = "excess snowfall due to snow capping" ;
		QSNWCPICE:units = "mm/s" ;
		QSNWCPICE:cell_methods = "time: mean" ;
		QSNWCPICE:_FillValue = 1.e+36f ;
		QSNWCPICE:missing_value = 1.e+36f ;
	float QSNWCPICE_NODYNLNDUSE(time, lndgrid) ;
		QSNWCPICE_NODYNLNDUSE:long_name = "excess snowfall due to snow capping not including correction for land use change" ;
		QSNWCPICE_NODYNLNDUSE:units = "mm H2O/s" ;
		QSNWCPICE_NODYNLNDUSE:cell_methods = "time: mean" ;
		QSNWCPICE_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QSNWCPICE_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QSOIL(time, lndgrid) ;
		QSOIL:long_name = "Ground evaporation (soil/snow evaporation + soil/snow sublimation - dew)" ;
		QSOIL:units = "mm/s" ;
		QSOIL:cell_methods = "time: mean" ;
		QSOIL:_FillValue = 1.e+36f ;
		QSOIL:missing_value = 1.e+36f ;
	float QVEGE(time, lndgrid) ;
		QVEGE:long_name = "canopy evaporation" ;
		QVEGE:units = "mm/s" ;
		QVEGE:cell_methods = "time: mean" ;
		QVEGE:_FillValue = 1.e+36f ;
		QVEGE:missing_value = 1.e+36f ;
	float QVEGT(time, lndgrid) ;
		QVEGT:long_name = "canopy transpiration" ;
		QVEGT:units = "mm/s" ;
		QVEGT:cell_methods = "time: mean" ;
		QVEGT:_FillValue = 1.e+36f ;
		QVEGT:missing_value = 1.e+36f ;
	float RAIN(time, lndgrid) ;
		RAIN:long_name = "atmospheric rain" ;
		RAIN:units = "mm/s" ;
		RAIN:cell_methods = "time: mean" ;
		RAIN:_FillValue = 1.e+36f ;
		RAIN:missing_value = 1.e+36f ;
	float RETRANSN(time, lndgrid) ;
		RETRANSN:long_name = "plant pool of retranslocated N" ;
		RETRANSN:units = "gN/m^2" ;
		RETRANSN:cell_methods = "time: mean" ;
		RETRANSN:_FillValue = 1.e+36f ;
		RETRANSN:missing_value = 1.e+36f ;
	float RETRANSN_TO_NPOOL(time, lndgrid) ;
		RETRANSN_TO_NPOOL:long_name = "deployment of retranslocated N" ;
		RETRANSN_TO_NPOOL:units = "gN/m^2/s" ;
		RETRANSN_TO_NPOOL:cell_methods = "time: mean" ;
		RETRANSN_TO_NPOOL:_FillValue = 1.e+36f ;
		RETRANSN_TO_NPOOL:missing_value = 1.e+36f ;
	float RH2M(time, lndgrid) ;
		RH2M:long_name = "2m relative humidity" ;
		RH2M:units = "%" ;
		RH2M:cell_methods = "time: mean" ;
		RH2M:_FillValue = 1.e+36f ;
		RH2M:missing_value = 1.e+36f ;
	float RH2M_R(time, lndgrid) ;
		RH2M_R:long_name = "Rural 2m specific humidity" ;
		RH2M_R:units = "%" ;
		RH2M_R:cell_methods = "time: mean" ;
		RH2M_R:_FillValue = 1.e+36f ;
		RH2M_R:missing_value = 1.e+36f ;
	float RH2M_U(time, lndgrid) ;
		RH2M_U:long_name = "Urban 2m relative humidity" ;
		RH2M_U:units = "%" ;
		RH2M_U:cell_methods = "time: mean" ;
		RH2M_U:_FillValue = 1.e+36f ;
		RH2M_U:missing_value = 1.e+36f ;
	float RR(time, lndgrid) ;
		RR:long_name = "root respiration (fine root MR + total root GR)" ;
		RR:units = "gC/m^2/s" ;
		RR:cell_methods = "time: mean" ;
		RR:_FillValue = 1.e+36f ;
		RR:missing_value = 1.e+36f ;
	float RSCANOPY(time, lndgrid) ;
		RSCANOPY:long_name = "canopy resistance" ;
		RSCANOPY:units = " s m-1" ;
		RSCANOPY:cell_methods = "time: mean" ;
		RSCANOPY:_FillValue = 1.e+36f ;
		RSCANOPY:missing_value = 1.e+36f ;
	float SABG(time, lndgrid) ;
		SABG:long_name = "solar rad absorbed by ground" ;
		SABG:units = "W/m^2" ;
		SABG:cell_methods = "time: mean" ;
		SABG:_FillValue = 1.e+36f ;
		SABG:missing_value = 1.e+36f ;
	float SABG_PEN(time, lndgrid) ;
		SABG_PEN:long_name = "Rural solar rad penetrating top soil or snow layer" ;
		SABG_PEN:units = "watt/m^2" ;
		SABG_PEN:cell_methods = "time: mean" ;
		SABG_PEN:_FillValue = 1.e+36f ;
		SABG_PEN:missing_value = 1.e+36f ;
	float SABV(time, lndgrid) ;
		SABV:long_name = "solar rad absorbed by veg" ;
		SABV:units = "W/m^2" ;
		SABV:cell_methods = "time: mean" ;
		SABV:_FillValue = 1.e+36f ;
		SABV:missing_value = 1.e+36f ;
	float SEEDC(time, lndgrid) ;
		SEEDC:long_name = "pool for seeding new Patches" ;
		SEEDC:units = "gC/m^2" ;
		SEEDC:cell_methods = "time: mean" ;
		SEEDC:_FillValue = 1.e+36f ;
		SEEDC:missing_value = 1.e+36f ;
	float SEEDN(time, lndgrid) ;
		SEEDN:long_name = "pool for seeding new PFTs" ;
		SEEDN:units = "gN/m^2" ;
		SEEDN:cell_methods = "time: mean" ;
		SEEDN:_FillValue = 1.e+36f ;
		SEEDN:missing_value = 1.e+36f ;
	float SMINN(time, lndgrid) ;
		SMINN:long_name = "soil mineral N" ;
		SMINN:units = "gN/m^2" ;
		SMINN:cell_methods = "time: mean" ;
		SMINN:_FillValue = 1.e+36f ;
		SMINN:missing_value = 1.e+36f ;
	float SMINN_TO_NPOOL(time, lndgrid) ;
		SMINN_TO_NPOOL:long_name = "deployment of soil mineral N uptake" ;
		SMINN_TO_NPOOL:units = "gN/m^2/s" ;
		SMINN_TO_NPOOL:cell_methods = "time: mean" ;
		SMINN_TO_NPOOL:_FillValue = 1.e+36f ;
		SMINN_TO_NPOOL:missing_value = 1.e+36f ;
	float SMINN_TO_PLANT(time, lndgrid) ;
		SMINN_TO_PLANT:long_name = "plant uptake of soil mineral N" ;
		SMINN_TO_PLANT:units = "gN/m^2/s" ;
		SMINN_TO_PLANT:cell_methods = "time: mean" ;
		SMINN_TO_PLANT:_FillValue = 1.e+36f ;
		SMINN_TO_PLANT:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L1(time, lndgrid) ;
		SMINN_TO_SOIL1N_L1:long_name = "mineral N flux for decomp. of LITR1to SOIL1" ;
		SMINN_TO_SOIL1N_L1:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L2(time, lndgrid) ;
		SMINN_TO_SOIL1N_L2:long_name = "mineral N flux for decomp. of LITR2to SOIL1" ;
		SMINN_TO_SOIL1N_L2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S2(time, lndgrid) ;
		SMINN_TO_SOIL1N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL1" ;
		SMINN_TO_SOIL1N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S3(time, lndgrid) ;
		SMINN_TO_SOIL1N_S3:long_name = "mineral N flux for decomp. of SOIL3to SOIL1" ;
		SMINN_TO_SOIL1N_S3:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_L3(time, lndgrid) ;
		SMINN_TO_SOIL2N_L3:long_name = "mineral N flux for decomp. of LITR3to SOIL2" ;
		SMINN_TO_SOIL2N_L3:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_L3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_L3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_L3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_S1(time, lndgrid) ;
		SMINN_TO_SOIL2N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL2" ;
		SMINN_TO_SOIL2N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S1(time, lndgrid) ;
		SMINN_TO_SOIL3N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL3" ;
		SMINN_TO_SOIL3N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S2(time, lndgrid) ;
		SMINN_TO_SOIL3N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL3" ;
		SMINN_TO_SOIL3N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S2:missing_value = 1.e+36f ;
	float SMIN_NH4(time, lndgrid) ;
		SMIN_NH4:long_name = "soil mineral NH4" ;
		SMIN_NH4:units = "gN/m^2" ;
		SMIN_NH4:cell_methods = "time: mean" ;
		SMIN_NH4:_FillValue = 1.e+36f ;
		SMIN_NH4:missing_value = 1.e+36f ;
	float SMIN_NH4_vr(time, levdcmp, lndgrid) ;
		SMIN_NH4_vr:long_name = "soil mineral NH4 (vert. res.)" ;
		SMIN_NH4_vr:units = "gN/m^3" ;
		SMIN_NH4_vr:cell_methods = "time: mean" ;
		SMIN_NH4_vr:_FillValue = 1.e+36f ;
		SMIN_NH4_vr:missing_value = 1.e+36f ;
	float SMIN_NO3(time, lndgrid) ;
		SMIN_NO3:long_name = "soil mineral NO3" ;
		SMIN_NO3:units = "gN/m^2" ;
		SMIN_NO3:cell_methods = "time: mean" ;
		SMIN_NO3:_FillValue = 1.e+36f ;
		SMIN_NO3:missing_value = 1.e+36f ;
	float SMIN_NO3_LEACHED(time, lndgrid) ;
		SMIN_NO3_LEACHED:long_name = "soil NO3 pool loss to leaching" ;
		SMIN_NO3_LEACHED:units = "gN/m^2/s" ;
		SMIN_NO3_LEACHED:cell_methods = "time: mean" ;
		SMIN_NO3_LEACHED:_FillValue = 1.e+36f ;
		SMIN_NO3_LEACHED:missing_value = 1.e+36f ;
	float SMIN_NO3_RUNOFF(time, lndgrid) ;
		SMIN_NO3_RUNOFF:long_name = "soil NO3 pool loss to runoff" ;
		SMIN_NO3_RUNOFF:units = "gN/m^2/s" ;
		SMIN_NO3_RUNOFF:cell_methods = "time: mean" ;
		SMIN_NO3_RUNOFF:_FillValue = 1.e+36f ;
		SMIN_NO3_RUNOFF:missing_value = 1.e+36f ;
	float SMIN_NO3_vr(time, levdcmp, lndgrid) ;
		SMIN_NO3_vr:long_name = "soil mineral NO3 (vert. res.)" ;
		SMIN_NO3_vr:units = "gN/m^3" ;
		SMIN_NO3_vr:cell_methods = "time: mean" ;
		SMIN_NO3_vr:_FillValue = 1.e+36f ;
		SMIN_NO3_vr:missing_value = 1.e+36f ;
	float SNOBCMCL(time, lndgrid) ;
		SNOBCMCL:long_name = "mass of BC in snow column" ;
		SNOBCMCL:units = "kg/m2" ;
		SNOBCMCL:cell_methods = "time: mean" ;
		SNOBCMCL:_FillValue = 1.e+36f ;
		SNOBCMCL:missing_value = 1.e+36f ;
	float SNOBCMSL(time, lndgrid) ;
		SNOBCMSL:long_name = "mass of BC in top snow layer" ;
		SNOBCMSL:units = "kg/m2" ;
		SNOBCMSL:cell_methods = "time: mean" ;
		SNOBCMSL:_FillValue = 1.e+36f ;
		SNOBCMSL:missing_value = 1.e+36f ;
	float SNODSTMCL(time, lndgrid) ;
		SNODSTMCL:long_name = "mass of dust in snow column" ;
		SNODSTMCL:units = "kg/m2" ;
		SNODSTMCL:cell_methods = "time: mean" ;
		SNODSTMCL:_FillValue = 1.e+36f ;
		SNODSTMCL:missing_value = 1.e+36f ;
	float SNODSTMSL(time, lndgrid) ;
		SNODSTMSL:long_name = "mass of dust in top snow layer" ;
		SNODSTMSL:units = "kg/m2" ;
		SNODSTMSL:cell_methods = "time: mean" ;
		SNODSTMSL:_FillValue = 1.e+36f ;
		SNODSTMSL:missing_value = 1.e+36f ;
	float SNOINTABS(time, lndgrid) ;
		SNOINTABS:long_name = "Percent of incoming solar absorbed by lower snow layers" ;
		SNOINTABS:units = "%" ;
		SNOINTABS:cell_methods = "time: mean" ;
		SNOINTABS:_FillValue = 1.e+36f ;
		SNOINTABS:missing_value = 1.e+36f ;
	float SNOOCMCL(time, lndgrid) ;
		SNOOCMCL:long_name = "mass of OC in snow column" ;
		SNOOCMCL:units = "kg/m2" ;
		SNOOCMCL:cell_methods = "time: mean" ;
		SNOOCMCL:_FillValue = 1.e+36f ;
		SNOOCMCL:missing_value = 1.e+36f ;
	float SNOOCMSL(time, lndgrid) ;
		SNOOCMSL:long_name = "mass of OC in top snow layer" ;
		SNOOCMSL:units = "kg/m2" ;
		SNOOCMSL:cell_methods = "time: mean" ;
		SNOOCMSL:_FillValue = 1.e+36f ;
		SNOOCMSL:missing_value = 1.e+36f ;
	float SNOW(time, lndgrid) ;
		SNOW:long_name = "atmospheric snow" ;
		SNOW:units = "mm/s" ;
		SNOW:cell_methods = "time: mean" ;
		SNOW:_FillValue = 1.e+36f ;
		SNOW:missing_value = 1.e+36f ;
	float SNOWDP(time, lndgrid) ;
		SNOWDP:long_name = "gridcell mean snow height" ;
		SNOWDP:units = "m" ;
		SNOWDP:cell_methods = "time: mean" ;
		SNOWDP:_FillValue = 1.e+36f ;
		SNOWDP:missing_value = 1.e+36f ;
	float SNOWICE(time, lndgrid) ;
		SNOWICE:long_name = "snow ice" ;
		SNOWICE:units = "kg/m2" ;
		SNOWICE:cell_methods = "time: mean" ;
		SNOWICE:_FillValue = 1.e+36f ;
		SNOWICE:missing_value = 1.e+36f ;
	float SNOWLIQ(time, lndgrid) ;
		SNOWLIQ:long_name = "snow liquid water" ;
		SNOWLIQ:units = "kg/m2" ;
		SNOWLIQ:cell_methods = "time: mean" ;
		SNOWLIQ:_FillValue = 1.e+36f ;
		SNOWLIQ:missing_value = 1.e+36f ;
	float SNOW_DEPTH(time, lndgrid) ;
		SNOW_DEPTH:long_name = "snow height of snow covered area" ;
		SNOW_DEPTH:units = "m" ;
		SNOW_DEPTH:cell_methods = "time: mean" ;
		SNOW_DEPTH:_FillValue = 1.e+36f ;
		SNOW_DEPTH:missing_value = 1.e+36f ;
	float SNOW_SINKS(time, lndgrid) ;
		SNOW_SINKS:long_name = "snow sinks (liquid water)" ;
		SNOW_SINKS:units = "mm/s" ;
		SNOW_SINKS:cell_methods = "time: mean" ;
		SNOW_SINKS:_FillValue = 1.e+36f ;
		SNOW_SINKS:missing_value = 1.e+36f ;
	float SNOW_SOURCES(time, lndgrid) ;
		SNOW_SOURCES:long_name = "snow sources (liquid water)" ;
		SNOW_SOURCES:units = "mm/s" ;
		SNOW_SOURCES:cell_methods = "time: mean" ;
		SNOW_SOURCES:_FillValue = 1.e+36f ;
		SNOW_SOURCES:missing_value = 1.e+36f ;
	float SOIL1C(time, lndgrid) ;
		SOIL1C:long_name = "SOIL1 C" ;
		SOIL1C:units = "gC/m^2" ;
		SOIL1C:cell_methods = "time: mean" ;
		SOIL1C:_FillValue = 1.e+36f ;
		SOIL1C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL2C(time, lndgrid) ;
		SOIL1C_TO_SOIL2C:long_name = "decomp. of soil 1 C to soil 2 C" ;
		SOIL1C_TO_SOIL2C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL2C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL2C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL2C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL3C(time, lndgrid) ;
		SOIL1C_TO_SOIL3C:long_name = "decomp. of soil 1 C to soil 3 C" ;
		SOIL1C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL1C_vr(time, levdcmp, lndgrid) ;
		SOIL1C_vr:long_name = "SOIL1 C (vertically resolved)" ;
		SOIL1C_vr:units = "gC/m^3" ;
		SOIL1C_vr:cell_methods = "time: mean" ;
		SOIL1C_vr:_FillValue = 1.e+36f ;
		SOIL1C_vr:missing_value = 1.e+36f ;
	float SOIL1N(time, lndgrid) ;
		SOIL1N:long_name = "SOIL1 N" ;
		SOIL1N:units = "gN/m^2" ;
		SOIL1N:cell_methods = "time: mean" ;
		SOIL1N:_FillValue = 1.e+36f ;
		SOIL1N:missing_value = 1.e+36f ;
	float SOIL1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL1N_TNDNCY_VERT_TRANS:long_name = "soil 1 N tendency due to vertical transport" ;
		SOIL1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL2N(time, lndgrid) ;
		SOIL1N_TO_SOIL2N:long_name = "decomp. of soil 1 N to soil 2 N" ;
		SOIL1N_TO_SOIL2N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL2N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL2N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL2N:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL3N(time, lndgrid) ;
		SOIL1N_TO_SOIL3N:long_name = "decomp. of soil 1 N to soil 3 N" ;
		SOIL1N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL1N_vr(time, levdcmp, lndgrid) ;
		SOIL1N_vr:long_name = "SOIL1 N (vertically resolved)" ;
		SOIL1N_vr:units = "gN/m^3" ;
		SOIL1N_vr:cell_methods = "time: mean" ;
		SOIL1N_vr:_FillValue = 1.e+36f ;
		SOIL1N_vr:missing_value = 1.e+36f ;
	float SOIL1_HR_S2(time, lndgrid) ;
		SOIL1_HR_S2:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S2:units = "gC/m^2/s" ;
		SOIL1_HR_S2:cell_methods = "time: mean" ;
		SOIL1_HR_S2:_FillValue = 1.e+36f ;
		SOIL1_HR_S2:missing_value = 1.e+36f ;
	float SOIL1_HR_S3(time, lndgrid) ;
		SOIL1_HR_S3:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S3:units = "gC/m^2/s" ;
		SOIL1_HR_S3:cell_methods = "time: mean" ;
		SOIL1_HR_S3:_FillValue = 1.e+36f ;
		SOIL1_HR_S3:missing_value = 1.e+36f ;
	float SOIL2C(time, lndgrid) ;
		SOIL2C:long_name = "SOIL2 C" ;
		SOIL2C:units = "gC/m^2" ;
		SOIL2C:cell_methods = "time: mean" ;
		SOIL2C:_FillValue = 1.e+36f ;
		SOIL2C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL1C(time, lndgrid) ;
		SOIL2C_TO_SOIL1C:long_name = "decomp. of soil 2 C to soil 1 C" ;
		SOIL2C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL3C(time, lndgrid) ;
		SOIL2C_TO_SOIL3C:long_name = "decomp. of soil 2 C to soil 3 C" ;
		SOIL2C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL2C_vr(time, levdcmp, lndgrid) ;
		SOIL2C_vr:long_name = "SOIL2 C (vertically resolved)" ;
		SOIL2C_vr:units = "gC/m^3" ;
		SOIL2C_vr:cell_methods = "time: mean" ;
		SOIL2C_vr:_FillValue = 1.e+36f ;
		SOIL2C_vr:missing_value = 1.e+36f ;
	float SOIL2N(time, lndgrid) ;
		SOIL2N:long_name = "SOIL2 N" ;
		SOIL2N:units = "gN/m^2" ;
		SOIL2N:cell_methods = "time: mean" ;
		SOIL2N:_FillValue = 1.e+36f ;
		SOIL2N:missing_value = 1.e+36f ;
	float SOIL2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL2N_TNDNCY_VERT_TRANS:long_name = "soil 2 N tendency due to vertical transport" ;
		SOIL2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL1N(time, lndgrid) ;
		SOIL2N_TO_SOIL1N:long_name = "decomp. of soil 2 N to soil 1 N" ;
		SOIL2N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL3N(time, lndgrid) ;
		SOIL2N_TO_SOIL3N:long_name = "decomp. of soil 2 N to soil 3 N" ;
		SOIL2N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL2N_vr(time, levdcmp, lndgrid) ;
		SOIL2N_vr:long_name = "SOIL2 N (vertically resolved)" ;
		SOIL2N_vr:units = "gN/m^3" ;
		SOIL2N_vr:cell_methods = "time: mean" ;
		SOIL2N_vr:_FillValue = 1.e+36f ;
		SOIL2N_vr:missing_value = 1.e+36f ;
	float SOIL2_HR_S1(time, lndgrid) ;
		SOIL2_HR_S1:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S1:units = "gC/m^2/s" ;
		SOIL2_HR_S1:cell_methods = "time: mean" ;
		SOIL2_HR_S1:_FillValue = 1.e+36f ;
		SOIL2_HR_S1:missing_value = 1.e+36f ;
	float SOIL2_HR_S3(time, lndgrid) ;
		SOIL2_HR_S3:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S3:units = "gC/m^2/s" ;
		SOIL2_HR_S3:cell_methods = "time: mean" ;
		SOIL2_HR_S3:_FillValue = 1.e+36f ;
		SOIL2_HR_S3:missing_value = 1.e+36f ;
	float SOIL3C(time, lndgrid) ;
		SOIL3C:long_name = "SOIL3 C" ;
		SOIL3C:units = "gC/m^2" ;
		SOIL3C:cell_methods = "time: mean" ;
		SOIL3C:_FillValue = 1.e+36f ;
		SOIL3C:missing_value = 1.e+36f ;
	float SOIL3C_TO_SOIL1C(time, lndgrid) ;
		SOIL3C_TO_SOIL1C:long_name = "decomp. of soil 3 C to soil 1 C" ;
		SOIL3C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL3C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL3C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL3C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL3C_vr(time, levdcmp, lndgrid) ;
		SOIL3C_vr:long_name = "SOIL3 C (vertically resolved)" ;
		SOIL3C_vr:units = "gC/m^3" ;
		SOIL3C_vr:cell_methods = "time: mean" ;
		SOIL3C_vr:_FillValue = 1.e+36f ;
		SOIL3C_vr:missing_value = 1.e+36f ;
	float SOIL3N(time, lndgrid) ;
		SOIL3N:long_name = "SOIL3 N" ;
		SOIL3N:units = "gN/m^2" ;
		SOIL3N:cell_methods = "time: mean" ;
		SOIL3N:_FillValue = 1.e+36f ;
		SOIL3N:missing_value = 1.e+36f ;
	float SOIL3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL3N_TNDNCY_VERT_TRANS:long_name = "soil 3 N tendency due to vertical transport" ;
		SOIL3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL3N_TO_SOIL1N(time, lndgrid) ;
		SOIL3N_TO_SOIL1N:long_name = "decomp. of soil 3 N to soil 1 N" ;
		SOIL3N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL3N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL3N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL3N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL3N_vr(time, levdcmp, lndgrid) ;
		SOIL3N_vr:long_name = "SOIL3 N (vertically resolved)" ;
		SOIL3N_vr:units = "gN/m^3" ;
		SOIL3N_vr:cell_methods = "time: mean" ;
		SOIL3N_vr:_FillValue = 1.e+36f ;
		SOIL3N_vr:missing_value = 1.e+36f ;
	float SOIL3_HR(time, lndgrid) ;
		SOIL3_HR:long_name = "Het. Resp. from soil 3" ;
		SOIL3_HR:units = "gC/m^2/s" ;
		SOIL3_HR:cell_methods = "time: mean" ;
		SOIL3_HR:_FillValue = 1.e+36f ;
		SOIL3_HR:missing_value = 1.e+36f ;
	float SOILC(time, lndgrid) ;
		SOILC:long_name = "soil C" ;
		SOILC:units = "gC/m^2" ;
		SOILC:cell_methods = "time: mean" ;
		SOILC:_FillValue = 1.e+36f ;
		SOILC:missing_value = 1.e+36f ;
	float SOILC_HR(time, lndgrid) ;
		SOILC_HR:long_name = "soil C heterotrophic respiration" ;
		SOILC_HR:units = "gC/m^2/s" ;
		SOILC_HR:cell_methods = "time: mean" ;
		SOILC_HR:_FillValue = 1.e+36f ;
		SOILC_HR:missing_value = 1.e+36f ;
	float SOILC_LOSS(time, lndgrid) ;
		SOILC_LOSS:long_name = "soil C loss" ;
		SOILC_LOSS:units = "gC/m^2/s" ;
		SOILC_LOSS:cell_methods = "time: mean" ;
		SOILC_LOSS:_FillValue = 1.e+36f ;
		SOILC_LOSS:missing_value = 1.e+36f ;
	float SOILICE(time, levgrnd, lndgrid) ;
		SOILICE:long_name = "soil ice (vegetated landunits only)" ;
		SOILICE:units = "kg/m2" ;
		SOILICE:cell_methods = "time: mean" ;
		SOILICE:_FillValue = 1.e+36f ;
		SOILICE:missing_value = 1.e+36f ;
	float SOILLIQ(time, levgrnd, lndgrid) ;
		SOILLIQ:long_name = "soil liquid water (vegetated landunits only)" ;
		SOILLIQ:units = "kg/m2" ;
		SOILLIQ:cell_methods = "time: mean" ;
		SOILLIQ:_FillValue = 1.e+36f ;
		SOILLIQ:missing_value = 1.e+36f ;
	float SOILPSI(time, levgrnd, lndgrid) ;
		SOILPSI:long_name = "soil water potential in each soil layer" ;
		SOILPSI:units = "MPa" ;
		SOILPSI:cell_methods = "time: mean" ;
		SOILPSI:_FillValue = 1.e+36f ;
		SOILPSI:missing_value = 1.e+36f ;
	float SOILWATER_10CM(time, lndgrid) ;
		SOILWATER_10CM:long_name = "soil liquid water + ice in top 10cm of soil (veg landunits only)" ;
		SOILWATER_10CM:units = "kg/m2" ;
		SOILWATER_10CM:cell_methods = "time: mean" ;
		SOILWATER_10CM:_FillValue = 1.e+36f ;
		SOILWATER_10CM:missing_value = 1.e+36f ;
	float SOMC_FIRE(time, lndgrid) ;
		SOMC_FIRE:long_name = "C loss due to peat burning" ;
		SOMC_FIRE:units = "gC/m^2/s" ;
		SOMC_FIRE:cell_methods = "time: mean" ;
		SOMC_FIRE:_FillValue = 1.e+36f ;
		SOMC_FIRE:missing_value = 1.e+36f ;
	float SOMHR(time, lndgrid) ;
		SOMHR:long_name = "soil organic matter heterotrophic respiration" ;
		SOMHR:units = "gC/m^2/s" ;
		SOMHR:cell_methods = "time: mean" ;
		SOMHR:_FillValue = 1.e+36f ;
		SOMHR:missing_value = 1.e+36f ;
	float SOM_C_LEACHED(time, lndgrid) ;
		SOM_C_LEACHED:long_name = "total flux of C from SOM pools due to leaching" ;
		SOM_C_LEACHED:units = "gC/m^2/s" ;
		SOM_C_LEACHED:cell_methods = "time: mean" ;
		SOM_C_LEACHED:_FillValue = 1.e+36f ;
		SOM_C_LEACHED:missing_value = 1.e+36f ;
	float SR(time, lndgrid) ;
		SR:long_name = "total soil respiration (HR + root resp)" ;
		SR:units = "gC/m^2/s" ;
		SR:cell_methods = "time: mean" ;
		SR:_FillValue = 1.e+36f ;
		SR:missing_value = 1.e+36f ;
	float STORVEGC(time, lndgrid) ;
		STORVEGC:long_name = "stored vegetation carbon, excluding cpool" ;
		STORVEGC:units = "gC/m^2" ;
		STORVEGC:cell_methods = "time: mean" ;
		STORVEGC:_FillValue = 1.e+36f ;
		STORVEGC:missing_value = 1.e+36f ;
	float STORVEGN(time, lndgrid) ;
		STORVEGN:long_name = "stored vegetation nitrogen" ;
		STORVEGN:units = "gN/m^2" ;
		STORVEGN:cell_methods = "time: mean" ;
		STORVEGN:_FillValue = 1.e+36f ;
		STORVEGN:missing_value = 1.e+36f ;
	float SUPPLEMENT_TO_SMINN(time, lndgrid) ;
		SUPPLEMENT_TO_SMINN:long_name = "supplemental N supply" ;
		SUPPLEMENT_TO_SMINN:units = "gN/m^2/s" ;
		SUPPLEMENT_TO_SMINN:cell_methods = "time: mean" ;
		SUPPLEMENT_TO_SMINN:_FillValue = 1.e+36f ;
		SUPPLEMENT_TO_SMINN:missing_value = 1.e+36f ;
	float SoilAlpha(time, lndgrid) ;
		SoilAlpha:long_name = "factor limiting ground evap" ;
		SoilAlpha:units = "unitless" ;
		SoilAlpha:cell_methods = "time: mean" ;
		SoilAlpha:_FillValue = 1.e+36f ;
		SoilAlpha:missing_value = 1.e+36f ;
	float SoilAlpha_U(time, lndgrid) ;
		SoilAlpha_U:long_name = "urban factor limiting ground evap" ;
		SoilAlpha_U:units = "unitless" ;
		SoilAlpha_U:cell_methods = "time: mean" ;
		SoilAlpha_U:_FillValue = 1.e+36f ;
		SoilAlpha_U:missing_value = 1.e+36f ;
	float TAUX(time, lndgrid) ;
		TAUX:long_name = "zonal surface stress" ;
		TAUX:units = "kg/m/s^2" ;
		TAUX:cell_methods = "time: mean" ;
		TAUX:_FillValue = 1.e+36f ;
		TAUX:missing_value = 1.e+36f ;
	float TAUY(time, lndgrid) ;
		TAUY:long_name = "meridional surface stress" ;
		TAUY:units = "kg/m/s^2" ;
		TAUY:cell_methods = "time: mean" ;
		TAUY:_FillValue = 1.e+36f ;
		TAUY:missing_value = 1.e+36f ;
	float TBOT(time, lndgrid) ;
		TBOT:long_name = "atmospheric air temperature" ;
		TBOT:units = "K" ;
		TBOT:cell_methods = "time: mean" ;
		TBOT:_FillValue = 1.e+36f ;
		TBOT:missing_value = 1.e+36f ;
	float TBUILD(time, lndgrid) ;
		TBUILD:long_name = "internal urban building temperature" ;
		TBUILD:units = "K" ;
		TBUILD:cell_methods = "time: mean" ;
		TBUILD:_FillValue = 1.e+36f ;
		TBUILD:missing_value = 1.e+36f ;
	float TG(time, lndgrid) ;
		TG:long_name = "ground temperature" ;
		TG:units = "K" ;
		TG:cell_methods = "time: mean" ;
		TG:_FillValue = 1.e+36f ;
		TG:missing_value = 1.e+36f ;
	float TG_R(time, lndgrid) ;
		TG_R:long_name = "Rural ground temperature" ;
		TG_R:units = "K" ;
		TG_R:cell_methods = "time: mean" ;
		TG_R:_FillValue = 1.e+36f ;
		TG_R:missing_value = 1.e+36f ;
	float TG_U(time, lndgrid) ;
		TG_U:long_name = "Urban ground temperature" ;
		TG_U:units = "K" ;
		TG_U:cell_methods = "time: mean" ;
		TG_U:_FillValue = 1.e+36f ;
		TG_U:missing_value = 1.e+36f ;
	float TH2OSFC(time, lndgrid) ;
		TH2OSFC:long_name = "surface water temperature" ;
		TH2OSFC:units = "K" ;
		TH2OSFC:cell_methods = "time: mean" ;
		TH2OSFC:_FillValue = 1.e+36f ;
		TH2OSFC:missing_value = 1.e+36f ;
	float THBOT(time, lndgrid) ;
		THBOT:long_name = "atmospheric air potential temperature" ;
		THBOT:units = "K" ;
		THBOT:cell_methods = "time: mean" ;
		THBOT:_FillValue = 1.e+36f ;
		THBOT:missing_value = 1.e+36f ;
	float TKE1(time, lndgrid) ;
		TKE1:long_name = "top lake level eddy thermal conductivity" ;
		TKE1:units = "W/(mK)" ;
		TKE1:cell_methods = "time: mean" ;
		TKE1:_FillValue = 1.e+36f ;
		TKE1:missing_value = 1.e+36f ;
	float TLAI(time, lndgrid) ;
		TLAI:long_name = "total projected leaf area index" ;
		TLAI:units = "none" ;
		TLAI:cell_methods = "time: mean" ;
		TLAI:_FillValue = 1.e+36f ;
		TLAI:missing_value = 1.e+36f ;
	float TLAKE(time, levlak, lndgrid) ;
		TLAKE:long_name = "lake temperature" ;
		TLAKE:units = "K" ;
		TLAKE:cell_methods = "time: mean" ;
		TLAKE:_FillValue = 1.e+36f ;
		TLAKE:missing_value = 1.e+36f ;
	float TOTCOLC(time, lndgrid) ;
		TOTCOLC:long_name = "total column carbon, incl veg and cpool" ;
		TOTCOLC:units = "gC/m^2" ;
		TOTCOLC:cell_methods = "time: mean" ;
		TOTCOLC:_FillValue = 1.e+36f ;
		TOTCOLC:missing_value = 1.e+36f ;
	float TOTCOLCH4(time, lndgrid) ;
		TOTCOLCH4:long_name = "total belowground CH4, (0 for non-lake special landunits)" ;
		TOTCOLCH4:units = "gC/m2" ;
		TOTCOLCH4:cell_methods = "time: mean" ;
		TOTCOLCH4:_FillValue = 1.e+36f ;
		TOTCOLCH4:missing_value = 1.e+36f ;
	float TOTCOLN(time, lndgrid) ;
		TOTCOLN:long_name = "total column-level N" ;
		TOTCOLN:units = "gN/m^2" ;
		TOTCOLN:cell_methods = "time: mean" ;
		TOTCOLN:_FillValue = 1.e+36f ;
		TOTCOLN:missing_value = 1.e+36f ;
	float TOTECOSYSC(time, lndgrid) ;
		TOTECOSYSC:long_name = "total ecosystem carbon, incl veg but excl cpool" ;
		TOTECOSYSC:units = "gC/m^2" ;
		TOTECOSYSC:cell_methods = "time: mean" ;
		TOTECOSYSC:_FillValue = 1.e+36f ;
		TOTECOSYSC:missing_value = 1.e+36f ;
	float TOTECOSYSN(time, lndgrid) ;
		TOTECOSYSN:long_name = "total ecosystem N" ;
		TOTECOSYSN:units = "gN/m^2" ;
		TOTECOSYSN:cell_methods = "time: mean" ;
		TOTECOSYSN:_FillValue = 1.e+36f ;
		TOTECOSYSN:missing_value = 1.e+36f ;
	float TOTLITC(time, lndgrid) ;
		TOTLITC:long_name = "total litter carbon" ;
		TOTLITC:units = "gC/m^2" ;
		TOTLITC:cell_methods = "time: mean" ;
		TOTLITC:_FillValue = 1.e+36f ;
		TOTLITC:missing_value = 1.e+36f ;
	float TOTLITC_1m(time, lndgrid) ;
		TOTLITC_1m:long_name = "total litter carbon to 1 meter depth" ;
		TOTLITC_1m:units = "gC/m^2" ;
		TOTLITC_1m:cell_methods = "time: mean" ;
		TOTLITC_1m:_FillValue = 1.e+36f ;
		TOTLITC_1m:missing_value = 1.e+36f ;
	float TOTLITN(time, lndgrid) ;
		TOTLITN:long_name = "total litter N" ;
		TOTLITN:units = "gN/m^2" ;
		TOTLITN:cell_methods = "time: mean" ;
		TOTLITN:_FillValue = 1.e+36f ;
		TOTLITN:missing_value = 1.e+36f ;
	float TOTLITN_1m(time, lndgrid) ;
		TOTLITN_1m:long_name = "total litter N to 1 meter" ;
		TOTLITN_1m:units = "gN/m^2" ;
		TOTLITN_1m:cell_methods = "time: mean" ;
		TOTLITN_1m:_FillValue = 1.e+36f ;
		TOTLITN_1m:missing_value = 1.e+36f ;
	float TOTPFTC(time, lndgrid) ;
		TOTPFTC:long_name = "total patch-level carbon, including cpool" ;
		TOTPFTC:units = "gC/m^2" ;
		TOTPFTC:cell_methods = "time: mean" ;
		TOTPFTC:_FillValue = 1.e+36f ;
		TOTPFTC:missing_value = 1.e+36f ;
	float TOTPFTN(time, lndgrid) ;
		TOTPFTN:long_name = "total PFT-level nitrogen" ;
		TOTPFTN:units = "gN/m^2" ;
		TOTPFTN:cell_methods = "time: mean" ;
		TOTPFTN:_FillValue = 1.e+36f ;
		TOTPFTN:missing_value = 1.e+36f ;
	float TOTPRODC(time, lndgrid) ;
		TOTPRODC:long_name = "total wood product C" ;
		TOTPRODC:units = "gC/m^2" ;
		TOTPRODC:cell_methods = "time: mean" ;
		TOTPRODC:_FillValue = 1.e+36f ;
		TOTPRODC:missing_value = 1.e+36f ;
	float TOTPRODN(time, lndgrid) ;
		TOTPRODN:long_name = "total wood product N" ;
		TOTPRODN:units = "gN/m^2" ;
		TOTPRODN:cell_methods = "time: mean" ;
		TOTPRODN:_FillValue = 1.e+36f ;
		TOTPRODN:missing_value = 1.e+36f ;
	float TOTSOMC(time, lndgrid) ;
		TOTSOMC:long_name = "total soil organic matter carbon" ;
		TOTSOMC:units = "gC/m^2" ;
		TOTSOMC:cell_methods = "time: mean" ;
		TOTSOMC:_FillValue = 1.e+36f ;
		TOTSOMC:missing_value = 1.e+36f ;
	float TOTSOMC_1m(time, lndgrid) ;
		TOTSOMC_1m:long_name = "total soil organic matter carbon to 1 meter depth" ;
		TOTSOMC_1m:units = "gC/m^2" ;
		TOTSOMC_1m:cell_methods = "time: mean" ;
		TOTSOMC_1m:_FillValue = 1.e+36f ;
		TOTSOMC_1m:missing_value = 1.e+36f ;
	float TOTSOMN(time, lndgrid) ;
		TOTSOMN:long_name = "total soil organic matter N" ;
		TOTSOMN:units = "gN/m^2" ;
		TOTSOMN:cell_methods = "time: mean" ;
		TOTSOMN:_FillValue = 1.e+36f ;
		TOTSOMN:missing_value = 1.e+36f ;
	float TOTSOMN_1m(time, lndgrid) ;
		TOTSOMN_1m:long_name = "total soil organic matter N to 1 meter" ;
		TOTSOMN_1m:units = "gN/m^2" ;
		TOTSOMN_1m:cell_methods = "time: mean" ;
		TOTSOMN_1m:_FillValue = 1.e+36f ;
		TOTSOMN_1m:missing_value = 1.e+36f ;
	float TOTVEGC(time, lndgrid) ;
		TOTVEGC:long_name = "total vegetation carbon, excluding cpool" ;
		TOTVEGC:units = "gC/m^2" ;
		TOTVEGC:cell_methods = "time: mean" ;
		TOTVEGC:_FillValue = 1.e+36f ;
		TOTVEGC:missing_value = 1.e+36f ;
	float TOTVEGN(time, lndgrid) ;
		TOTVEGN:long_name = "total vegetation nitrogen" ;
		TOTVEGN:units = "gN/m^2" ;
		TOTVEGN:cell_methods = "time: mean" ;
		TOTVEGN:_FillValue = 1.e+36f ;
		TOTVEGN:missing_value = 1.e+36f ;
	float TREFMNAV(time, lndgrid) ;
		TREFMNAV:long_name = "daily minimum of average 2-m temperature" ;
		TREFMNAV:units = "K" ;
		TREFMNAV:cell_methods = "time: mean" ;
		TREFMNAV:_FillValue = 1.e+36f ;
		TREFMNAV:missing_value = 1.e+36f ;
	float TREFMNAV_R(time, lndgrid) ;
		TREFMNAV_R:long_name = "Rural daily minimum of average 2-m temperature" ;
		TREFMNAV_R:units = "K" ;
		TREFMNAV_R:cell_methods = "time: mean" ;
		TREFMNAV_R:_FillValue = 1.e+36f ;
		TREFMNAV_R:missing_value = 1.e+36f ;
	float TREFMNAV_U(time, lndgrid) ;
		TREFMNAV_U:long_name = "Urban daily minimum of average 2-m temperature" ;
		TREFMNAV_U:units = "K" ;
		TREFMNAV_U:cell_methods = "time: mean" ;
		TREFMNAV_U:_FillValue = 1.e+36f ;
		TREFMNAV_U:missing_value = 1.e+36f ;
	float TREFMXAV(time, lndgrid) ;
		TREFMXAV:long_name = "daily maximum of average 2-m temperature" ;
		TREFMXAV:units = "K" ;
		TREFMXAV:cell_methods = "time: mean" ;
		TREFMXAV:_FillValue = 1.e+36f ;
		TREFMXAV:missing_value = 1.e+36f ;
	float TREFMXAV_R(time, lndgrid) ;
		TREFMXAV_R:long_name = "Rural daily maximum of average 2-m temperature" ;
		TREFMXAV_R:units = "K" ;
		TREFMXAV_R:cell_methods = "time: mean" ;
		TREFMXAV_R:_FillValue = 1.e+36f ;
		TREFMXAV_R:missing_value = 1.e+36f ;
	float TREFMXAV_U(time, lndgrid) ;
		TREFMXAV_U:long_name = "Urban daily maximum of average 2-m temperature" ;
		TREFMXAV_U:units = "K" ;
		TREFMXAV_U:cell_methods = "time: mean" ;
		TREFMXAV_U:_FillValue = 1.e+36f ;
		TREFMXAV_U:missing_value = 1.e+36f ;
	float TSA(time, lndgrid) ;
		TSA:long_name = "2m air temperature" ;
		TSA:units = "K" ;
		TSA:cell_methods = "time: mean" ;
		TSA:_FillValue = 1.e+36f ;
		TSA:missing_value = 1.e+36f ;
	float TSAI(time, lndgrid) ;
		TSAI:long_name = "total projected stem area index" ;
		TSAI:units = "none" ;
		TSAI:cell_methods = "time: mean" ;
		TSAI:_FillValue = 1.e+36f ;
		TSAI:missing_value = 1.e+36f ;
	float TSA_R(time, lndgrid) ;
		TSA_R:long_name = "Rural 2m air temperature" ;
		TSA_R:units = "K" ;
		TSA_R:cell_methods = "time: mean" ;
		TSA_R:_FillValue = 1.e+36f ;
		TSA_R:missing_value = 1.e+36f ;
	float TSA_U(time, lndgrid) ;
		TSA_U:long_name = "Urban 2m air temperature" ;
		TSA_U:units = "K" ;
		TSA_U:cell_methods = "time: mean" ;
		TSA_U:_FillValue = 1.e+36f ;
		TSA_U:missing_value = 1.e+36f ;
	float TSOI(time, levgrnd, lndgrid) ;
		TSOI:long_name = "soil temperature (vegetated landunits only)" ;
		TSOI:units = "K" ;
		TSOI:cell_methods = "time: mean" ;
		TSOI:_FillValue = 1.e+36f ;
		TSOI:missing_value = 1.e+36f ;
	float TSOI_10CM(time, lndgrid) ;
		TSOI_10CM:long_name = "soil temperature in top 10cm of soil" ;
		TSOI_10CM:units = "K" ;
		TSOI_10CM:cell_methods = "time: mean" ;
		TSOI_10CM:_FillValue = 1.e+36f ;
		TSOI_10CM:missing_value = 1.e+36f ;
	float TSOI_ICE(time, levgrnd, lndgrid) ;
		TSOI_ICE:long_name = "soil temperature (ice landunits only)" ;
		TSOI_ICE:units = "K" ;
		TSOI_ICE:cell_methods = "time: mean" ;
		TSOI_ICE:_FillValue = 1.e+36f ;
		TSOI_ICE:missing_value = 1.e+36f ;
	float TV(time, lndgrid) ;
		TV:long_name = "vegetation temperature" ;
		TV:units = "K" ;
		TV:cell_methods = "time: mean" ;
		TV:_FillValue = 1.e+36f ;
		TV:missing_value = 1.e+36f ;
	float TWS(time, lndgrid) ;
		TWS:long_name = "total water storage" ;
		TWS:units = "mm" ;
		TWS:cell_methods = "time: mean" ;
		TWS:_FillValue = 1.e+36f ;
		TWS:missing_value = 1.e+36f ;
	float T_SCALAR(time, levdcmp, lndgrid) ;
		T_SCALAR:long_name = "temperature inhibition of decomposition" ;
		T_SCALAR:units = "unitless" ;
		T_SCALAR:cell_methods = "time: mean" ;
		T_SCALAR:_FillValue = 1.e+36f ;
		T_SCALAR:missing_value = 1.e+36f ;
	float U10(time, lndgrid) ;
		U10:long_name = "10-m wind" ;
		U10:units = "m/s" ;
		U10:cell_methods = "time: mean" ;
		U10:_FillValue = 1.e+36f ;
		U10:missing_value = 1.e+36f ;
	float URBAN_AC(time, lndgrid) ;
		URBAN_AC:long_name = "urban air conditioning flux" ;
		URBAN_AC:units = "W/m^2" ;
		URBAN_AC:cell_methods = "time: mean" ;
		URBAN_AC:_FillValue = 1.e+36f ;
		URBAN_AC:missing_value = 1.e+36f ;
	float URBAN_HEAT(time, lndgrid) ;
		URBAN_HEAT:long_name = "urban heating flux" ;
		URBAN_HEAT:units = "W/m^2" ;
		URBAN_HEAT:cell_methods = "time: mean" ;
		URBAN_HEAT:_FillValue = 1.e+36f ;
		URBAN_HEAT:missing_value = 1.e+36f ;
	float VOCFLXT(time, lndgrid) ;
		VOCFLXT:long_name = "total VOC flux into atmosphere" ;
		VOCFLXT:units = "moles/m2/sec" ;
		VOCFLXT:cell_methods = "time: mean" ;
		VOCFLXT:_FillValue = 1.e+36f ;
		VOCFLXT:missing_value = 1.e+36f ;
	float VOLR(time, lndgrid) ;
		VOLR:long_name = "river channel water storage" ;
		VOLR:units = "m3" ;
		VOLR:cell_methods = "time: mean" ;
		VOLR:_FillValue = 1.e+36f ;
		VOLR:missing_value = 1.e+36f ;
	float WA(time, lndgrid) ;
		WA:long_name = "water in the unconfined aquifer (vegetated landunits only)" ;
		WA:units = "mm" ;
		WA:cell_methods = "time: mean" ;
		WA:_FillValue = 1.e+36f ;
		WA:missing_value = 1.e+36f ;
	float WASTEHEAT(time, lndgrid) ;
		WASTEHEAT:long_name = "sensible heat flux from heating/cooling sources of urban waste heat" ;
		WASTEHEAT:units = "W/m^2" ;
		WASTEHEAT:cell_methods = "time: mean" ;
		WASTEHEAT:_FillValue = 1.e+36f ;
		WASTEHEAT:missing_value = 1.e+36f ;
	float WF(time, lndgrid) ;
		WF:long_name = "soil water as frac. of whc for top 0.05 m" ;
		WF:units = "proportion" ;
		WF:cell_methods = "time: mean" ;
		WF:_FillValue = 1.e+36f ;
		WF:missing_value = 1.e+36f ;
	float WIND(time, lndgrid) ;
		WIND:long_name = "atmospheric wind velocity magnitude" ;
		WIND:units = "m/s" ;
		WIND:cell_methods = "time: mean" ;
		WIND:_FillValue = 1.e+36f ;
		WIND:missing_value = 1.e+36f ;
	float WOODC(time, lndgrid) ;
		WOODC:long_name = "wood C" ;
		WOODC:units = "gC/m^2" ;
		WOODC:cell_methods = "time: mean" ;
		WOODC:_FillValue = 1.e+36f ;
		WOODC:missing_value = 1.e+36f ;
	float WOODC_ALLOC(time, lndgrid) ;
		WOODC_ALLOC:long_name = "wood C eallocation" ;
		WOODC_ALLOC:units = "gC/m^2/s" ;
		WOODC_ALLOC:cell_methods = "time: mean" ;
		WOODC_ALLOC:_FillValue = 1.e+36f ;
		WOODC_ALLOC:missing_value = 1.e+36f ;
	float WOODC_LOSS(time, lndgrid) ;
		WOODC_LOSS:long_name = "wood C loss" ;
		WOODC_LOSS:units = "gC/m^2/s" ;
		WOODC_LOSS:cell_methods = "time: mean" ;
		WOODC_LOSS:_FillValue = 1.e+36f ;
		WOODC_LOSS:missing_value = 1.e+36f ;
	float WOOD_HARVESTC(time, lndgrid) ;
		WOOD_HARVESTC:long_name = "wood harvest carbon (to product pools)" ;
		WOOD_HARVESTC:units = "gC/m^2/s" ;
		WOOD_HARVESTC:cell_methods = "time: mean" ;
		WOOD_HARVESTC:_FillValue = 1.e+36f ;
		WOOD_HARVESTC:missing_value = 1.e+36f ;
	float WOOD_HARVESTN(time, lndgrid) ;
		WOOD_HARVESTN:long_name = "wood harvest N (to product pools)" ;
		WOOD_HARVESTN:units = "gN/m^2/s" ;
		WOOD_HARVESTN:cell_methods = "time: mean" ;
		WOOD_HARVESTN:_FillValue = 1.e+36f ;
		WOOD_HARVESTN:missing_value = 1.e+36f ;
	float WTGQ(time, lndgrid) ;
		WTGQ:long_name = "surface tracer conductance" ;
		WTGQ:units = "m/s" ;
		WTGQ:cell_methods = "time: mean" ;
		WTGQ:_FillValue = 1.e+36f ;
		WTGQ:missing_value = 1.e+36f ;
	float W_SCALAR(time, levdcmp, lndgrid) ;
		W_SCALAR:long_name = "Moisture (dryness) inhibition of decomposition" ;
		W_SCALAR:units = "unitless" ;
		W_SCALAR:cell_methods = "time: mean" ;
		W_SCALAR:_FillValue = 1.e+36f ;
		W_SCALAR:missing_value = 1.e+36f ;
	float XSMRPOOL(time, lndgrid) ;
		XSMRPOOL:long_name = "temporary photosynthate C pool" ;
		XSMRPOOL:units = "gC/m^2" ;
		XSMRPOOL:cell_methods = "time: mean" ;
		XSMRPOOL:_FillValue = 1.e+36f ;
		XSMRPOOL:missing_value = 1.e+36f ;
	float XSMRPOOL_RECOVER(time, lndgrid) ;
		XSMRPOOL_RECOVER:long_name = "C flux assigned to recovery of negative xsmrpool" ;
		XSMRPOOL_RECOVER:units = "gC/m^2/s" ;
		XSMRPOOL_RECOVER:cell_methods = "time: mean" ;
		XSMRPOOL_RECOVER:_FillValue = 1.e+36f ;
		XSMRPOOL_RECOVER:missing_value = 1.e+36f ;
	float ZBOT(time, lndgrid) ;
		ZBOT:long_name = "atmospheric reference height" ;
		ZBOT:units = "m" ;
		ZBOT:cell_methods = "time: mean" ;
		ZBOT:_FillValue = 1.e+36f ;
		ZBOT:missing_value = 1.e+36f ;
	float ZWT(time, lndgrid) ;
		ZWT:long_name = "water table depth (vegetated landunits only)" ;
		ZWT:units = "m" ;
		ZWT:cell_methods = "time: mean" ;
		ZWT:_FillValue = 1.e+36f ;
		ZWT:missing_value = 1.e+36f ;
	float ZWT_CH4_UNSAT(time, lndgrid) ;
		ZWT_CH4_UNSAT:long_name = "depth of water table for methane production used in non-inundated area" ;
		ZWT_CH4_UNSAT:units = "m" ;
		ZWT_CH4_UNSAT:cell_methods = "time: mean" ;
		ZWT_CH4_UNSAT:_FillValue = 1.e+36f ;
		ZWT_CH4_UNSAT:missing_value = 1.e+36f ;
	float ZWT_PERCH(time, lndgrid) ;
		ZWT_PERCH:long_name = "perched water table depth (vegetated landunits only)" ;
		ZWT_PERCH:units = "m" ;
		ZWT_PERCH:cell_methods = "time: mean" ;
		ZWT_PERCH:_FillValue = 1.e+36f ;
		ZWT_PERCH:missing_value = 1.e+36f ;
	float o2_decomp_depth_unsat(time, levgrnd, lndgrid) ;
		o2_decomp_depth_unsat:long_name = "o2_decomp_depth_unsat" ;
		o2_decomp_depth_unsat:units = "mol/m3/2" ;
		o2_decomp_depth_unsat:cell_methods = "time: mean" ;
		o2_decomp_depth_unsat:_FillValue = 1.e+36f ;
		o2_decomp_depth_unsat:missing_value = 1.e+36f ;

// global attributes:
		:title = "CLM History file information" ;
		:comment = "NOTE: None of the variables are weighted by land fraction!" ;
		:Conventions = "CF-1.0" ;
		:history = "created on 07/19/16 09:53:11" ;
		:source = "Community Land Model CLM4.0" ;
		:hostname = "userdefined" ;
		:username = "gbisht" ;
		:version = "" ;
		:revision_id = "$Id: histFileMod.F90 42903 2012-12-21 15:32:10Z muszala $" ;
		:case_title = "UNSET" ;
		:case_id = "ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-1" ;
		:Surface_dataset = "surfdata_13x26pt_US-Brw_simyr1850.nc" ;
		:Initial_conditions_dataset = "arbitrary initialization" ;
		:PFT_physiological_constants_dataset = "clm_params.c140423.nc" ;
		:ltype_vegetated_or_bare_soil = 1 ;
		:ltype_crop = 2 ;
		:ltype_landice = 3 ;
		:ltype_landice_multiple_elevation_classes = 4 ;
		:ltype_deep_lake = 5 ;
		:ltype_wetland = 6 ;
		:ltype_urban_tbd = 7 ;
		:ltype_urban_hd = 8 ;
		:ltype_urban_md = 9 ;
		:Time_constant_3Dvars_filename = "./ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-1.clm2.h0.0001-12-01-00000.nc" ;
		:Time_constant_3Dvars = "ZSOI:DZSOI:WATSAT:SUCSAT:BSW:HKSAT:ZLAKE:DZLAKE" ;
data:

 levgrnd = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 levlak = 0.05, 0.6, 2.1, 4.6, 8.1, 12.6, 18.6, 25.6, 34.325, 44.775 ;

 levdcmp = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 time = 1 ;

 mcdate = 11202 ;

 mcsec = 0 ;

 mdcur = 1 ;

 mscur = 0 ;

 nstep = 48 ;

 time_bounds =
  0, 1 ;

 date_written =
  "07/19/16" ;

 time_written =
  "09:53:11" ;

 lon = -156.6089, -156.6089, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6083, -156.6082, -156.608, -156.608, -156.6078, -156.6078, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, 
    -156.6069, -156.6069, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6063, -156.6062, -156.6089, -156.6089, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6083, -156.6082, -156.608, -156.608, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6074, -156.6073, 
    -156.6071, -156.6071, -156.6069, -156.6069, -156.6067, -156.6066, 
    -156.6065, -156.6064, -156.6063, -156.6062, -156.6089, -156.6089, 
    -156.6087, -156.6086, -156.6085, -156.6084, -156.6083, -156.6082, 
    -156.608, -156.608, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6074, -156.6073, -156.6071, -156.6071, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6065, -156.6064, -156.6062, -156.6062, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6082, -156.6082, -156.608, -156.608, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6071, -156.6071, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6062, -156.6062, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6082, -156.6082, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6073, -156.6073, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6067, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6062, -156.6089, -156.6088, 
    -156.6087, -156.6086, -156.6084, -156.6084, -156.6082, -156.6082, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6073, -156.6073, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6064, -156.6064, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6084, -156.6084, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6073, -156.6073, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6064, -156.6064, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6084, -156.6084, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6075, -156.6075, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6061, -156.6089, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6084, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6075, -156.6075, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6066, -156.6066, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6086, -156.6086, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6075, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6066, -156.6066, -156.6064, -156.6063, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6086, -156.6086, 
    -156.6084, -156.6083, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6077, -156.6077, -156.6075, -156.6074, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6068, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6063, -156.6062, -156.6061, -156.6088, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6083, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6077, -156.6077, -156.6075, -156.6074, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6068, -156.6068, 
    -156.6066, -156.6065, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6088, -156.6088, -156.6086, -156.6085, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.6079, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6068, -156.6068, -156.6066, -156.6065, -156.6064, -156.6063, 
    -156.6062, -156.6061 ;

 lat = 71.27904, 71.27901, 71.27903, 71.27901, 71.27901, 71.27903, 71.27901, 
    71.27903, 71.279, 71.27902, 71.27902, 71.279, 71.27899, 71.27901, 
    71.27901, 71.27899, 71.27899, 71.27901, 71.27898, 71.27901, 71.27901, 
    71.27898, 71.27901, 71.27898, 71.27898, 71.279, 71.27911, 71.27908, 
    71.27911, 71.27908, 71.27908, 71.2791, 71.27908, 71.2791, 71.2791, 
    71.27907, 71.27907, 71.27909, 71.27909, 71.27907, 71.27909, 71.27906, 
    71.27906, 71.27908, 71.27906, 71.27908, 71.27905, 71.27908, 71.27908, 
    71.27905, 71.27908, 71.27905, 71.27915, 71.27918, 71.27915, 71.27917, 
    71.27917, 71.27915, 71.27917, 71.27914, 71.27914, 71.27917, 71.27914, 
    71.27917, 71.27916, 71.27914, 71.27914, 71.27916, 71.27914, 71.27916, 
    71.27913, 71.27915, 71.27913, 71.27915, 71.27915, 71.27912, 71.27914, 
    71.27912, 71.27923, 71.27925, 71.27923, 71.27925, 71.27924, 71.27922, 
    71.27922, 71.27924, 71.27921, 71.27924, 71.27921, 71.27924, 71.27924, 
    71.27921, 71.27921, 71.27923, 71.27923, 71.27921, 71.27923, 71.2792, 
    71.27922, 71.2792, 71.27922, 71.2792, 71.27922, 71.27919, 71.27932, 
    71.2793, 71.2793, 71.27932, 71.2793, 71.27932, 71.27931, 71.27929, 
    71.27929, 71.27931, 71.27931, 71.27928, 71.27928, 71.2793, 71.27928, 
    71.2793, 71.27927, 71.2793, 71.27927, 71.2793, 71.2793, 71.27927, 
    71.27929, 71.27927, 71.27927, 71.27929, 71.27937, 71.2794, 71.27937, 
    71.27939, 71.27939, 71.27937, 71.27937, 71.27939, 71.27938, 71.27936, 
    71.27936, 71.27938, 71.27935, 71.27937, 71.27935, 71.27937, 71.27935, 
    71.27937, 71.27934, 71.27937, 71.27937, 71.27934, 71.27937, 71.27934, 
    71.27934, 71.27936, 71.27944, 71.27946, 71.27946, 71.27944, 71.27946, 
    71.27943, 71.27943, 71.27946, 71.27946, 71.27943, 71.27945, 71.27943, 
    71.27943, 71.27945, 71.27942, 71.27944, 71.27942, 71.27944, 71.27942, 
    71.27944, 71.27943, 71.27941, 71.27943, 71.27941, 71.27943, 71.2794, 
    71.27951, 71.27953, 71.27951, 71.27953, 71.27953, 71.27951, 71.2795, 
    71.27953, 71.27953, 71.2795, 71.27953, 71.2795, 71.2795, 71.27952, 
    71.2795, 71.27952, 71.27949, 71.27951, 71.27949, 71.27951, 71.27951, 
    71.27949, 71.27951, 71.27948, 71.27948, 71.2795, 71.27959, 71.27961, 
    71.27961, 71.27958, 71.2796, 71.27958, 71.27958, 71.2796, 71.2796, 
    71.27957, 71.27957, 71.27959, 71.27957, 71.27959, 71.27959, 71.27956, 
    71.27959, 71.27956, 71.27956, 71.27959, 71.27958, 71.27956, 71.27958, 
    71.27956, 71.27958, 71.27955, 71.27966, 71.27968, 71.27968, 71.27966, 
    71.27968, 71.27965, 71.27967, 71.27965, 71.27967, 71.27965, 71.27967, 
    71.27964, 71.27966, 71.27964, 71.27964, 71.27966, 71.27963, 71.27966, 
    71.27966, 71.27963, 71.27963, 71.27966, 71.27962, 71.27965, 71.27962, 
    71.27965, 71.27973, 71.27975, 71.27975, 71.27972, 71.27975, 71.27972, 
    71.27972, 71.27975, 71.27974, 71.27972, 71.27974, 71.27972, 71.27974, 
    71.27971, 71.27973, 71.27971, 71.27973, 71.27971, 71.27972, 71.2797, 
    71.2797, 71.27972, 71.27972, 71.27969, 71.27972, 71.27969, 71.27982, 
    71.2798, 71.2798, 71.27982, 71.27982, 71.27979, 71.27982, 71.27979, 
    71.27982, 71.27979, 71.27979, 71.27981, 71.27981, 71.27979, 71.27981, 
    71.27978, 71.2798, 71.27978, 71.27978, 71.2798, 71.27977, 71.27979, 
    71.27977, 71.27979, 71.27977, 71.27979, 71.2799, 71.27987, 71.27987, 
    71.27989, 71.27987, 71.27989, 71.27988, 71.27986, 71.27986, 71.27988, 
    71.27988, 71.27985, 71.27988, 71.27985, 71.27985, 71.27988, 71.27988, 
    71.27985, 71.27987, 71.27985, 71.27985, 71.27987, 71.27984, 71.27986, 
    71.27984, 71.27985 ;

 area = 9.902211e-05, 9.902174e-05, 9.902174e-05, 9.902209e-05, 9.902172e-05, 
    9.902208e-05, 9.902207e-05, 9.902169e-05, 9.902168e-05, 9.902204e-05, 
    9.902203e-05, 9.902166e-05, 9.902201e-05, 9.902164e-05, 9.902163e-05, 
    9.902199e-05, 9.902198e-05, 9.902161e-05, 9.902196e-05, 9.902159e-05, 
    9.902158e-05, 9.902194e-05, 9.902156e-05, 9.902192e-05, 9.902155e-05, 
    4.951087e-05, 9.902174e-05, 9.902138e-05, 9.902137e-05, 9.902173e-05, 
    9.902172e-05, 9.902135e-05, 9.90217e-05, 9.902133e-05, 9.902168e-05, 
    9.902132e-05, 9.90213e-05, 9.902166e-05, 9.902164e-05, 9.902128e-05, 
    9.902163e-05, 9.902126e-05, 9.902161e-05, 9.902124e-05, 9.902123e-05, 
    9.902159e-05, 9.902121e-05, 9.902157e-05, 9.902119e-05, 9.902156e-05, 
    9.902118e-05, 9.902155e-05, 9.902102e-05, 9.902138e-05, 9.902137e-05, 
    9.9021e-05, 9.902135e-05, 9.902099e-05, 9.902097e-05, 9.902133e-05, 
    9.902132e-05, 9.902095e-05, 9.90213e-05, 9.902093e-05, 9.902128e-05, 
    9.902092e-05, 9.902126e-05, 9.90209e-05, 9.902124e-05, 9.902088e-05, 
    9.902123e-05, 9.902086e-05, 9.902084e-05, 9.902121e-05, 9.902119e-05, 
    9.902083e-05, 9.902118e-05, 9.902081e-05, 9.902065e-05, 9.902102e-05, 
    9.9021e-05, 9.902064e-05, 9.902099e-05, 9.902062e-05, 9.902097e-05, 
    9.90206e-05, 9.902095e-05, 9.902059e-05, 9.902094e-05, 9.902057e-05, 
    9.902092e-05, 9.902055e-05, 9.902054e-05, 9.90209e-05, 9.902052e-05, 
    9.902088e-05, 9.902086e-05, 9.90205e-05, 9.902048e-05, 9.902084e-05, 
    9.902046e-05, 9.902083e-05, 9.902046e-05, 9.902081e-05, 9.902029e-05, 
    9.902065e-05, 9.902064e-05, 9.902028e-05, 9.902062e-05, 9.902026e-05, 
    9.902024e-05, 9.90206e-05, 9.902059e-05, 9.902022e-05, 9.90202e-05, 
    9.902057e-05, 9.902019e-05, 9.902055e-05, 9.902054e-05, 9.902017e-05, 
    9.902052e-05, 9.902015e-05, 9.902014e-05, 9.90205e-05, 9.902048e-05, 
    9.902012e-05, 9.902046e-05, 9.90201e-05, 9.902046e-05, 9.902009e-05, 
    9.901992e-05, 9.902028e-05, 9.901991e-05, 9.902028e-05, 9.902026e-05, 
    9.901989e-05, 9.901988e-05, 9.902024e-05, 9.902022e-05, 9.901986e-05, 
    9.90202e-05, 9.901984e-05, 9.901982e-05, 9.902019e-05, 9.90198e-05, 
    9.902017e-05, 9.901979e-05, 9.902015e-05, 9.901977e-05, 9.902013e-05, 
    9.902012e-05, 9.901975e-05, 9.90201e-05, 9.901973e-05, 9.901972e-05, 
    9.902009e-05, 9.901955e-05, 9.901992e-05, 9.901991e-05, 9.901955e-05, 
    9.90199e-05, 9.901953e-05, 9.901951e-05, 9.901988e-05, 9.901986e-05, 
    9.901949e-05, 9.901984e-05, 9.901947e-05, 9.901946e-05, 9.901982e-05, 
    9.901944e-05, 9.90198e-05, 9.901942e-05, 9.901979e-05, 9.90194e-05, 
    9.901977e-05, 9.901975e-05, 9.901939e-05, 9.901974e-05, 9.901937e-05, 
    9.901972e-05, 9.901936e-05, 9.901919e-05, 9.901955e-05, 9.901918e-05, 
    9.901955e-05, 9.901953e-05, 9.901916e-05, 9.901915e-05, 9.901951e-05, 
    9.90195e-05, 9.901913e-05, 9.901911e-05, 9.901947e-05, 9.90191e-05, 
    9.901946e-05, 9.901907e-05, 9.901944e-05, 9.901906e-05, 9.901942e-05, 
    9.901904e-05, 9.90194e-05, 9.901939e-05, 9.901902e-05, 9.901937e-05, 
    9.9019e-05, 9.901899e-05, 9.901936e-05, 9.901919e-05, 9.901883e-05, 
    9.901882e-05, 9.901918e-05, 9.90188e-05, 9.901916e-05, 9.901915e-05, 
    9.901878e-05, 9.901877e-05, 9.901913e-05, 9.901911e-05, 9.901875e-05, 
    9.901873e-05, 9.90191e-05, 9.901871e-05, 9.901907e-05, 9.90187e-05, 
    9.901906e-05, 9.901867e-05, 9.901904e-05, 9.901902e-05, 9.901866e-05, 
    9.901901e-05, 9.901864e-05, 9.901863e-05, 9.901899e-05, 9.901846e-05, 
    9.901883e-05, 9.901846e-05, 9.901882e-05, 9.90188e-05, 9.901843e-05, 
    9.901842e-05, 9.901878e-05, 9.90184e-05, 9.901876e-05, 9.901838e-05, 
    9.901875e-05, 9.901873e-05, 9.901836e-05, 9.901835e-05, 9.901871e-05, 
    9.90187e-05, 9.901833e-05, 9.901867e-05, 9.901831e-05, 9.901866e-05, 
    9.90183e-05, 9.901864e-05, 9.901827e-05, 9.901863e-05, 9.901827e-05, 
    9.90181e-05, 9.901846e-05, 9.901809e-05, 9.901846e-05, 9.901843e-05, 
    9.901807e-05, 9.901842e-05, 9.901806e-05, 9.901803e-05, 9.90184e-05, 
    9.901802e-05, 9.901838e-05, 9.901837e-05, 9.9018e-05, 9.901798e-05, 
    9.901835e-05, 9.901797e-05, 9.901833e-05, 9.901795e-05, 9.901831e-05, 
    9.901793e-05, 9.90183e-05, 9.901827e-05, 9.901791e-05, 9.901827e-05, 
    9.90179e-05, 9.90181e-05, 9.901774e-05, 9.901809e-05, 9.901772e-05, 
    9.901771e-05, 9.901807e-05, 9.901769e-05, 9.901806e-05, 9.901803e-05, 
    9.901767e-05, 9.901766e-05, 9.901802e-05, 9.9018e-05, 9.901763e-05, 
    9.901798e-05, 9.901762e-05, 9.90176e-05, 9.901796e-05, 9.901758e-05, 
    9.901795e-05, 9.901757e-05, 9.901793e-05, 9.901791e-05, 9.901755e-05, 
    9.90179e-05, 9.901754e-05, 9.901774e-05, 9.901737e-05, 9.901773e-05, 
    9.901736e-05, 9.901734e-05, 9.901771e-05, 9.901733e-05, 9.901768e-05, 
    9.901731e-05, 9.901767e-05, 9.901766e-05, 9.901728e-05, 9.901727e-05, 
    9.901763e-05, 9.901762e-05, 9.901726e-05, 9.901723e-05, 9.90176e-05, 
    9.901722e-05, 9.901758e-05, 9.901757e-05, 9.90172e-05, 9.901755e-05, 
    9.901718e-05, 9.901718e-05, 9.901754e-05 ;

 topo = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0 ;

 landfrac = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 landmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 pftmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 ACTUAL_IMMOB =
  5.20049e-14, 5.213718e-14, 5.211149e-14, 5.221808e-14, 5.215898e-14, 
    5.222874e-14, 5.203175e-14, 5.214241e-14, 5.207179e-14, 5.201684e-14, 
    5.242459e-14, 5.222284e-14, 5.263398e-14, 5.250555e-14, 5.282794e-14, 
    5.261398e-14, 5.287104e-14, 5.282182e-14, 5.297001e-14, 5.292758e-14, 
    5.311679e-14, 5.298958e-14, 5.321482e-14, 5.308646e-14, 5.310653e-14, 
    5.298538e-14, 5.226351e-14, 5.239947e-14, 5.225544e-14, 5.227484e-14, 
    5.226615e-14, 5.216018e-14, 5.210672e-14, 5.199481e-14, 5.201514e-14, 
    5.209735e-14, 5.228357e-14, 5.222042e-14, 5.237959e-14, 5.2376e-14, 
    5.255292e-14, 5.247318e-14, 5.277016e-14, 5.268585e-14, 5.292935e-14, 
    5.286815e-14, 5.292647e-14, 5.290879e-14, 5.29267e-14, 5.283694e-14, 
    5.28754e-14, 5.27964e-14, 5.248811e-14, 5.257879e-14, 5.23081e-14, 
    5.214496e-14, 5.203659e-14, 5.19596e-14, 5.197049e-14, 5.199123e-14, 
    5.209783e-14, 5.219801e-14, 5.227428e-14, 5.232526e-14, 5.237548e-14, 
    5.252724e-14, 5.260758e-14, 5.278718e-14, 5.275483e-14, 5.280965e-14, 
    5.286207e-14, 5.294995e-14, 5.29355e-14, 5.297419e-14, 5.280824e-14, 
    5.291854e-14, 5.273639e-14, 5.278623e-14, 5.238897e-14, 5.223747e-14, 
    5.217287e-14, 5.211642e-14, 5.197886e-14, 5.207386e-14, 5.203642e-14, 
    5.212552e-14, 5.218208e-14, 5.215412e-14, 5.232666e-14, 5.225961e-14, 
    5.261234e-14, 5.246054e-14, 5.285596e-14, 5.276147e-14, 5.28786e-14, 
    5.281885e-14, 5.292119e-14, 5.282909e-14, 5.29886e-14, 5.302328e-14, 
    5.299958e-14, 5.309065e-14, 5.282398e-14, 5.292645e-14, 5.215333e-14, 
    5.215789e-14, 5.217915e-14, 5.208566e-14, 5.207994e-14, 5.199425e-14, 
    5.207052e-14, 5.210297e-14, 5.218537e-14, 5.223406e-14, 5.228033e-14, 
    5.2382e-14, 5.249542e-14, 5.265388e-14, 5.27676e-14, 5.284375e-14, 
    5.279707e-14, 5.283828e-14, 5.279221e-14, 5.277061e-14, 5.301028e-14, 
    5.287575e-14, 5.307756e-14, 5.306641e-14, 5.29751e-14, 5.306766e-14, 
    5.216109e-14, 5.213484e-14, 5.204361e-14, 5.211501e-14, 5.198491e-14, 
    5.205773e-14, 5.209958e-14, 5.226097e-14, 5.229644e-14, 5.232927e-14, 
    5.239412e-14, 5.247727e-14, 5.262297e-14, 5.274961e-14, 5.286512e-14, 
    5.285667e-14, 5.285964e-14, 5.288541e-14, 5.282154e-14, 5.28959e-14, 
    5.290836e-14, 5.287575e-14, 5.306491e-14, 5.301091e-14, 5.306617e-14, 
    5.303102e-14, 5.214338e-14, 5.218755e-14, 5.216368e-14, 5.220855e-14, 
    5.217693e-14, 5.231742e-14, 5.235951e-14, 5.25563e-14, 5.247562e-14, 
    5.260404e-14, 5.248868e-14, 5.250912e-14, 5.260816e-14, 5.249493e-14, 
    5.27426e-14, 5.257469e-14, 5.288642e-14, 5.271889e-14, 5.28969e-14, 
    5.286462e-14, 5.291808e-14, 5.296591e-14, 5.302609e-14, 5.313698e-14, 
    5.311132e-14, 5.320402e-14, 5.225338e-14, 5.23106e-14, 5.230559e-14, 
    5.236546e-14, 5.240972e-14, 5.250561e-14, 5.26592e-14, 5.260147e-14, 
    5.270746e-14, 5.272871e-14, 5.256771e-14, 5.266656e-14, 5.23489e-14, 
    5.240025e-14, 5.23697e-14, 5.225788e-14, 5.261474e-14, 5.243172e-14, 
    5.276947e-14, 5.26705e-14, 5.295909e-14, 5.281563e-14, 5.309718e-14, 
    5.321724e-14, 5.333024e-14, 5.346198e-14, 5.234185e-14, 5.230298e-14, 
    5.237259e-14, 5.246877e-14, 5.255804e-14, 5.267654e-14, 5.268867e-14, 
    5.271085e-14, 5.27683e-14, 5.281657e-14, 5.271783e-14, 5.282868e-14, 
    5.241209e-14, 5.263062e-14, 5.228825e-14, 5.239142e-14, 5.246312e-14, 
    5.24317e-14, 5.259488e-14, 5.26333e-14, 5.278925e-14, 5.270868e-14, 
    5.318759e-14, 5.297597e-14, 5.356227e-14, 5.339874e-14, 5.228939e-14, 
    5.234173e-14, 5.252365e-14, 5.243713e-14, 5.268446e-14, 5.274524e-14, 
    5.279465e-14, 5.285774e-14, 5.286457e-14, 5.290192e-14, 5.284069e-14, 
    5.289952e-14, 5.267679e-14, 5.277638e-14, 5.250291e-14, 5.256951e-14, 
    5.253889e-14, 5.250527e-14, 5.260901e-14, 5.271937e-14, 5.272178e-14, 
    5.275714e-14, 5.285662e-14, 5.268546e-14, 5.321478e-14, 5.288811e-14, 
    5.239877e-14, 5.24994e-14, 5.251382e-14, 5.247485e-14, 5.273915e-14, 
    5.264345e-14, 5.290102e-14, 5.283148e-14, 5.294541e-14, 5.288881e-14, 
    5.288047e-14, 5.280774e-14, 5.276241e-14, 5.264783e-14, 5.255453e-14, 
    5.24805e-14, 5.249773e-14, 5.257902e-14, 5.272613e-14, 5.286516e-14, 
    5.283472e-14, 5.293676e-14, 5.266654e-14, 5.277991e-14, 5.273609e-14, 
    5.285031e-14, 5.259993e-14, 5.281303e-14, 5.254538e-14, 5.256888e-14, 
    5.264155e-14, 5.278756e-14, 5.281991e-14, 5.285435e-14, 5.283311e-14, 
    5.272988e-14, 5.271298e-14, 5.263979e-14, 5.261956e-14, 5.256377e-14, 
    5.251753e-14, 5.255976e-14, 5.260409e-14, 5.272994e-14, 5.284321e-14, 
    5.296658e-14, 5.299677e-14, 5.314058e-14, 5.302346e-14, 5.321659e-14, 
    5.305232e-14, 5.333657e-14, 5.282544e-14, 5.304758e-14, 5.264487e-14, 
    5.268834e-14, 5.276687e-14, 5.294686e-14, 5.284978e-14, 5.296333e-14, 
    5.271232e-14, 5.25818e-14, 5.254806e-14, 5.2485e-14, 5.254951e-14, 
    5.254426e-14, 5.260595e-14, 5.258614e-14, 5.273412e-14, 5.265465e-14, 
    5.288025e-14, 5.296245e-14, 5.319429e-14, 5.333613e-14, 5.34804e-14, 
    5.3544e-14, 5.356335e-14, 5.357144e-14 ;

 AGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX_LASTYEAR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 AR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_CROP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_PEATF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BCDEP =
  9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15 ;

 BGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BTRAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BUILDHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4PROD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_DIFF_SAT =
  -7.438852e-15, -7.432389e-15, -7.433646e-15, -7.428435e-15, -7.431327e-15, 
    -7.427914e-15, -7.437543e-15, -7.432131e-15, -7.435586e-15, 
    -7.438272e-15, -7.418334e-15, -7.428204e-15, -7.408229e-15, 
    -7.414502e-15, -7.398768e-15, -7.409201e-15, -7.396668e-15, 
    -7.399073e-15, -7.391849e-15, -7.393917e-15, -7.384681e-15, 
    -7.390894e-15, -7.379908e-15, -7.386166e-15, -7.385185e-15, 
    -7.391099e-15, -7.42622e-15, -7.419561e-15, -7.426614e-15, -7.425663e-15, 
    -7.426091e-15, -7.431265e-15, -7.433871e-15, -7.439349e-15, 
    -7.438355e-15, -7.434334e-15, -7.425237e-15, -7.428326e-15, 
    -7.420554e-15, -7.420729e-15, -7.412191e-15, -7.415983e-15, 
    -7.401592e-15, -7.405707e-15, -7.393831e-15, -7.396814e-15, 
    -7.393971e-15, -7.394833e-15, -7.393959e-15, -7.398335e-15, 
    -7.396459e-15, -7.400313e-15, -7.415253e-15, -7.410927e-15, -7.42404e-15, 
    -7.431999e-15, -7.437305e-15, -7.441069e-15, -7.440536e-15, 
    -7.439521e-15, -7.434311e-15, -7.429421e-15, -7.425696e-15, 
    -7.423206e-15, -7.420755e-15, -7.413431e-15, -7.409517e-15, 
    -7.400758e-15, -7.402342e-15, -7.399663e-15, -7.397112e-15, 
    -7.392825e-15, -7.39353e-15, -7.391642e-15, -7.399737e-15, -7.394354e-15, 
    -7.403243e-15, -7.40081e-15, -7.420071e-15, -7.427493e-15, -7.430637e-15, 
    -7.433404e-15, -7.440127e-15, -7.435482e-15, -7.437313e-15, 
    -7.432962e-15, -7.430198e-15, -7.431566e-15, -7.423138e-15, 
    -7.426412e-15, -7.409285e-15, -7.416596e-15, -7.397409e-15, 
    -7.402018e-15, -7.396305e-15, -7.39922e-15, -7.394226e-15, -7.39872e-15, 
    -7.390941e-15, -7.389247e-15, -7.390404e-15, -7.385966e-15, 
    -7.398969e-15, -7.393969e-15, -7.431604e-15, -7.43138e-15, -7.430342e-15, 
    -7.434905e-15, -7.435186e-15, -7.439376e-15, -7.435649e-15, 
    -7.434061e-15, -7.430039e-15, -7.427659e-15, -7.425399e-15, 
    -7.420434e-15, -7.414893e-15, -7.407262e-15, -7.401719e-15, 
    -7.398005e-15, -7.400283e-15, -7.398272e-15, -7.400519e-15, 
    -7.401574e-15, -7.389881e-15, -7.396441e-15, -7.386604e-15, 
    -7.387149e-15, -7.391597e-15, -7.387088e-15, -7.431224e-15, 
    -7.432507e-15, -7.436963e-15, -7.433476e-15, -7.439833e-15, 
    -7.436272e-15, -7.434224e-15, -7.42634e-15, -7.424614e-15, -7.423009e-15, 
    -7.419843e-15, -7.415784e-15, -7.408771e-15, -7.402593e-15, 
    -7.396963e-15, -7.397376e-15, -7.397231e-15, -7.395972e-15, 
    -7.399088e-15, -7.395462e-15, -7.394852e-15, -7.396444e-15, 
    -7.387222e-15, -7.389854e-15, -7.387161e-15, -7.388875e-15, 
    -7.432091e-15, -7.429932e-15, -7.431098e-15, -7.428904e-15, 
    -7.430448e-15, -7.423581e-15, -7.421525e-15, -7.41202e-15, -7.415862e-15, 
    -7.409693e-15, -7.415226e-15, -7.414328e-15, -7.409482e-15, 
    -7.415024e-15, -7.40293e-15, -7.41112e-15, -7.395923e-15, -7.404081e-15, 
    -7.395412e-15, -7.396988e-15, -7.394382e-15, -7.392046e-15, 
    -7.389114e-15, -7.383704e-15, -7.384957e-15, -7.380439e-15, 
    -7.426716e-15, -7.423918e-15, -7.424168e-15, -7.421243e-15, -7.41908e-15, 
    -7.414503e-15, -7.407005e-15, -7.409824e-15, -7.404654e-15, 
    -7.403616e-15, -7.411473e-15, -7.406644e-15, -7.422048e-15, 
    -7.419536e-15, -7.421034e-15, -7.426494e-15, -7.40917e-15, -7.418e-15, 
    -7.401626e-15, -7.406454e-15, -7.392379e-15, -7.39937e-15, -7.385646e-15, 
    -7.379784e-15, -7.37429e-15, -7.367862e-15, -7.422395e-15, -7.424295e-15, 
    -7.420896e-15, -7.416192e-15, -7.411942e-15, -7.40616e-15, -7.40557e-15, 
    -7.404487e-15, -7.401686e-15, -7.399331e-15, -7.404141e-15, 
    -7.398741e-15, -7.418947e-15, -7.408397e-15, -7.425011e-15, 
    -7.419966e-15, -7.416471e-15, -7.418007e-15, -7.410147e-15, 
    -7.408272e-15, -7.400659e-15, -7.404594e-15, -7.381227e-15, 
    -7.391549e-15, -7.362985e-15, -7.370945e-15, -7.424959e-15, 
    -7.422403e-15, -7.413617e-15, -7.417742e-15, -7.405775e-15, 
    -7.402809e-15, -7.400401e-15, -7.39732e-15, -7.39699e-15, -7.395166e-15, 
    -7.398155e-15, -7.395285e-15, -7.406147e-15, -7.40129e-15, -7.414636e-15, 
    -7.411382e-15, -7.412879e-15, -7.414521e-15, -7.409457e-15, 
    -7.404064e-15, -7.403955e-15, -7.402226e-15, -7.397349e-15, 
    -7.405727e-15, -7.379887e-15, -7.395817e-15, -7.419617e-15, 
    -7.414797e-15, -7.414101e-15, -7.415904e-15, -7.403105e-15, 
    -7.407774e-15, -7.395212e-15, -7.398604e-15, -7.393048e-15, 
    -7.395807e-15, -7.396214e-15, -7.399762e-15, -7.401971e-15, 
    -7.407559e-15, -7.412113e-15, -7.415628e-15, -7.414888e-15, 
    -7.410917e-15, -7.403736e-15, -7.396957e-15, -7.398441e-15, -7.39347e-15, 
    -7.406649e-15, -7.401115e-15, -7.403252e-15, -7.397684e-15, 
    -7.409898e-15, -7.39948e-15, -7.412563e-15, -7.411415e-15, -7.407867e-15, 
    -7.400737e-15, -7.399168e-15, -7.397485e-15, -7.398524e-15, 
    -7.403555e-15, -7.404382e-15, -7.407954e-15, -7.408939e-15, 
    -7.411665e-15, -7.413922e-15, -7.411859e-15, -7.409693e-15, 
    -7.403555e-15, -7.398028e-15, -7.392012e-15, -7.390544e-15, 
    -7.383516e-15, -7.389229e-15, -7.379797e-15, -7.387804e-15, 
    -7.373961e-15, -7.398884e-15, -7.38805e-15, -7.407707e-15, -7.405587e-15, 
    -7.401747e-15, -7.392967e-15, -7.39771e-15, -7.392166e-15, -7.404415e-15, 
    -7.410777e-15, -7.412431e-15, -7.415407e-15, -7.412361e-15, 
    -7.412617e-15, -7.409607e-15, -7.410574e-15, -7.403351e-15, 
    -7.407229e-15, -7.396222e-15, -7.392211e-15, -7.38091e-15, -7.373994e-15, 
    -7.366975e-15, -7.363877e-15, -7.362936e-15, -7.362542e-15 ;

 CH4_SURF_DIFF_UNSAT =
  4.975673e-14, 4.923995e-14, 4.934057e-14, 4.892274e-14, 4.915469e-14, 
    4.888088e-14, 4.965213e-14, 4.921937e-14, 4.949579e-14, 4.971033e-14, 
    4.810867e-14, 4.890409e-14, 4.727853e-14, 4.778878e-14, 4.650419e-14, 
    4.735798e-14, 4.633153e-14, 4.652897e-14, 4.593426e-14, 4.610485e-14, 
    4.534177e-14, 4.585547e-14, 4.494506e-14, 4.546463e-14, 4.538342e-14, 
    4.587238e-14, 4.874442e-14, 4.820788e-14, 4.877613e-14, 4.869975e-14, 
    4.873405e-14, 4.914987e-14, 4.935895e-14, 4.979622e-14, 4.971694e-14, 
    4.939577e-14, 4.866539e-14, 4.891376e-14, 4.828726e-14, 4.830144e-14, 
    4.760096e-14, 4.791725e-14, 4.673565e-14, 4.70723e-14, 4.609774e-14, 
    4.634333e-14, 4.610926e-14, 4.618028e-14, 4.610834e-14, 4.64684e-14, 
    4.631422e-14, 4.663074e-14, 4.785807e-14, 4.749815e-14, 4.85689e-14, 
    4.920911e-14, 4.963316e-14, 4.993331e-14, 4.989091e-14, 4.981004e-14, 
    4.939389e-14, 4.900171e-14, 4.870216e-14, 4.850146e-14, 4.830348e-14, 
    4.770232e-14, 4.738356e-14, 4.666744e-14, 4.679698e-14, 4.657754e-14, 
    4.636775e-14, 4.601485e-14, 4.6073e-14, 4.591732e-14, 4.658339e-14, 
    4.614098e-14, 4.687071e-14, 4.667142e-14, 4.824929e-14, 4.884681e-14, 
    4.909983e-14, 4.932122e-14, 4.98583e-14, 4.948758e-14, 4.963382e-14, 
    4.928576e-14, 4.906415e-14, 4.917381e-14, 4.849597e-14, 4.875982e-14, 
    4.736464e-14, 4.796715e-14, 4.639223e-14, 4.677041e-14, 4.630148e-14, 
    4.654094e-14, 4.613041e-14, 4.649993e-14, 4.585938e-14, 4.571955e-14, 
    4.581511e-14, 4.544786e-14, 4.652038e-14, 4.610923e-14, 4.917686e-14, 
    4.915898e-14, 4.907569e-14, 4.944149e-14, 4.946385e-14, 4.979838e-14, 
    4.950078e-14, 4.937386e-14, 4.905132e-14, 4.886018e-14, 4.867829e-14, 
    4.827764e-14, 4.782898e-14, 4.719946e-14, 4.674592e-14, 4.64412e-14, 
    4.662814e-14, 4.646311e-14, 4.664756e-14, 4.673397e-14, 4.577193e-14, 
    4.631276e-14, 4.550073e-14, 4.554577e-14, 4.591361e-14, 4.554069e-14, 
    4.914643e-14, 4.92493e-14, 4.960581e-14, 4.932688e-14, 4.983477e-14, 
    4.955063e-14, 4.9387e-14, 4.875424e-14, 4.861496e-14, 4.84856e-14, 
    4.822989e-14, 4.790108e-14, 4.732251e-14, 4.681767e-14, 4.635555e-14, 
    4.638946e-14, 4.637752e-14, 4.627409e-14, 4.653013e-14, 4.623203e-14, 
    4.618192e-14, 4.631286e-14, 4.55518e-14, 4.576957e-14, 4.554672e-14, 
    4.568856e-14, 4.921587e-14, 4.904273e-14, 4.913631e-14, 4.896028e-14, 
    4.908429e-14, 4.853204e-14, 4.83661e-14, 4.758729e-14, 4.790754e-14, 
    4.739776e-14, 4.785587e-14, 4.777463e-14, 4.738097e-14, 4.783101e-14, 
    4.684549e-14, 4.751415e-14, 4.627007e-14, 4.693994e-14, 4.6228e-14, 
    4.635755e-14, 4.614304e-14, 4.595066e-14, 4.570839e-14, 4.52604e-14, 
    4.536426e-14, 4.498901e-14, 4.87843e-14, 4.855905e-14, 4.857895e-14, 
    4.834297e-14, 4.816821e-14, 4.77887e-14, 4.717838e-14, 4.740817e-14, 
    4.698615e-14, 4.690128e-14, 4.754237e-14, 4.714898e-14, 4.840817e-14, 
    4.820535e-14, 4.832618e-14, 4.87665e-14, 4.735516e-14, 4.808103e-14, 
    4.67384e-14, 4.713339e-14, 4.597809e-14, 4.655355e-14, 4.542138e-14, 
    4.493501e-14, 4.447634e-14, 4.393854e-14, 4.843605e-14, 4.858925e-14, 
    4.83149e-14, 4.793446e-14, 4.758068e-14, 4.710931e-14, 4.706104e-14, 
    4.697254e-14, 4.674317e-14, 4.655005e-14, 4.694449e-14, 4.650161e-14, 
    4.815815e-14, 4.729205e-14, 4.864707e-14, 4.824019e-14, 4.795693e-14, 
    4.808131e-14, 4.743443e-14, 4.728162e-14, 4.66592e-14, 4.698127e-14, 
    4.505512e-14, 4.590991e-14, 4.352822e-14, 4.419688e-14, 4.864272e-14, 
    4.843661e-14, 4.771697e-14, 4.805987e-14, 4.707783e-14, 4.683523e-14, 
    4.663781e-14, 4.638502e-14, 4.635775e-14, 4.620779e-14, 4.645346e-14, 
    4.621752e-14, 4.71083e-14, 4.671081e-14, 4.779944e-14, 4.753509e-14, 
    4.765677e-14, 4.77901e-14, 4.737826e-14, 4.693827e-14, 4.692896e-14, 
    4.678761e-14, 4.638849e-14, 4.707384e-14, 4.494431e-14, 4.626235e-14, 
    4.821155e-14, 4.781295e-14, 4.775609e-14, 4.791074e-14, 4.685956e-14, 
    4.724113e-14, 4.621146e-14, 4.649037e-14, 4.603316e-14, 4.62605e-14, 
    4.629392e-14, 4.658543e-14, 4.676664e-14, 4.722364e-14, 4.759458e-14, 
    4.788836e-14, 4.781997e-14, 4.749728e-14, 4.691134e-14, 4.635524e-14, 
    4.64772e-14, 4.606796e-14, 4.714921e-14, 4.66966e-14, 4.687165e-14, 
    4.641486e-14, 4.741425e-14, 4.656329e-14, 4.763104e-14, 4.753771e-14, 
    4.72487e-14, 4.666579e-14, 4.653671e-14, 4.639859e-14, 4.648385e-14, 
    4.689646e-14, 4.696401e-14, 4.725575e-14, 4.733616e-14, 4.755804e-14, 
    4.774147e-14, 4.757386e-14, 4.739765e-14, 4.689633e-14, 4.644323e-14, 
    4.59479e-14, 4.582651e-14, 4.524534e-14, 4.571845e-14, 4.493692e-14, 
    4.560138e-14, 4.444972e-14, 4.651399e-14, 4.562108e-14, 4.723556e-14, 
    4.706239e-14, 4.67486e-14, 4.602694e-14, 4.641702e-14, 4.596078e-14, 
    4.696667e-14, 4.748609e-14, 4.762034e-14, 4.78705e-14, 4.761463e-14, 
    4.763544e-14, 4.739041e-14, 4.74692e-14, 4.687966e-14, 4.719659e-14, 
    4.629473e-14, 4.596442e-14, 4.502834e-14, 4.445201e-14, 4.386365e-14, 
    4.360325e-14, 4.352393e-14, 4.349075e-14 ;

 CH4_SURF_EBUL_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_EBUL_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_CTRUNC =
  1.931904e-23, 1.931903e-23, 1.931903e-23, 1.931903e-23, 1.931903e-23, 
    1.931903e-23, 1.931904e-23, 1.931903e-23, 1.931903e-23, 1.931904e-23, 
    1.931902e-23, 1.931903e-23, 1.9319e-23, 1.931901e-23, 1.931899e-23, 
    1.9319e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 
    1.931898e-23, 1.931898e-23, 1.931897e-23, 1.931898e-23, 1.931898e-23, 
    1.931898e-23, 1.931902e-23, 1.931902e-23, 1.931903e-23, 1.931902e-23, 
    1.931902e-23, 1.931903e-23, 1.931903e-23, 1.931904e-23, 1.931904e-23, 
    1.931903e-23, 1.931902e-23, 1.931903e-23, 1.931902e-23, 1.931902e-23, 
    1.931901e-23, 1.931901e-23, 1.9319e-23, 1.9319e-23, 1.931899e-23, 
    1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 
    1.931899e-23, 1.9319e-23, 1.931901e-23, 1.931901e-23, 1.931902e-23, 
    1.931903e-23, 1.931904e-23, 1.931904e-23, 1.931904e-23, 1.931904e-23, 
    1.931903e-23, 1.931903e-23, 1.931902e-23, 1.931902e-23, 1.931902e-23, 
    1.931901e-23, 1.9319e-23, 1.9319e-23, 1.9319e-23, 1.931899e-23, 
    1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931898e-23, 1.931899e-23, 
    1.931899e-23, 1.9319e-23, 1.9319e-23, 1.931902e-23, 1.931903e-23, 
    1.931903e-23, 1.931903e-23, 1.931904e-23, 1.931903e-23, 1.931904e-23, 
    1.931903e-23, 1.931903e-23, 1.931903e-23, 1.931902e-23, 1.931902e-23, 
    1.9319e-23, 1.931901e-23, 1.931899e-23, 1.9319e-23, 1.931899e-23, 
    1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931898e-23, 1.931898e-23, 
    1.931898e-23, 1.931898e-23, 1.931899e-23, 1.931899e-23, 1.931903e-23, 
    1.931903e-23, 1.931903e-23, 1.931903e-23, 1.931903e-23, 1.931904e-23, 
    1.931903e-23, 1.931903e-23, 1.931903e-23, 1.931903e-23, 1.931902e-23, 
    1.931902e-23, 1.931901e-23, 1.9319e-23, 1.9319e-23, 1.931899e-23, 
    1.9319e-23, 1.931899e-23, 1.9319e-23, 1.9319e-23, 1.931898e-23, 
    1.931899e-23, 1.931898e-23, 1.931898e-23, 1.931898e-23, 1.931898e-23, 
    1.931903e-23, 1.931903e-23, 1.931904e-23, 1.931903e-23, 1.931904e-23, 
    1.931903e-23, 1.931903e-23, 1.931902e-23, 1.931902e-23, 1.931902e-23, 
    1.931902e-23, 1.931901e-23, 1.9319e-23, 1.9319e-23, 1.931899e-23, 
    1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 
    1.931899e-23, 1.931899e-23, 1.931898e-23, 1.931898e-23, 1.931898e-23, 
    1.931898e-23, 1.931903e-23, 1.931903e-23, 1.931903e-23, 1.931903e-23, 
    1.931903e-23, 1.931902e-23, 1.931902e-23, 1.931901e-23, 1.931901e-23, 
    1.9319e-23, 1.931901e-23, 1.931901e-23, 1.9319e-23, 1.931901e-23, 
    1.9319e-23, 1.931901e-23, 1.931899e-23, 1.9319e-23, 1.931899e-23, 
    1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931898e-23, 1.931898e-23, 
    1.931898e-23, 1.931897e-23, 1.931903e-23, 1.931902e-23, 1.931902e-23, 
    1.931902e-23, 1.931902e-23, 1.931901e-23, 1.9319e-23, 1.931901e-23, 
    1.9319e-23, 1.9319e-23, 1.931901e-23, 1.9319e-23, 1.931902e-23, 
    1.931902e-23, 1.931902e-23, 1.931903e-23, 1.9319e-23, 1.931901e-23, 
    1.9319e-23, 1.9319e-23, 1.931899e-23, 1.931899e-23, 1.931898e-23, 
    1.931897e-23, 1.931897e-23, 1.931896e-23, 1.931902e-23, 1.931902e-23, 
    1.931902e-23, 1.931901e-23, 1.931901e-23, 1.9319e-23, 1.9319e-23, 
    1.9319e-23, 1.9319e-23, 1.931899e-23, 1.9319e-23, 1.931899e-23, 
    1.931902e-23, 1.9319e-23, 1.931902e-23, 1.931902e-23, 1.931901e-23, 
    1.931901e-23, 1.931901e-23, 1.9319e-23, 1.9319e-23, 1.9319e-23, 
    1.931897e-23, 1.931898e-23, 1.931895e-23, 1.931896e-23, 1.931902e-23, 
    1.931902e-23, 1.931901e-23, 1.931901e-23, 1.9319e-23, 1.9319e-23, 
    1.9319e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 
    1.931899e-23, 1.9319e-23, 1.9319e-23, 1.931901e-23, 1.931901e-23, 
    1.931901e-23, 1.931901e-23, 1.9319e-23, 1.9319e-23, 1.9319e-23, 
    1.9319e-23, 1.931899e-23, 1.9319e-23, 1.931897e-23, 1.931899e-23, 
    1.931902e-23, 1.931901e-23, 1.931901e-23, 1.931901e-23, 1.9319e-23, 
    1.9319e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 
    1.931899e-23, 1.931899e-23, 1.9319e-23, 1.9319e-23, 1.931901e-23, 
    1.931901e-23, 1.931901e-23, 1.931901e-23, 1.9319e-23, 1.931899e-23, 
    1.931899e-23, 1.931899e-23, 1.9319e-23, 1.9319e-23, 1.9319e-23, 
    1.931899e-23, 1.931901e-23, 1.931899e-23, 1.931901e-23, 1.931901e-23, 
    1.9319e-23, 1.9319e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 
    1.9319e-23, 1.9319e-23, 1.9319e-23, 1.9319e-23, 1.931901e-23, 
    1.931901e-23, 1.931901e-23, 1.9319e-23, 1.9319e-23, 1.931899e-23, 
    1.931899e-23, 1.931898e-23, 1.931898e-23, 1.931898e-23, 1.931897e-23, 
    1.931898e-23, 1.931897e-23, 1.931899e-23, 1.931898e-23, 1.9319e-23, 
    1.9319e-23, 1.9319e-23, 1.931899e-23, 1.931899e-23, 1.931899e-23, 
    1.9319e-23, 1.931901e-23, 1.931901e-23, 1.931901e-23, 1.931901e-23, 
    1.931901e-23, 1.9319e-23, 1.931901e-23, 1.9319e-23, 1.9319e-23, 
    1.931899e-23, 1.931899e-23, 1.931897e-23, 1.931897e-23, 1.931896e-23, 
    1.931895e-23, 1.931895e-23, 1.931895e-23 ;

 COL_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_NTRUNC =
  1.975319e-24, 1.975318e-24, 1.975318e-24, 1.975317e-24, 1.975317e-24, 
    1.975317e-24, 1.975318e-24, 1.975318e-24, 1.975318e-24, 1.975319e-24, 
    1.975315e-24, 1.975317e-24, 1.975314e-24, 1.975315e-24, 1.975312e-24, 
    1.975314e-24, 1.975312e-24, 1.975312e-24, 1.975311e-24, 1.975311e-24, 
    1.97531e-24, 1.975311e-24, 1.975309e-24, 1.97531e-24, 1.97531e-24, 
    1.975311e-24, 1.975317e-24, 1.975316e-24, 1.975317e-24, 1.975317e-24, 
    1.975317e-24, 1.975317e-24, 1.975318e-24, 1.975319e-24, 1.975319e-24, 
    1.975318e-24, 1.975317e-24, 1.975317e-24, 1.975316e-24, 1.975316e-24, 
    1.975314e-24, 1.975315e-24, 1.975313e-24, 1.975313e-24, 1.975311e-24, 
    1.975312e-24, 1.975311e-24, 1.975312e-24, 1.975311e-24, 1.975312e-24, 
    1.975312e-24, 1.975312e-24, 1.975315e-24, 1.975314e-24, 1.975316e-24, 
    1.975318e-24, 1.975318e-24, 1.975319e-24, 1.975319e-24, 1.975319e-24, 
    1.975318e-24, 1.975317e-24, 1.975317e-24, 1.975316e-24, 1.975316e-24, 
    1.975315e-24, 1.975314e-24, 1.975313e-24, 1.975313e-24, 1.975312e-24, 
    1.975312e-24, 1.975311e-24, 1.975311e-24, 1.975311e-24, 1.975312e-24, 
    1.975312e-24, 1.975313e-24, 1.975313e-24, 1.975316e-24, 1.975317e-24, 
    1.975317e-24, 1.975318e-24, 1.975319e-24, 1.975318e-24, 1.975318e-24, 
    1.975318e-24, 1.975317e-24, 1.975318e-24, 1.975316e-24, 1.975317e-24, 
    1.975314e-24, 1.975315e-24, 1.975312e-24, 1.975313e-24, 1.975312e-24, 
    1.975312e-24, 1.975312e-24, 1.975312e-24, 1.975311e-24, 1.975311e-24, 
    1.975311e-24, 1.97531e-24, 1.975312e-24, 1.975311e-24, 1.975318e-24, 
    1.975317e-24, 1.975317e-24, 1.975318e-24, 1.975318e-24, 1.975319e-24, 
    1.975318e-24, 1.975318e-24, 1.975317e-24, 1.975317e-24, 1.975317e-24, 
    1.975316e-24, 1.975315e-24, 1.975314e-24, 1.975313e-24, 1.975312e-24, 
    1.975312e-24, 1.975312e-24, 1.975313e-24, 1.975313e-24, 1.975311e-24, 
    1.975312e-24, 1.97531e-24, 1.97531e-24, 1.975311e-24, 1.97531e-24, 
    1.975317e-24, 1.975318e-24, 1.975318e-24, 1.975318e-24, 1.975319e-24, 
    1.975318e-24, 1.975318e-24, 1.975317e-24, 1.975316e-24, 1.975316e-24, 
    1.975316e-24, 1.975315e-24, 1.975314e-24, 1.975313e-24, 1.975312e-24, 
    1.975312e-24, 1.975312e-24, 1.975312e-24, 1.975312e-24, 1.975312e-24, 
    1.975312e-24, 1.975312e-24, 1.97531e-24, 1.975311e-24, 1.97531e-24, 
    1.975311e-24, 1.975318e-24, 1.975317e-24, 1.975317e-24, 1.975317e-24, 
    1.975317e-24, 1.975316e-24, 1.975316e-24, 1.975314e-24, 1.975315e-24, 
    1.975314e-24, 1.975315e-24, 1.975315e-24, 1.975314e-24, 1.975315e-24, 
    1.975313e-24, 1.975314e-24, 1.975312e-24, 1.975313e-24, 1.975312e-24, 
    1.975312e-24, 1.975312e-24, 1.975311e-24, 1.975311e-24, 1.97531e-24, 
    1.97531e-24, 1.975309e-24, 1.975317e-24, 1.975316e-24, 1.975316e-24, 
    1.975316e-24, 1.975316e-24, 1.975315e-24, 1.975314e-24, 1.975314e-24, 
    1.975313e-24, 1.975313e-24, 1.975314e-24, 1.975314e-24, 1.975316e-24, 
    1.975316e-24, 1.975316e-24, 1.975317e-24, 1.975314e-24, 1.975315e-24, 
    1.975313e-24, 1.975313e-24, 1.975311e-24, 1.975312e-24, 1.97531e-24, 
    1.975309e-24, 1.975308e-24, 1.975307e-24, 1.975316e-24, 1.975316e-24, 
    1.975316e-24, 1.975315e-24, 1.975314e-24, 1.975313e-24, 1.975313e-24, 
    1.975313e-24, 1.975313e-24, 1.975312e-24, 1.975313e-24, 1.975312e-24, 
    1.975315e-24, 1.975314e-24, 1.975316e-24, 1.975316e-24, 1.975315e-24, 
    1.975315e-24, 1.975314e-24, 1.975314e-24, 1.975313e-24, 1.975313e-24, 
    1.975309e-24, 1.975311e-24, 1.975307e-24, 1.975308e-24, 1.975316e-24, 
    1.975316e-24, 1.975315e-24, 1.975315e-24, 1.975313e-24, 1.975313e-24, 
    1.975312e-24, 1.975312e-24, 1.975312e-24, 1.975312e-24, 1.975312e-24, 
    1.975312e-24, 1.975313e-24, 1.975313e-24, 1.975315e-24, 1.975314e-24, 
    1.975315e-24, 1.975315e-24, 1.975314e-24, 1.975313e-24, 1.975313e-24, 
    1.975313e-24, 1.975312e-24, 1.975313e-24, 1.975309e-24, 1.975312e-24, 
    1.975316e-24, 1.975315e-24, 1.975315e-24, 1.975315e-24, 1.975313e-24, 
    1.975314e-24, 1.975312e-24, 1.975312e-24, 1.975311e-24, 1.975312e-24, 
    1.975312e-24, 1.975312e-24, 1.975313e-24, 1.975314e-24, 1.975314e-24, 
    1.975315e-24, 1.975315e-24, 1.975314e-24, 1.975313e-24, 1.975312e-24, 
    1.975312e-24, 1.975311e-24, 1.975314e-24, 1.975313e-24, 1.975313e-24, 
    1.975312e-24, 1.975314e-24, 1.975312e-24, 1.975314e-24, 1.975314e-24, 
    1.975314e-24, 1.975313e-24, 1.975312e-24, 1.975312e-24, 1.975312e-24, 
    1.975313e-24, 1.975313e-24, 1.975314e-24, 1.975314e-24, 1.975314e-24, 
    1.975315e-24, 1.975314e-24, 1.975314e-24, 1.975313e-24, 1.975312e-24, 
    1.975311e-24, 1.975311e-24, 1.97531e-24, 1.975311e-24, 1.975309e-24, 
    1.97531e-24, 1.975308e-24, 1.975312e-24, 1.975311e-24, 1.975314e-24, 
    1.975313e-24, 1.975313e-24, 1.975311e-24, 1.975312e-24, 1.975311e-24, 
    1.975313e-24, 1.975314e-24, 1.975314e-24, 1.975315e-24, 1.975314e-24, 
    1.975314e-24, 1.975314e-24, 1.975314e-24, 1.975313e-24, 1.975314e-24, 
    1.975312e-24, 1.975311e-24, 1.975309e-24, 1.975308e-24, 1.975307e-24, 
    1.975307e-24, 1.975307e-24, 1.975307e-24 ;

 CONC_CH4_SAT =
  3.550062e-08, 3.549992e-08, 3.550007e-08, 3.549946e-08, 3.549982e-08, 
    3.54994e-08, 3.55005e-08, 3.549988e-08, 3.550029e-08, 3.550059e-08, 
    3.549816e-08, 3.549944e-08, 3.549736e-08, 3.549821e-08, 3.549607e-08, 
    3.549747e-08, 3.549578e-08, 3.549615e-08, 3.549513e-08, 3.549543e-08, 
    3.549399e-08, 3.549499e-08, 3.549328e-08, 3.549425e-08, 3.549409e-08, 
    3.549502e-08, 3.549923e-08, 3.549831e-08, 3.549927e-08, 3.549914e-08, 
    3.549921e-08, 3.54998e-08, 3.550005e-08, 3.55007e-08, 3.550059e-08, 
    3.550013e-08, 3.549909e-08, 3.549948e-08, 3.549856e-08, 3.549858e-08, 
    3.549792e-08, 3.549798e-08, 3.54965e-08, 3.549707e-08, 3.549542e-08, 
    3.549584e-08, 3.549543e-08, 3.549556e-08, 3.549543e-08, 3.549605e-08, 
    3.549578e-08, 3.549633e-08, 3.549788e-08, 3.549774e-08, 3.549896e-08, 
    3.549982e-08, 3.550047e-08, 3.550088e-08, 3.550083e-08, 3.55007e-08, 
    3.550013e-08, 3.54996e-08, 3.549918e-08, 3.549888e-08, 3.549858e-08, 
    3.5498e-08, 3.549753e-08, 3.549637e-08, 3.549662e-08, 3.549622e-08, 
    3.549588e-08, 3.549526e-08, 3.549537e-08, 3.549508e-08, 3.549625e-08, 
    3.549547e-08, 3.549675e-08, 3.54964e-08, 3.549837e-08, 3.549938e-08, 
    3.549968e-08, 3.550004e-08, 3.550078e-08, 3.550026e-08, 3.550046e-08, 
    3.550001e-08, 3.549969e-08, 3.549985e-08, 3.549887e-08, 3.549926e-08, 
    3.54975e-08, 3.549804e-08, 3.549592e-08, 3.549657e-08, 3.549577e-08, 
    3.549619e-08, 3.549546e-08, 3.549611e-08, 3.549499e-08, 3.549472e-08, 
    3.54949e-08, 3.549425e-08, 3.549615e-08, 3.549542e-08, 3.549985e-08, 
    3.549982e-08, 3.549971e-08, 3.55002e-08, 3.550023e-08, 3.55007e-08, 
    3.55003e-08, 3.550011e-08, 3.549968e-08, 3.54994e-08, 3.549913e-08, 
    3.549853e-08, 3.549782e-08, 3.549725e-08, 3.549652e-08, 3.549602e-08, 
    3.549634e-08, 3.549605e-08, 3.549637e-08, 3.549652e-08, 3.549481e-08, 
    3.549577e-08, 3.549434e-08, 3.549443e-08, 3.549507e-08, 3.549442e-08, 
    3.549981e-08, 3.549996e-08, 3.550043e-08, 3.550007e-08, 3.550075e-08, 
    3.550036e-08, 3.550011e-08, 3.549922e-08, 3.549905e-08, 3.549884e-08, 
    3.549847e-08, 3.549795e-08, 3.549746e-08, 3.549663e-08, 3.549587e-08, 
    3.549593e-08, 3.54959e-08, 3.549572e-08, 3.549616e-08, 3.549565e-08, 
    3.549555e-08, 3.549579e-08, 3.549444e-08, 3.549483e-08, 3.549443e-08, 
    3.549469e-08, 3.549991e-08, 3.549966e-08, 3.54998e-08, 3.549954e-08, 
    3.549971e-08, 3.549888e-08, 3.549863e-08, 3.549786e-08, 3.549796e-08, 
    3.549757e-08, 3.549789e-08, 3.549819e-08, 3.549749e-08, 3.549829e-08, 
    3.549665e-08, 3.549773e-08, 3.549571e-08, 3.549678e-08, 3.549564e-08, 
    3.549587e-08, 3.54955e-08, 3.549514e-08, 3.549472e-08, 3.549388e-08, 
    3.549408e-08, 3.549338e-08, 3.549929e-08, 3.549894e-08, 3.5499e-08, 
    3.549864e-08, 3.549836e-08, 3.549822e-08, 3.549723e-08, 3.549762e-08, 
    3.549694e-08, 3.549679e-08, 3.549784e-08, 3.549717e-08, 3.549872e-08, 
    3.549838e-08, 3.54986e-08, 3.549925e-08, 3.54975e-08, 3.54982e-08, 
    3.549651e-08, 3.549717e-08, 3.549519e-08, 3.549617e-08, 3.549419e-08, 
    3.549322e-08, 3.549241e-08, 3.549129e-08, 3.549877e-08, 3.549901e-08, 
    3.54986e-08, 3.549797e-08, 3.549789e-08, 3.549712e-08, 3.549706e-08, 
    3.54969e-08, 3.549653e-08, 3.54962e-08, 3.549683e-08, 3.549612e-08, 
    3.549825e-08, 3.549741e-08, 3.549908e-08, 3.549843e-08, 3.549802e-08, 
    3.549823e-08, 3.549767e-08, 3.549742e-08, 3.549636e-08, 3.549693e-08, 
    3.549344e-08, 3.549503e-08, 3.54905e-08, 3.549182e-08, 3.549909e-08, 
    3.549878e-08, 3.549809e-08, 3.54982e-08, 3.549708e-08, 3.549667e-08, 
    3.549636e-08, 3.54959e-08, 3.549587e-08, 3.54956e-08, 3.549604e-08, 
    3.549562e-08, 3.549712e-08, 3.549647e-08, 3.549825e-08, 3.549781e-08, 
    3.549802e-08, 3.549823e-08, 3.549758e-08, 3.549681e-08, 3.549684e-08, 
    3.549658e-08, 3.549577e-08, 3.549708e-08, 3.549315e-08, 3.549557e-08, 
    3.549845e-08, 3.549821e-08, 3.549817e-08, 3.549798e-08, 3.549671e-08, 
    3.549734e-08, 3.549561e-08, 3.54961e-08, 3.54953e-08, 3.54957e-08, 
    3.549576e-08, 3.549626e-08, 3.549656e-08, 3.54973e-08, 3.549791e-08, 
    3.549795e-08, 3.549828e-08, 3.549775e-08, 3.549678e-08, 3.549585e-08, 
    3.549605e-08, 3.549536e-08, 3.54972e-08, 3.549643e-08, 3.549671e-08, 
    3.549596e-08, 3.549762e-08, 3.549609e-08, 3.549798e-08, 3.549783e-08, 
    3.549735e-08, 3.549635e-08, 3.549618e-08, 3.549592e-08, 3.549609e-08, 
    3.549676e-08, 3.549688e-08, 3.549738e-08, 3.549749e-08, 3.549787e-08, 
    3.549816e-08, 3.549788e-08, 3.549758e-08, 3.549678e-08, 3.5496e-08, 
    3.549513e-08, 3.549493e-08, 3.549378e-08, 3.549466e-08, 3.549313e-08, 
    3.549435e-08, 3.549224e-08, 3.549606e-08, 3.549447e-08, 3.549735e-08, 
    3.549706e-08, 3.549649e-08, 3.549524e-08, 3.549597e-08, 3.549513e-08, 
    3.549689e-08, 3.549771e-08, 3.549796e-08, 3.549791e-08, 3.549795e-08, 
    3.549799e-08, 3.54976e-08, 3.549773e-08, 3.549675e-08, 3.549728e-08, 
    3.549575e-08, 3.549515e-08, 3.549344e-08, 3.549232e-08, 3.54912e-08, 
    3.549067e-08, 3.549052e-08, 3.549044e-08,
  6.548689e-11, 6.558122e-11, 6.556294e-11, 6.563884e-11, 6.559682e-11, 
    6.564645e-11, 6.550611e-11, 6.558489e-11, 6.553466e-11, 6.54955e-11, 
    6.578561e-11, 6.564225e-11, 6.593551e-11, 6.584423e-11, 6.607349e-11, 
    6.59212e-11, 6.610418e-11, 6.60693e-11, 6.61747e-11, 6.614453e-11, 
    6.627872e-11, 6.618862e-11, 6.634846e-11, 6.625732e-11, 6.627152e-11, 
    6.618561e-11, 6.567131e-11, 6.576772e-11, 6.566555e-11, 6.567932e-11, 
    6.567318e-11, 6.559762e-11, 6.555938e-11, 6.54798e-11, 6.549429e-11, 
    6.555281e-11, 6.568551e-11, 6.564062e-11, 6.575405e-11, 6.57515e-11, 
    6.587796e-11, 6.582067e-11, 6.603255e-11, 6.597262e-11, 6.61458e-11, 
    6.610227e-11, 6.614372e-11, 6.613118e-11, 6.614388e-11, 6.608004e-11, 
    6.610739e-11, 6.605124e-11, 6.583126e-11, 6.589634e-11, 6.570304e-11, 
    6.558656e-11, 6.550953e-11, 6.545467e-11, 6.546243e-11, 6.547718e-11, 
    6.555315e-11, 6.562465e-11, 6.567903e-11, 6.571534e-11, 6.575113e-11, 
    6.585939e-11, 6.591672e-11, 6.604457e-11, 6.602168e-11, 6.606057e-11, 
    6.609794e-11, 6.61604e-11, 6.615015e-11, 6.617761e-11, 6.605967e-11, 
    6.613802e-11, 6.60086e-11, 6.604401e-11, 6.576021e-11, 6.565277e-11, 
    6.560649e-11, 6.556643e-11, 6.546837e-11, 6.553608e-11, 6.550938e-11, 
    6.5573e-11, 6.561329e-11, 6.55934e-11, 6.571634e-11, 6.566855e-11, 
    6.592012e-11, 6.581158e-11, 6.609359e-11, 6.602639e-11, 6.61097e-11, 
    6.606724e-11, 6.613993e-11, 6.607451e-11, 6.618787e-11, 6.621245e-11, 
    6.619565e-11, 6.626041e-11, 6.607087e-11, 6.614366e-11, 6.559281e-11, 
    6.559605e-11, 6.561122e-11, 6.554447e-11, 6.554042e-11, 6.547936e-11, 
    6.553375e-11, 6.555684e-11, 6.561568e-11, 6.565033e-11, 6.56833e-11, 
    6.575572e-11, 6.583639e-11, 6.594975e-11, 6.603074e-11, 6.608494e-11, 
    6.605176e-11, 6.608105e-11, 6.604828e-11, 6.603294e-11, 6.62032e-11, 
    6.610761e-11, 6.625109e-11, 6.624318e-11, 6.617824e-11, 6.624408e-11, 
    6.559834e-11, 6.557966e-11, 6.551455e-11, 6.556551e-11, 6.547272e-11, 
    6.55246e-11, 6.555435e-11, 6.566941e-11, 6.569481e-11, 6.571815e-11, 
    6.576438e-11, 6.582357e-11, 6.592777e-11, 6.60179e-11, 6.610015e-11, 
    6.609414e-11, 6.609625e-11, 6.611453e-11, 6.606913e-11, 6.612199e-11, 
    6.61308e-11, 6.610767e-11, 6.624212e-11, 6.620375e-11, 6.624302e-11, 
    6.621805e-11, 6.558575e-11, 6.56172e-11, 6.56002e-11, 6.563213e-11, 
    6.560958e-11, 6.57096e-11, 6.573955e-11, 6.588023e-11, 6.582237e-11, 
    6.591428e-11, 6.58317e-11, 6.584677e-11, 6.591698e-11, 6.583674e-11, 
    6.601281e-11, 6.589326e-11, 6.611525e-11, 6.599582e-11, 6.61227e-11, 
    6.609979e-11, 6.613779e-11, 6.617173e-11, 6.621453e-11, 6.629321e-11, 
    6.627503e-11, 6.634087e-11, 6.566412e-11, 6.57048e-11, 6.570134e-11, 
    6.574397e-11, 6.577545e-11, 6.584433e-11, 6.59536e-11, 6.591257e-11, 
    6.5988e-11, 6.600308e-11, 6.588856e-11, 6.595879e-11, 6.57321e-11, 
    6.576857e-11, 6.574695e-11, 6.566726e-11, 6.592186e-11, 6.579099e-11, 
    6.603206e-11, 6.596167e-11, 6.616688e-11, 6.606479e-11, 6.626499e-11, 
    6.635002e-11, 6.64305e-11, 6.652373e-11, 6.572712e-11, 6.569948e-11, 
    6.574907e-11, 6.581739e-11, 6.588161e-11, 6.596594e-11, 6.597463e-11, 
    6.599037e-11, 6.603129e-11, 6.606561e-11, 6.599524e-11, 6.607422e-11, 
    6.577678e-11, 6.593322e-11, 6.568891e-11, 6.576226e-11, 6.581342e-11, 
    6.57911e-11, 6.590791e-11, 6.593524e-11, 6.604607e-11, 6.598887e-11, 
    6.632894e-11, 6.617873e-11, 6.659501e-11, 6.647893e-11, 6.568979e-11, 
    6.572708e-11, 6.585707e-11, 6.579499e-11, 6.597163e-11, 6.601483e-11, 
    6.605004e-11, 6.609481e-11, 6.609973e-11, 6.612625e-11, 6.608277e-11, 
    6.612458e-11, 6.596612e-11, 6.603701e-11, 6.584244e-11, 6.588979e-11, 
    6.586805e-11, 6.584411e-11, 6.591795e-11, 6.599631e-11, 6.599819e-11, 
    6.602325e-11, 6.609348e-11, 6.597235e-11, 6.634793e-11, 6.611595e-11, 
    6.576771e-11, 6.583972e-11, 6.585015e-11, 6.582189e-11, 6.60105e-11, 
    6.594241e-11, 6.612563e-11, 6.607621e-11, 6.615721e-11, 6.611696e-11, 
    6.611103e-11, 6.605932e-11, 6.602706e-11, 6.594549e-11, 6.58791e-11, 
    6.582593e-11, 6.583874e-11, 6.589652e-11, 6.600115e-11, 6.610008e-11, 
    6.60784e-11, 6.615106e-11, 6.595888e-11, 6.603944e-11, 6.600825e-11, 
    6.608958e-11, 6.591144e-11, 6.606258e-11, 6.587267e-11, 6.588939e-11, 
    6.594106e-11, 6.604477e-11, 6.606798e-11, 6.60924e-11, 6.607737e-11, 
    6.600383e-11, 6.599187e-11, 6.593985e-11, 6.592538e-11, 6.588576e-11, 
    6.585285e-11, 6.588288e-11, 6.591434e-11, 6.600395e-11, 6.608446e-11, 
    6.617219e-11, 6.619371e-11, 6.629549e-11, 6.621238e-11, 6.634918e-11, 
    6.623248e-11, 6.643454e-11, 6.607161e-11, 6.622945e-11, 6.594347e-11, 
    6.59744e-11, 6.603009e-11, 6.615802e-11, 6.60892e-11, 6.616977e-11, 
    6.599141e-11, 6.589841e-11, 6.587457e-11, 6.582909e-11, 6.58756e-11, 
    6.587187e-11, 6.591579e-11, 6.590169e-11, 6.600693e-11, 6.595043e-11, 
    6.611083e-11, 6.616919e-11, 6.63339e-11, 6.64345e-11, 6.653703e-11, 
    6.658212e-11, 6.659585e-11, 6.660159e-11,
  3.353199e-14, 3.362921e-14, 3.361035e-14, 3.368868e-14, 3.364528e-14, 
    3.369653e-14, 3.355177e-14, 3.363301e-14, 3.358119e-14, 3.354084e-14, 
    3.384051e-14, 3.369219e-14, 3.399543e-14, 3.390071e-14, 3.413886e-14, 
    3.398059e-14, 3.41708e-14, 3.413446e-14, 3.424425e-14, 3.421281e-14, 
    3.435289e-14, 3.425876e-14, 3.442577e-14, 3.43305e-14, 3.434534e-14, 
    3.425563e-14, 3.372219e-14, 3.382199e-14, 3.371624e-14, 3.373048e-14, 
    3.372413e-14, 3.364612e-14, 3.360672e-14, 3.352467e-14, 3.353959e-14, 
    3.359991e-14, 3.373689e-14, 3.369049e-14, 3.380773e-14, 3.380509e-14, 
    3.393568e-14, 3.387671e-14, 3.409623e-14, 3.403392e-14, 3.421412e-14, 
    3.416878e-14, 3.421196e-14, 3.419889e-14, 3.421213e-14, 3.414564e-14, 
    3.417412e-14, 3.411566e-14, 3.388769e-14, 3.395475e-14, 3.375499e-14, 
    3.363476e-14, 3.355531e-14, 3.349881e-14, 3.350679e-14, 3.352199e-14, 
    3.360027e-14, 3.3674e-14, 3.373016e-14, 3.37677e-14, 3.380471e-14, 
    3.391649e-14, 3.397593e-14, 3.410875e-14, 3.408492e-14, 3.41254e-14, 
    3.416427e-14, 3.422935e-14, 3.421866e-14, 3.424729e-14, 3.412443e-14, 
    3.420604e-14, 3.407131e-14, 3.410814e-14, 3.381423e-14, 3.370303e-14, 
    3.365531e-14, 3.361395e-14, 3.351292e-14, 3.358266e-14, 3.355516e-14, 
    3.362071e-14, 3.366229e-14, 3.364174e-14, 3.376872e-14, 3.371933e-14, 
    3.397945e-14, 3.386731e-14, 3.415974e-14, 3.408982e-14, 3.417652e-14, 
    3.41323e-14, 3.420802e-14, 3.413988e-14, 3.4258e-14, 3.428366e-14, 
    3.426611e-14, 3.433369e-14, 3.413609e-14, 3.421191e-14, 3.364114e-14, 
    3.364449e-14, 3.366014e-14, 3.359132e-14, 3.358714e-14, 3.352424e-14, 
    3.358026e-14, 3.360407e-14, 3.366474e-14, 3.370052e-14, 3.373458e-14, 
    3.380947e-14, 3.389303e-14, 3.40102e-14, 3.409435e-14, 3.415073e-14, 
    3.411619e-14, 3.414668e-14, 3.411258e-14, 3.409662e-14, 3.427401e-14, 
    3.417435e-14, 3.432397e-14, 3.431571e-14, 3.424795e-14, 3.431665e-14, 
    3.364685e-14, 3.362757e-14, 3.356047e-14, 3.361298e-14, 3.351739e-14, 
    3.357083e-14, 3.360152e-14, 3.372025e-14, 3.374647e-14, 3.377061e-14, 
    3.381842e-14, 3.387972e-14, 3.398738e-14, 3.4081e-14, 3.416656e-14, 
    3.41603e-14, 3.41625e-14, 3.418155e-14, 3.413428e-14, 3.418932e-14, 
    3.41985e-14, 3.41744e-14, 3.43146e-14, 3.427455e-14, 3.431553e-14, 
    3.428948e-14, 3.363385e-14, 3.366631e-14, 3.364876e-14, 3.368173e-14, 
    3.365846e-14, 3.376179e-14, 3.379277e-14, 3.393807e-14, 3.387848e-14, 
    3.397338e-14, 3.388814e-14, 3.390335e-14, 3.397624e-14, 3.389294e-14, 
    3.407574e-14, 3.39516e-14, 3.418229e-14, 3.40581e-14, 3.419006e-14, 
    3.416619e-14, 3.420578e-14, 3.424117e-14, 3.42858e-14, 3.436799e-14, 
    3.434899e-14, 3.441781e-14, 3.371476e-14, 3.375682e-14, 3.375321e-14, 
    3.37973e-14, 3.382989e-14, 3.390081e-14, 3.401418e-14, 3.397158e-14, 
    3.40499e-14, 3.406559e-14, 3.394666e-14, 3.401958e-14, 3.378504e-14, 
    3.38228e-14, 3.38004e-14, 3.371802e-14, 3.398125e-14, 3.384601e-14, 
    3.409572e-14, 3.402256e-14, 3.423611e-14, 3.41298e-14, 3.43385e-14, 
    3.442744e-14, 3.451163e-14, 3.460945e-14, 3.377988e-14, 3.375129e-14, 
    3.380258e-14, 3.387335e-14, 3.393947e-14, 3.4027e-14, 3.403601e-14, 
    3.405238e-14, 3.409491e-14, 3.413061e-14, 3.405746e-14, 3.413957e-14, 
    3.383135e-14, 3.399303e-14, 3.374039e-14, 3.381627e-14, 3.386922e-14, 
    3.384609e-14, 3.396674e-14, 3.39951e-14, 3.411031e-14, 3.405081e-14, 
    3.440539e-14, 3.42485e-14, 3.468428e-14, 3.456244e-14, 3.374128e-14, 
    3.377983e-14, 3.391404e-14, 3.385011e-14, 3.40329e-14, 3.407781e-14, 
    3.41144e-14, 3.416102e-14, 3.416613e-14, 3.419376e-14, 3.414847e-14, 
    3.419201e-14, 3.402718e-14, 3.410086e-14, 3.389884e-14, 3.394795e-14, 
    3.392539e-14, 3.390057e-14, 3.397716e-14, 3.405858e-14, 3.406049e-14, 
    3.408657e-14, 3.415977e-14, 3.403364e-14, 3.442534e-14, 3.418314e-14, 
    3.382187e-14, 3.389607e-14, 3.390685e-14, 3.387797e-14, 3.40733e-14, 
    3.400256e-14, 3.419311e-14, 3.414164e-14, 3.422602e-14, 3.418408e-14, 
    3.41779e-14, 3.412407e-14, 3.409051e-14, 3.400577e-14, 3.393687e-14, 
    3.388215e-14, 3.389501e-14, 3.395494e-14, 3.40636e-14, 3.416652e-14, 
    3.414395e-14, 3.421961e-14, 3.401965e-14, 3.410341e-14, 3.407098e-14, 
    3.415556e-14, 3.397041e-14, 3.412757e-14, 3.393018e-14, 3.394752e-14, 
    3.400116e-14, 3.410898e-14, 3.413308e-14, 3.415851e-14, 3.414285e-14, 
    3.406639e-14, 3.405394e-14, 3.399989e-14, 3.398489e-14, 3.394376e-14, 
    3.390963e-14, 3.394077e-14, 3.397344e-14, 3.406649e-14, 3.415026e-14, 
    3.424165e-14, 3.426408e-14, 3.437044e-14, 3.428363e-14, 3.442665e-14, 
    3.430471e-14, 3.451597e-14, 3.413693e-14, 3.430146e-14, 3.400365e-14, 
    3.403577e-14, 3.40937e-14, 3.422691e-14, 3.415517e-14, 3.423915e-14, 
    3.405346e-14, 3.395693e-14, 3.393216e-14, 3.388544e-14, 3.393322e-14, 
    3.392935e-14, 3.397491e-14, 3.396028e-14, 3.406958e-14, 3.401088e-14, 
    3.41777e-14, 3.423853e-14, 3.441053e-14, 3.451587e-14, 3.462336e-14, 
    3.467072e-14, 3.468515e-14, 3.469117e-14,
  5.203943e-18, 5.226065e-18, 5.221734e-18, 5.239728e-18, 5.229756e-18, 
    5.241533e-18, 5.208395e-18, 5.226939e-18, 5.215042e-18, 5.205932e-18, 
    5.274674e-18, 5.240535e-18, 5.310368e-18, 5.288511e-18, 5.343519e-18, 
    5.306946e-18, 5.350911e-18, 5.342495e-18, 5.367917e-18, 5.360632e-18, 
    5.393124e-18, 5.37128e-18, 5.410047e-18, 5.387922e-18, 5.391369e-18, 
    5.370555e-18, 5.247429e-18, 5.270409e-18, 5.246061e-18, 5.249337e-18, 
    5.247875e-18, 5.22995e-18, 5.220906e-18, 5.202291e-18, 5.205652e-18, 
    5.219341e-18, 5.250811e-18, 5.240142e-18, 5.267109e-18, 5.266501e-18, 
    5.296575e-18, 5.282999e-18, 5.333654e-18, 5.31925e-18, 5.360936e-18, 
    5.350437e-18, 5.360437e-18, 5.357409e-18, 5.360477e-18, 5.345083e-18, 
    5.351675e-18, 5.338147e-18, 5.285532e-18, 5.300975e-18, 5.254975e-18, 
    5.227347e-18, 5.209192e-18, 5.196469e-18, 5.198266e-18, 5.201688e-18, 
    5.219422e-18, 5.236352e-18, 5.249259e-18, 5.257895e-18, 5.266413e-18, 
    5.292158e-18, 5.305866e-18, 5.336552e-18, 5.331036e-18, 5.340402e-18, 
    5.349394e-18, 5.364466e-18, 5.361988e-18, 5.368625e-18, 5.340175e-18, 
    5.359067e-18, 5.327889e-18, 5.336407e-18, 5.268621e-18, 5.243024e-18, 
    5.232066e-18, 5.222563e-18, 5.199647e-18, 5.215382e-18, 5.20916e-18, 
    5.22411e-18, 5.23366e-18, 5.228941e-18, 5.258131e-18, 5.246771e-18, 
    5.306678e-18, 5.280837e-18, 5.348345e-18, 5.332171e-18, 5.352228e-18, 
    5.341996e-18, 5.359524e-18, 5.343748e-18, 5.371105e-18, 5.377056e-18, 
    5.372986e-18, 5.388661e-18, 5.342871e-18, 5.360427e-18, 5.228803e-18, 
    5.229572e-18, 5.233167e-18, 5.217369e-18, 5.216409e-18, 5.202193e-18, 
    5.214827e-18, 5.220294e-18, 5.234222e-18, 5.242447e-18, 5.250277e-18, 
    5.267511e-18, 5.286764e-18, 5.313775e-18, 5.333217e-18, 5.346259e-18, 
    5.338268e-18, 5.345322e-18, 5.337433e-18, 5.333741e-18, 5.374819e-18, 
    5.35173e-18, 5.386405e-18, 5.384488e-18, 5.368779e-18, 5.384704e-18, 
    5.230114e-18, 5.225686e-18, 5.210356e-18, 5.222338e-18, 5.200652e-18, 
    5.21269e-18, 5.219711e-18, 5.246985e-18, 5.25301e-18, 5.258566e-18, 
    5.269571e-18, 5.283692e-18, 5.308506e-18, 5.330134e-18, 5.349922e-18, 
    5.348473e-18, 5.348982e-18, 5.353395e-18, 5.342452e-18, 5.355193e-18, 
    5.357322e-18, 5.35174e-18, 5.384231e-18, 5.374943e-18, 5.384447e-18, 
    5.378402e-18, 5.227128e-18, 5.234585e-18, 5.230553e-18, 5.23813e-18, 
    5.232783e-18, 5.256541e-18, 5.263672e-18, 5.29713e-18, 5.283408e-18, 
    5.305274e-18, 5.285635e-18, 5.289118e-18, 5.305942e-18, 5.286716e-18, 
    5.32892e-18, 5.300253e-18, 5.353566e-18, 5.324848e-18, 5.355365e-18, 
    5.349836e-18, 5.359003e-18, 5.367205e-18, 5.377551e-18, 5.396626e-18, 
    5.392211e-18, 5.408195e-18, 5.245719e-18, 5.255394e-18, 5.254562e-18, 
    5.264709e-18, 5.272213e-18, 5.28853e-18, 5.314693e-18, 5.304855e-18, 
    5.322942e-18, 5.326569e-18, 5.299105e-18, 5.315942e-18, 5.261889e-18, 
    5.270585e-18, 5.265422e-18, 5.24647e-18, 5.307094e-18, 5.27593e-18, 
    5.333535e-18, 5.316626e-18, 5.366033e-18, 5.34142e-18, 5.389777e-18, 
    5.410441e-18, 5.430011e-18, 5.452797e-18, 5.2607e-18, 5.25412e-18, 
    5.265922e-18, 5.282229e-18, 5.297447e-18, 5.317653e-18, 5.319733e-18, 
    5.323516e-18, 5.333345e-18, 5.341604e-18, 5.324693e-18, 5.343677e-18, 
    5.272562e-18, 5.30981e-18, 5.251615e-18, 5.269082e-18, 5.281276e-18, 
    5.275946e-18, 5.303737e-18, 5.310284e-18, 5.336911e-18, 5.323152e-18, 
    5.40532e-18, 5.368909e-18, 5.470238e-18, 5.441843e-18, 5.251817e-18, 
    5.260687e-18, 5.291584e-18, 5.276871e-18, 5.319014e-18, 5.329394e-18, 
    5.337854e-18, 5.348643e-18, 5.349824e-18, 5.356223e-18, 5.345736e-18, 
    5.355817e-18, 5.317696e-18, 5.334722e-18, 5.288075e-18, 5.299403e-18, 
    5.294198e-18, 5.288475e-18, 5.306142e-18, 5.324954e-18, 5.325389e-18, 
    5.331421e-18, 5.348372e-18, 5.319186e-18, 5.409964e-18, 5.353781e-18, 
    5.270363e-18, 5.287444e-18, 5.289923e-18, 5.283288e-18, 5.328351e-18, 
    5.312008e-18, 5.356072e-18, 5.344157e-18, 5.363693e-18, 5.353979e-18, 
    5.352549e-18, 5.340091e-18, 5.332331e-18, 5.312751e-18, 5.296848e-18, 
    5.284252e-18, 5.287193e-18, 5.301018e-18, 5.326113e-18, 5.349916e-18, 
    5.344694e-18, 5.362207e-18, 5.315954e-18, 5.335315e-18, 5.327818e-18, 
    5.347379e-18, 5.304587e-18, 5.340919e-18, 5.295303e-18, 5.299303e-18, 
    5.311684e-18, 5.336606e-18, 5.342175e-18, 5.348063e-18, 5.344436e-18, 
    5.326757e-18, 5.323877e-18, 5.311391e-18, 5.307929e-18, 5.298435e-18, 
    5.290563e-18, 5.297747e-18, 5.305288e-18, 5.326778e-18, 5.346153e-18, 
    5.367317e-18, 5.372514e-18, 5.397204e-18, 5.377057e-18, 5.410271e-18, 
    5.381959e-18, 5.431036e-18, 5.343076e-18, 5.381194e-18, 5.312259e-18, 
    5.319678e-18, 5.333072e-18, 5.363907e-18, 5.347287e-18, 5.366742e-18, 
    5.323767e-18, 5.301479e-18, 5.295758e-18, 5.285011e-18, 5.296004e-18, 
    5.295112e-18, 5.305623e-18, 5.302247e-18, 5.327492e-18, 5.313927e-18, 
    5.352504e-18, 5.366597e-18, 5.406507e-18, 5.431002e-18, 5.456029e-18, 
    5.467072e-18, 5.470438e-18, 5.471844e-18,
  2.57918e-22, 2.593651e-22, 2.590815e-22, 2.602603e-22, 2.596067e-22, 
    2.603786e-22, 2.582088e-22, 2.594225e-22, 2.586434e-22, 2.580478e-22, 
    2.625542e-22, 2.603132e-22, 2.649261e-22, 2.634686e-22, 2.671406e-22, 
    2.64698e-22, 2.676349e-22, 2.670717e-22, 2.68773e-22, 2.682851e-22, 
    2.704638e-22, 2.689983e-22, 2.715997e-22, 2.701144e-22, 2.703458e-22, 
    2.689498e-22, 2.60765e-22, 2.622741e-22, 2.606753e-22, 2.608903e-22, 
    2.607942e-22, 2.596196e-22, 2.590276e-22, 2.578098e-22, 2.580295e-22, 
    2.589249e-22, 2.60987e-22, 2.602871e-22, 2.620563e-22, 2.620163e-22, 
    2.640059e-22, 2.631019e-22, 2.664806e-22, 2.655184e-22, 2.683055e-22, 
    2.676028e-22, 2.682721e-22, 2.680693e-22, 2.682748e-22, 2.672448e-22, 
    2.676857e-22, 2.667809e-22, 2.632707e-22, 2.642994e-22, 2.6126e-22, 
    2.594496e-22, 2.58261e-22, 2.574295e-22, 2.57547e-22, 2.577706e-22, 
    2.589302e-22, 2.600388e-22, 2.608849e-22, 2.614514e-22, 2.620105e-22, 
    2.637123e-22, 2.646258e-22, 2.666745e-22, 2.663057e-22, 2.669319e-22, 
    2.675331e-22, 2.685419e-22, 2.68376e-22, 2.688206e-22, 2.669165e-22, 
    2.681806e-22, 2.660953e-22, 2.666646e-22, 2.621568e-22, 2.604761e-22, 
    2.597586e-22, 2.591358e-22, 2.576372e-22, 2.586658e-22, 2.582589e-22, 
    2.592369e-22, 2.598624e-22, 2.595532e-22, 2.614669e-22, 2.607218e-22, 
    2.6468e-22, 2.629584e-22, 2.674629e-22, 2.663815e-22, 2.677227e-22, 
    2.670381e-22, 2.682111e-22, 2.671553e-22, 2.689866e-22, 2.693856e-22, 
    2.691128e-22, 2.701636e-22, 2.670967e-22, 2.682716e-22, 2.595442e-22, 
    2.595946e-22, 2.598301e-22, 2.587958e-22, 2.587329e-22, 2.578035e-22, 
    2.586294e-22, 2.589872e-22, 2.598991e-22, 2.604383e-22, 2.609518e-22, 
    2.620828e-22, 2.63353e-22, 2.651533e-22, 2.664514e-22, 2.673233e-22, 
    2.667889e-22, 2.672606e-22, 2.667331e-22, 2.664863e-22, 2.692357e-22, 
    2.676895e-22, 2.700123e-22, 2.698837e-22, 2.688309e-22, 2.698982e-22, 
    2.596301e-22, 2.593401e-22, 2.58337e-22, 2.591208e-22, 2.577028e-22, 
    2.584897e-22, 2.589492e-22, 2.607361e-22, 2.61131e-22, 2.614956e-22, 
    2.622179e-22, 2.631481e-22, 2.648016e-22, 2.662456e-22, 2.675683e-22, 
    2.674714e-22, 2.675054e-22, 2.678008e-22, 2.670687e-22, 2.679211e-22, 
    2.680637e-22, 2.6769e-22, 2.698665e-22, 2.692438e-22, 2.69881e-22, 
    2.694756e-22, 2.594345e-22, 2.59923e-22, 2.596589e-22, 2.601553e-22, 
    2.598051e-22, 2.61363e-22, 2.618311e-22, 2.640433e-22, 2.631292e-22, 
    2.645861e-22, 2.632775e-22, 2.635091e-22, 2.646313e-22, 2.633488e-22, 
    2.661647e-22, 2.642516e-22, 2.678122e-22, 2.658931e-22, 2.679326e-22, 
    2.675626e-22, 2.68176e-22, 2.687254e-22, 2.694186e-22, 2.706984e-22, 
    2.70402e-22, 2.714751e-22, 2.606527e-22, 2.612876e-22, 2.612327e-22, 
    2.618987e-22, 2.623916e-22, 2.634697e-22, 2.652144e-22, 2.645579e-22, 
    2.657649e-22, 2.660072e-22, 2.641744e-22, 2.652979e-22, 2.617138e-22, 
    2.62285e-22, 2.619456e-22, 2.607022e-22, 2.647076e-22, 2.626361e-22, 
    2.664727e-22, 2.653434e-22, 2.686469e-22, 2.670001e-22, 2.702386e-22, 
    2.716266e-22, 2.729416e-22, 2.744764e-22, 2.616356e-22, 2.612037e-22, 
    2.619783e-22, 2.63051e-22, 2.640641e-22, 2.65412e-22, 2.655507e-22, 
    2.658034e-22, 2.664599e-22, 2.670119e-22, 2.658822e-22, 2.671506e-22, 
    2.624154e-22, 2.648887e-22, 2.610395e-22, 2.621863e-22, 2.629874e-22, 
    2.626368e-22, 2.644832e-22, 2.6492e-22, 2.666985e-22, 2.65779e-22, 
    2.712827e-22, 2.6884e-22, 2.756519e-22, 2.737384e-22, 2.610527e-22, 
    2.616346e-22, 2.636735e-22, 2.626976e-22, 2.655027e-22, 2.66196e-22, 
    2.667612e-22, 2.674829e-22, 2.675618e-22, 2.679901e-22, 2.672883e-22, 
    2.679628e-22, 2.654148e-22, 2.66552e-22, 2.634393e-22, 2.641944e-22, 
    2.638473e-22, 2.63466e-22, 2.646437e-22, 2.658997e-22, 2.659284e-22, 
    2.663315e-22, 2.674662e-22, 2.655141e-22, 2.715954e-22, 2.678279e-22, 
    2.622699e-22, 2.633979e-22, 2.635626e-22, 2.63121e-22, 2.661263e-22, 
    2.650352e-22, 2.679799e-22, 2.671827e-22, 2.684901e-22, 2.678398e-22, 
    2.677441e-22, 2.669108e-22, 2.663922e-22, 2.650848e-22, 2.640241e-22, 
    2.631852e-22, 2.633806e-22, 2.643022e-22, 2.659771e-22, 2.675681e-22, 
    2.672189e-22, 2.683906e-22, 2.652984e-22, 2.665917e-22, 2.660909e-22, 
    2.673982e-22, 2.645401e-22, 2.669675e-22, 2.639209e-22, 2.641876e-22, 
    2.650135e-22, 2.666784e-22, 2.670501e-22, 2.674441e-22, 2.672014e-22, 
    2.6602e-22, 2.658275e-22, 2.649939e-22, 2.647631e-22, 2.641297e-22, 
    2.636051e-22, 2.640839e-22, 2.64587e-22, 2.660212e-22, 2.673164e-22, 
    2.68733e-22, 2.69081e-22, 2.707379e-22, 2.693862e-22, 2.716161e-22, 
    2.697159e-22, 2.730118e-22, 2.671112e-22, 2.696638e-22, 2.650518e-22, 
    2.65547e-22, 2.664421e-22, 2.68505e-22, 2.673921e-22, 2.686948e-22, 
    2.658201e-22, 2.643331e-22, 2.639513e-22, 2.632358e-22, 2.639677e-22, 
    2.639083e-22, 2.64609e-22, 2.643838e-22, 2.660689e-22, 2.651631e-22, 
    2.677412e-22, 2.686849e-22, 2.713619e-22, 2.730088e-22, 2.746936e-22, 
    2.754382e-22, 2.756652e-22, 2.7576e-22,
  4.169368e-27, 4.198372e-27, 4.192702e-27, 4.216297e-27, 4.203196e-27, 
    4.218689e-27, 4.175216e-27, 4.199521e-27, 4.183952e-27, 4.171975e-27, 
    4.262769e-27, 4.217365e-27, 4.310965e-27, 4.28131e-27, 4.356103e-27, 
    4.306325e-27, 4.366193e-27, 4.354691e-27, 4.38944e-27, 4.379468e-27, 
    4.424059e-27, 4.394049e-27, 4.447339e-27, 4.416895e-27, 4.421637e-27, 
    4.393057e-27, 4.226502e-27, 4.257089e-27, 4.224688e-27, 4.229041e-27, 
    4.227093e-27, 4.203456e-27, 4.191633e-27, 4.167187e-27, 4.171606e-27, 
    4.189578e-27, 4.231e-27, 4.216834e-27, 4.252651e-27, 4.25184e-27, 
    4.292234e-27, 4.27386e-27, 4.342632e-27, 4.323018e-27, 4.379884e-27, 
    4.365532e-27, 4.379205e-27, 4.37506e-27, 4.379259e-27, 4.358223e-27, 
    4.367226e-27, 4.348756e-27, 4.277292e-27, 4.298205e-27, 4.236525e-27, 
    4.200068e-27, 4.176267e-27, 4.15954e-27, 4.161902e-27, 4.166402e-27, 
    4.189683e-27, 4.211835e-27, 4.228927e-27, 4.240397e-27, 4.251724e-27, 
    4.286277e-27, 4.304852e-27, 4.346592e-27, 4.339063e-27, 4.351841e-27, 
    4.364107e-27, 4.38472e-27, 4.381326e-27, 4.390418e-27, 4.351521e-27, 
    4.377337e-27, 4.334773e-27, 4.346383e-27, 4.254713e-27, 4.220657e-27, 
    4.206243e-27, 4.193788e-27, 4.163717e-27, 4.184402e-27, 4.176226e-27, 
    4.195806e-27, 4.208308e-27, 4.202125e-27, 4.240711e-27, 4.225627e-27, 
    4.305954e-27, 4.270948e-27, 4.362675e-27, 4.340609e-27, 4.367979e-27, 
    4.354003e-27, 4.37796e-27, 4.356395e-27, 4.393812e-27, 4.401978e-27, 
    4.396395e-27, 4.417899e-27, 4.355199e-27, 4.379196e-27, 4.201948e-27, 
    4.202955e-27, 4.207661e-27, 4.186999e-27, 4.185743e-27, 4.167061e-27, 
    4.183672e-27, 4.19082e-27, 4.209041e-27, 4.219892e-27, 4.230282e-27, 
    4.25319e-27, 4.278967e-27, 4.315586e-27, 4.342036e-27, 4.359824e-27, 
    4.348917e-27, 4.358544e-27, 4.34778e-27, 4.342744e-27, 4.39891e-27, 
    4.367305e-27, 4.414801e-27, 4.412168e-27, 4.39063e-27, 4.412464e-27, 
    4.203664e-27, 4.197866e-27, 4.177797e-27, 4.193486e-27, 4.165035e-27, 
    4.18087e-27, 4.190064e-27, 4.225922e-27, 4.233909e-27, 4.241294e-27, 
    4.255929e-27, 4.274799e-27, 4.308426e-27, 4.337841e-27, 4.364825e-27, 
    4.362846e-27, 4.363542e-27, 4.369575e-27, 4.354629e-27, 4.372032e-27, 
    4.374949e-27, 4.367312e-27, 4.411814e-27, 4.399071e-27, 4.412111e-27, 
    4.403813e-27, 4.199752e-27, 4.209519e-27, 4.204238e-27, 4.21417e-27, 
    4.207163e-27, 4.238614e-27, 4.248097e-27, 4.293e-27, 4.274417e-27, 
    4.304041e-27, 4.277427e-27, 4.282132e-27, 4.30497e-27, 4.278872e-27, 
    4.336197e-27, 4.297241e-27, 4.369809e-27, 4.330665e-27, 4.372268e-27, 
    4.364708e-27, 4.377239e-27, 4.388471e-27, 4.402648e-27, 4.428858e-27, 
    4.422784e-27, 4.444779e-27, 4.22423e-27, 4.237084e-27, 4.235969e-27, 
    4.249459e-27, 4.259451e-27, 4.281329e-27, 4.316827e-27, 4.303461e-27, 
    4.32804e-27, 4.33298e-27, 4.295657e-27, 4.318529e-27, 4.245715e-27, 
    4.257296e-27, 4.250411e-27, 4.225233e-27, 4.306514e-27, 4.264414e-27, 
    4.342471e-27, 4.319453e-27, 4.386866e-27, 4.353234e-27, 4.419438e-27, 
    4.447897e-27, 4.474879e-27, 4.506449e-27, 4.24413e-27, 4.235381e-27, 
    4.25107e-27, 4.272832e-27, 4.293416e-27, 4.320851e-27, 4.323675e-27, 
    4.328825e-27, 4.342206e-27, 4.353469e-27, 4.330437e-27, 4.356298e-27, 
    4.25995e-27, 4.310198e-27, 4.23206e-27, 4.255298e-27, 4.271538e-27, 
    4.264424e-27, 4.301939e-27, 4.31083e-27, 4.347079e-27, 4.328325e-27, 
    4.440845e-27, 4.390821e-27, 4.530648e-27, 4.491265e-27, 4.232323e-27, 
    4.244108e-27, 4.285476e-27, 4.265655e-27, 4.322697e-27, 4.336827e-27, 
    4.348353e-27, 4.363087e-27, 4.364693e-27, 4.373443e-27, 4.359108e-27, 
    4.372883e-27, 4.32091e-27, 4.344086e-27, 4.280711e-27, 4.296068e-27, 
    4.289004e-27, 4.281252e-27, 4.305205e-27, 4.330794e-27, 4.331371e-27, 
    4.339594e-27, 4.36277e-27, 4.32293e-27, 4.447276e-27, 4.370153e-27, 
    4.256982e-27, 4.279878e-27, 4.283219e-27, 4.274247e-27, 4.335408e-27, 
    4.313177e-27, 4.373234e-27, 4.356954e-27, 4.383657e-27, 4.370371e-27, 
    4.368417e-27, 4.351405e-27, 4.340828e-27, 4.314189e-27, 4.292604e-27, 
    4.275551e-27, 4.279516e-27, 4.29826e-27, 4.33237e-27, 4.364825e-27, 
    4.357698e-27, 4.381624e-27, 4.318537e-27, 4.344901e-27, 4.334689e-27, 
    4.361355e-27, 4.303099e-27, 4.352587e-27, 4.290501e-27, 4.295927e-27, 
    4.312737e-27, 4.346673e-27, 4.354248e-27, 4.362294e-27, 4.357334e-27, 
    4.333243e-27, 4.329318e-27, 4.312334e-27, 4.307639e-27, 4.294747e-27, 
    4.28408e-27, 4.293818e-27, 4.304056e-27, 4.333265e-27, 4.359687e-27, 
    4.388627e-27, 4.39574e-27, 4.429682e-27, 4.401999e-27, 4.447702e-27, 
    4.408766e-27, 4.476343e-27, 4.355509e-27, 4.407682e-27, 4.313512e-27, 
    4.323599e-27, 4.341852e-27, 4.383974e-27, 4.36123e-27, 4.387851e-27, 
    4.329166e-27, 4.298894e-27, 4.29112e-27, 4.276581e-27, 4.291453e-27, 
    4.290244e-27, 4.3045e-27, 4.299917e-27, 4.334238e-27, 4.31578e-27, 
    4.368361e-27, 4.387648e-27, 4.44246e-27, 4.476268e-27, 4.510908e-27, 
    4.526241e-27, 4.530918e-27, 4.532872e-27,
  2.174826e-32, 2.193216e-32, 2.189626e-32, 2.204576e-32, 2.19627e-32, 
    2.206095e-32, 2.17854e-32, 2.193945e-32, 2.184089e-32, 2.176481e-32, 
    2.234141e-32, 2.205254e-32, 2.264944e-32, 2.245911e-32, 2.293989e-32, 
    2.261965e-32, 2.300493e-32, 2.293074e-32, 2.315497e-32, 2.309056e-32, 
    2.3379e-32, 2.318475e-32, 2.352991e-32, 2.333257e-32, 2.33633e-32, 
    2.317834e-32, 2.211056e-32, 2.230524e-32, 2.209904e-32, 2.212672e-32, 
    2.211432e-32, 2.196436e-32, 2.188953e-32, 2.173439e-32, 2.176246e-32, 
    2.18765e-32, 2.213917e-32, 2.204915e-32, 2.227686e-32, 2.22717e-32, 
    2.252916e-32, 2.241189e-32, 2.285307e-32, 2.272685e-32, 2.309325e-32, 
    2.300063e-32, 2.308887e-32, 2.30621e-32, 2.308922e-32, 2.295352e-32, 
    2.301157e-32, 2.28925e-32, 2.243364e-32, 2.256748e-32, 2.217428e-32, 
    2.194295e-32, 2.179209e-32, 2.168585e-32, 2.170084e-32, 2.172942e-32, 
    2.187717e-32, 2.201743e-32, 2.212596e-32, 2.219889e-32, 2.227096e-32, 
    2.249103e-32, 2.261018e-32, 2.287859e-32, 2.283008e-32, 2.29124e-32, 
    2.299144e-32, 2.312448e-32, 2.310256e-32, 2.31613e-32, 2.291031e-32, 
    2.307683e-32, 2.280245e-32, 2.287722e-32, 2.229012e-32, 2.207342e-32, 
    2.198205e-32, 2.190314e-32, 2.171237e-32, 2.184375e-32, 2.179184e-32, 
    2.191589e-32, 2.199508e-32, 2.195591e-32, 2.220089e-32, 2.2105e-32, 
    2.261725e-32, 2.239345e-32, 2.298221e-32, 2.284004e-32, 2.301641e-32, 
    2.29263e-32, 2.308084e-32, 2.294172e-32, 2.318323e-32, 2.323604e-32, 
    2.319993e-32, 2.333904e-32, 2.293401e-32, 2.308882e-32, 2.195479e-32, 
    2.196117e-32, 2.199097e-32, 2.186019e-32, 2.185223e-32, 2.17336e-32, 
    2.183912e-32, 2.188436e-32, 2.199971e-32, 2.206857e-32, 2.213459e-32, 
    2.228031e-32, 2.244427e-32, 2.267911e-32, 2.284923e-32, 2.296382e-32, 
    2.289353e-32, 2.295557e-32, 2.28862e-32, 2.285377e-32, 2.321621e-32, 
    2.301208e-32, 2.331899e-32, 2.330194e-32, 2.316268e-32, 2.330386e-32, 
    2.196566e-32, 2.192893e-32, 2.180181e-32, 2.190121e-32, 2.172073e-32, 
    2.182135e-32, 2.187959e-32, 2.21069e-32, 2.215763e-32, 2.220461e-32, 
    2.229774e-32, 2.241783e-32, 2.26331e-32, 2.282223e-32, 2.299607e-32, 
    2.29833e-32, 2.298779e-32, 2.302671e-32, 2.293034e-32, 2.304257e-32, 
    2.306141e-32, 2.301212e-32, 2.329965e-32, 2.321722e-32, 2.330158e-32, 
    2.324788e-32, 2.194088e-32, 2.200275e-32, 2.196929e-32, 2.203224e-32, 
    2.198783e-32, 2.218759e-32, 2.224793e-32, 2.253411e-32, 2.241542e-32, 
    2.260495e-32, 2.243449e-32, 2.246438e-32, 2.261097e-32, 2.244362e-32, 
    2.281168e-32, 2.256134e-32, 2.302823e-32, 2.277612e-32, 2.304409e-32, 
    2.299531e-32, 2.307616e-32, 2.314872e-32, 2.324035e-32, 2.341006e-32, 
    2.337069e-32, 2.351328e-32, 2.209612e-32, 2.217784e-32, 2.217073e-32, 
    2.225655e-32, 2.232017e-32, 2.245922e-32, 2.268707e-32, 2.26012e-32, 
    2.275915e-32, 2.279093e-32, 2.25511e-32, 2.269802e-32, 2.223274e-32, 
    2.230648e-32, 2.226262e-32, 2.210251e-32, 2.262084e-32, 2.235182e-32, 
    2.285203e-32, 2.270394e-32, 2.313835e-32, 2.292138e-32, 2.334902e-32, 
    2.353357e-32, 2.370877e-32, 2.391436e-32, 2.222264e-32, 2.216699e-32, 
    2.22668e-32, 2.24054e-32, 2.253674e-32, 2.271294e-32, 2.273108e-32, 
    2.27642e-32, 2.285031e-32, 2.292286e-32, 2.27746e-32, 2.294109e-32, 
    2.232344e-32, 2.264449e-32, 2.214589e-32, 2.229376e-32, 2.239719e-32, 
    2.235185e-32, 2.259142e-32, 2.264852e-32, 2.288172e-32, 2.276098e-32, 
    2.348783e-32, 2.316394e-32, 2.407219e-32, 2.381543e-32, 2.214755e-32, 
    2.222249e-32, 2.248583e-32, 2.235969e-32, 2.272479e-32, 2.281569e-32, 
    2.288989e-32, 2.298488e-32, 2.299522e-32, 2.305168e-32, 2.295921e-32, 
    2.304806e-32, 2.271331e-32, 2.286242e-32, 2.245527e-32, 2.255375e-32, 
    2.250842e-32, 2.245872e-32, 2.261239e-32, 2.277691e-32, 2.278058e-32, 
    2.283351e-32, 2.298297e-32, 2.272628e-32, 2.352963e-32, 2.303057e-32, 
    2.230444e-32, 2.245005e-32, 2.247134e-32, 2.241433e-32, 2.280656e-32, 
    2.266361e-32, 2.305032e-32, 2.294531e-32, 2.311761e-32, 2.303185e-32, 
    2.301925e-32, 2.290956e-32, 2.284145e-32, 2.267012e-32, 2.253153e-32, 
    2.242258e-32, 2.24477e-32, 2.256783e-32, 2.278703e-32, 2.299609e-32, 
    2.295014e-32, 2.310448e-32, 2.269805e-32, 2.286769e-32, 2.280195e-32, 
    2.29737e-32, 2.259889e-32, 2.291731e-32, 2.251803e-32, 2.255283e-32, 
    2.266078e-32, 2.287913e-32, 2.292788e-32, 2.297977e-32, 2.294777e-32, 
    2.279265e-32, 2.276738e-32, 2.265819e-32, 2.262804e-32, 2.254526e-32, 
    2.247685e-32, 2.253931e-32, 2.260504e-32, 2.279277e-32, 2.296296e-32, 
    2.314973e-32, 2.319568e-32, 2.341547e-32, 2.323623e-32, 2.353241e-32, 
    2.32801e-32, 2.371842e-32, 2.293608e-32, 2.327301e-32, 2.266575e-32, 
    2.273058e-32, 2.284807e-32, 2.311972e-32, 2.297289e-32, 2.314475e-32, 
    2.27664e-32, 2.257192e-32, 2.2522e-32, 2.242912e-32, 2.252413e-32, 
    2.251637e-32, 2.260786e-32, 2.257844e-32, 2.279903e-32, 2.268033e-32, 
    2.301889e-32, 2.314342e-32, 2.349825e-32, 2.371786e-32, 2.394336e-32, 
    2.40434e-32, 2.407393e-32, 2.408669e-32,
  3.736255e-38, 3.775949e-38, 3.768196e-38, 3.800503e-38, 3.782544e-38, 
    3.803774e-38, 3.744268e-38, 3.777527e-38, 3.756251e-38, 3.73982e-38, 
    3.864394e-38, 3.801962e-38, 3.931198e-38, 3.889861e-38, 3.994617e-38, 
    3.924721e-38, 4.009003e-38, 3.992606e-38, 4.042417e-38, 4.028054e-38, 
    4.092578e-38, 4.049066e-38, 4.126516e-38, 4.082153e-38, 4.089048e-38, 
    4.047635e-38, 3.814463e-38, 3.856556e-38, 3.811979e-38, 3.817949e-38, 
    3.815274e-38, 3.782906e-38, 3.766751e-38, 3.733258e-38, 3.739315e-38, 
    3.763934e-38, 3.820637e-38, 3.801226e-38, 3.850388e-38, 3.849271e-38, 
    3.905051e-38, 3.879645e-38, 3.975607e-38, 3.94805e-38, 4.028653e-38, 
    4.008041e-38, 4.027678e-38, 4.021715e-38, 4.027756e-38, 3.997596e-38, 
    4.010474e-38, 3.984232e-38, 3.884349e-38, 3.913374e-38, 3.828215e-38, 
    3.77829e-38, 3.745714e-38, 3.722794e-38, 3.726025e-38, 3.732189e-38, 
    3.764079e-38, 3.794382e-38, 3.817781e-38, 3.833527e-38, 3.84911e-38, 
    3.896793e-38, 3.922657e-38, 3.981193e-38, 3.970581e-38, 3.988593e-38, 
    4.005998e-38, 4.035618e-38, 4.030729e-38, 4.043833e-38, 3.98813e-38, 
    4.025e-38, 3.964544e-38, 3.980888e-38, 3.853282e-38, 3.806456e-38, 
    3.786741e-38, 3.769682e-38, 3.72851e-38, 3.756871e-38, 3.74566e-38, 
    3.772432e-38, 3.789547e-38, 3.781075e-38, 3.833958e-38, 3.813261e-38, 
    3.924196e-38, 3.875662e-38, 4.003947e-38, 3.972758e-38, 4.011549e-38, 
    3.99163e-38, 4.025893e-38, 3.995008e-38, 4.048729e-38, 4.060535e-38, 
    4.052461e-38, 4.083599e-38, 3.99332e-38, 4.027671e-38, 3.780834e-38, 
    3.782214e-38, 3.788658e-38, 3.760415e-38, 3.758699e-38, 3.733088e-38, 
    3.755869e-38, 3.765628e-38, 3.790547e-38, 3.80541e-38, 3.819644e-38, 
    3.851136e-38, 3.886653e-38, 3.937653e-38, 3.974767e-38, 3.999858e-38, 
    3.984455e-38, 3.998043e-38, 3.982853e-38, 3.975758e-38, 4.056102e-38, 
    4.01059e-38, 4.079104e-38, 4.075282e-38, 4.044143e-38, 4.075712e-38, 
    3.783185e-38, 3.775247e-38, 3.747812e-38, 3.769262e-38, 3.730312e-38, 
    3.752035e-38, 3.764602e-38, 3.813676e-38, 3.824615e-38, 3.834765e-38, 
    3.854908e-38, 3.880931e-38, 3.927639e-38, 3.96887e-38, 4.007024e-38, 
    4.004187e-38, 4.005185e-38, 4.013841e-38, 3.992516e-38, 4.017369e-38, 
    4.021564e-38, 4.010594e-38, 4.07477e-38, 4.056321e-38, 4.0752e-38, 
    4.063179e-38, 3.777827e-38, 3.791206e-38, 3.783969e-38, 3.797588e-38, 
    3.787982e-38, 3.831093e-38, 3.844137e-38, 3.906132e-38, 3.880411e-38, 
    3.921518e-38, 3.884532e-38, 3.891004e-38, 3.922838e-38, 3.886505e-38, 
    3.96657e-38, 3.912046e-38, 4.014178e-38, 3.95881e-38, 4.017707e-38, 
    4.006857e-38, 4.024846e-38, 4.041025e-38, 4.061495e-38, 4.099545e-38, 
    4.090702e-38, 4.122763e-38, 3.811347e-38, 3.828985e-38, 3.827443e-38, 
    3.845994e-38, 3.85977e-38, 3.889881e-38, 3.939383e-38, 3.920695e-38, 
    3.955092e-38, 3.96203e-38, 3.90981e-38, 3.941772e-38, 3.840847e-38, 
    3.856812e-38, 3.847309e-38, 3.812727e-38, 3.924974e-38, 3.866636e-38, 
    3.975381e-38, 3.943058e-38, 4.038712e-38, 3.990561e-38, 4.08584e-38, 
    4.127349e-38, 4.166918e-38, 4.213624e-38, 3.838662e-38, 3.826636e-38, 
    3.84821e-38, 3.87825e-38, 3.906695e-38, 3.945019e-38, 3.94897e-38, 
    3.956197e-38, 3.975001e-38, 3.990878e-38, 3.958471e-38, 3.99487e-38, 
    3.860495e-38, 3.930116e-38, 3.822086e-38, 3.854058e-38, 3.876473e-38, 
    3.866637e-38, 3.918569e-38, 3.930987e-38, 3.981877e-38, 3.955491e-38, 
    4.117047e-38, 4.044431e-38, 4.249641e-38, 4.191119e-38, 3.822439e-38, 
    3.838627e-38, 3.895655e-38, 3.868336e-38, 3.947599e-38, 3.967439e-38, 
    3.983659e-38, 4.004542e-38, 4.006836e-38, 4.019398e-38, 3.99884e-38, 
    4.018589e-38, 3.945101e-38, 3.977652e-38, 3.889025e-38, 3.91039e-38, 
    3.900548e-38, 3.889772e-38, 3.923129e-38, 3.958976e-38, 3.959769e-38, 
    3.971335e-38, 4.004146e-38, 3.947925e-38, 4.126481e-38, 4.014726e-38, 
    3.856359e-38, 3.887905e-38, 3.892509e-38, 3.880171e-38, 3.965445e-38, 
    3.934274e-38, 4.019095e-38, 3.995796e-38, 4.034084e-38, 4.014983e-38, 
    4.01218e-38, 3.987965e-38, 3.973067e-38, 3.935694e-38, 3.905567e-38, 
    3.881955e-38, 3.887388e-38, 3.913449e-38, 3.961185e-38, 4.007034e-38, 
    3.996859e-38, 4.031157e-38, 3.941772e-38, 3.978806e-38, 3.964441e-38, 
    4.002055e-38, 3.920195e-38, 3.989687e-38, 3.902631e-38, 3.910187e-38, 
    3.933659e-38, 3.981316e-38, 3.991977e-38, 4.003407e-38, 3.996334e-38, 
    3.962409e-38, 3.956891e-38, 3.933092e-38, 3.926536e-38, 3.908543e-38, 
    3.893701e-38, 3.907253e-38, 3.921535e-38, 3.962433e-38, 3.999672e-38, 
    4.041253e-38, 4.05151e-38, 4.100775e-38, 4.060588e-38, 4.127108e-38, 
    4.070428e-38, 4.169129e-38, 3.993789e-38, 4.068823e-38, 3.934738e-38, 
    3.948862e-38, 3.974521e-38, 4.034565e-38, 4.001875e-38, 4.040146e-38, 
    3.956677e-38, 3.914341e-38, 3.903494e-38, 3.88337e-38, 3.903957e-38, 
    3.902273e-38, 3.922144e-38, 3.915748e-38, 3.963799e-38, 3.937912e-38, 
    4.012103e-38, 4.039848e-38, 4.119381e-38, 4.168986e-38, 4.220219e-38, 
    4.243053e-38, 4.250034e-38, 4.252955e-38,
  2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.522337e-44, 2.382207e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.662467e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 2.662467e-44, 
    2.522337e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.522337e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.382207e-44, 2.522337e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.522337e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.522337e-44, 2.382207e-44, 
    2.522337e-44, 2.382207e-44, 2.382207e-44, 2.522337e-44, 2.382207e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.522337e-44, 2.382207e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.382207e-44, 2.522337e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 
    2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.662467e-44, 2.522337e-44, 2.662467e-44, 2.662467e-44, 2.382207e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.382207e-44, 2.522337e-44, 
    2.522337e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 
    2.382207e-44, 2.382207e-44, 2.382207e-44, 2.382207e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.382207e-44, 2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.382207e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.662467e-44, 2.522337e-44, 2.662467e-44, 
    2.522337e-44, 2.662467e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.382207e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 2.522337e-44, 
    2.522337e-44, 2.522337e-44, 2.662467e-44, 2.662467e-44, 2.662467e-44, 
    2.662467e-44, 2.662467e-44, 2.662467e-44,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_CH4_UNSAT =
  2.094769e-05, 2.075876e-05, 2.079554e-05, 2.06428e-05, 2.072758e-05, 
    2.062749e-05, 2.090945e-05, 2.075124e-05, 2.085229e-05, 2.093072e-05, 
    2.034526e-05, 2.063597e-05, 2.004191e-05, 2.022837e-05, 1.975897e-05, 
    2.007095e-05, 1.969588e-05, 1.976801e-05, 1.955073e-05, 1.961305e-05, 
    1.933432e-05, 1.952195e-05, 1.918941e-05, 1.937919e-05, 1.934953e-05, 
    1.952812e-05, 2.05776e-05, 2.038152e-05, 2.058919e-05, 2.056128e-05, 
    2.057381e-05, 2.072582e-05, 2.080227e-05, 2.096212e-05, 2.093314e-05, 
    2.081572e-05, 2.054872e-05, 2.06395e-05, 2.041049e-05, 2.041567e-05, 
    2.015973e-05, 2.027526e-05, 1.984352e-05, 1.996653e-05, 1.961045e-05, 
    1.970018e-05, 1.961467e-05, 1.964061e-05, 1.961433e-05, 1.974588e-05, 
    1.968955e-05, 1.980519e-05, 2.025363e-05, 2.012216e-05, 2.051345e-05, 
    2.07475e-05, 2.090251e-05, 2.101225e-05, 2.099675e-05, 2.096718e-05, 
    2.081504e-05, 2.067165e-05, 2.056215e-05, 2.048878e-05, 2.041642e-05, 
    2.01968e-05, 2.008029e-05, 1.981861e-05, 1.986593e-05, 1.978576e-05, 
    1.97091e-05, 1.958017e-05, 1.960142e-05, 1.954455e-05, 1.978789e-05, 
    1.962626e-05, 1.989287e-05, 1.982005e-05, 2.039666e-05, 2.061503e-05, 
    2.070755e-05, 2.078847e-05, 2.098483e-05, 2.084929e-05, 2.090275e-05, 
    2.077549e-05, 2.069448e-05, 2.073456e-05, 2.048678e-05, 2.058323e-05, 
    2.007338e-05, 2.02935e-05, 1.971805e-05, 1.985622e-05, 1.968489e-05, 
    1.977238e-05, 1.962239e-05, 1.975739e-05, 1.952338e-05, 1.94723e-05, 
    1.950721e-05, 1.937305e-05, 1.976487e-05, 1.961466e-05, 2.073568e-05, 
    2.072915e-05, 2.06987e-05, 2.083244e-05, 2.084061e-05, 2.096291e-05, 
    2.085411e-05, 2.080771e-05, 2.068979e-05, 2.061991e-05, 2.055342e-05, 
    2.040698e-05, 2.024301e-05, 2.001301e-05, 1.984728e-05, 1.973594e-05, 
    1.980423e-05, 1.974394e-05, 1.981134e-05, 1.98429e-05, 1.949144e-05, 
    1.968902e-05, 1.939236e-05, 1.940881e-05, 1.954319e-05, 1.940696e-05, 
    2.072456e-05, 2.076216e-05, 2.089251e-05, 2.079053e-05, 2.097622e-05, 
    2.087234e-05, 2.081252e-05, 2.05812e-05, 2.053027e-05, 2.048299e-05, 
    2.038952e-05, 2.026935e-05, 2.005797e-05, 1.98735e-05, 1.970464e-05, 
    1.971703e-05, 1.971267e-05, 1.967489e-05, 1.976843e-05, 1.965952e-05, 
    1.964121e-05, 1.968905e-05, 1.941102e-05, 1.949057e-05, 1.940916e-05, 
    1.946097e-05, 2.074994e-05, 2.068665e-05, 2.072086e-05, 2.065651e-05, 
    2.070185e-05, 2.049998e-05, 2.043933e-05, 2.015475e-05, 2.027171e-05, 
    2.008548e-05, 2.025282e-05, 2.02232e-05, 2.007936e-05, 2.02438e-05, 
    1.988367e-05, 2.012802e-05, 1.967342e-05, 1.99182e-05, 1.965805e-05, 
    1.970537e-05, 1.9627e-05, 1.955672e-05, 1.946822e-05, 1.930459e-05, 
    1.934251e-05, 1.920545e-05, 2.059217e-05, 2.050985e-05, 2.051711e-05, 
    2.043085e-05, 2.036698e-05, 2.022833e-05, 2.00053e-05, 2.008927e-05, 
    1.993505e-05, 1.990404e-05, 2.013831e-05, 1.999456e-05, 2.045469e-05, 
    2.038057e-05, 2.042472e-05, 2.058568e-05, 2.006991e-05, 2.033513e-05, 
    1.984453e-05, 1.998886e-05, 1.956675e-05, 1.9777e-05, 1.936338e-05, 
    1.918575e-05, 1.901821e-05, 1.882184e-05, 2.046488e-05, 2.052087e-05, 
    2.042059e-05, 2.028156e-05, 2.015231e-05, 1.998006e-05, 1.996242e-05, 
    1.993008e-05, 1.984627e-05, 1.977571e-05, 1.991984e-05, 1.975801e-05, 
    2.036334e-05, 2.004684e-05, 2.054202e-05, 2.039331e-05, 2.028977e-05, 
    2.033522e-05, 2.009886e-05, 2.004302e-05, 1.98156e-05, 1.993327e-05, 
    1.922962e-05, 1.954185e-05, 1.8672e-05, 1.891617e-05, 2.054042e-05, 
    2.046508e-05, 2.020213e-05, 2.032738e-05, 1.996855e-05, 1.987991e-05, 
    1.980777e-05, 1.971542e-05, 1.970545e-05, 1.965066e-05, 1.974042e-05, 
    1.965422e-05, 1.997969e-05, 1.983445e-05, 2.023226e-05, 2.013565e-05, 
    2.018012e-05, 2.022884e-05, 2.007834e-05, 1.991757e-05, 1.991415e-05, 
    1.986251e-05, 1.971674e-05, 1.996709e-05, 1.918918e-05, 1.967064e-05, 
    2.038282e-05, 2.023722e-05, 2.021642e-05, 2.027287e-05, 1.98888e-05, 
    2.002823e-05, 1.9652e-05, 1.97539e-05, 1.958686e-05, 1.966992e-05, 
    1.968213e-05, 1.978863e-05, 1.985485e-05, 2.002184e-05, 2.015739e-05, 
    2.026469e-05, 2.023976e-05, 2.012184e-05, 1.990773e-05, 1.970454e-05, 
    1.97491e-05, 1.959957e-05, 1.999464e-05, 1.982926e-05, 1.989322e-05, 
    1.972632e-05, 2.009149e-05, 1.978059e-05, 2.017071e-05, 2.013661e-05, 
    2.0031e-05, 1.981801e-05, 1.977083e-05, 1.972038e-05, 1.975152e-05, 
    1.990229e-05, 1.992697e-05, 2.003357e-05, 2.006296e-05, 2.014404e-05, 
    2.021107e-05, 2.014982e-05, 2.008543e-05, 1.990223e-05, 1.973668e-05, 
    1.955572e-05, 1.951137e-05, 1.929911e-05, 1.947192e-05, 1.918649e-05, 
    1.942919e-05, 1.900853e-05, 1.976256e-05, 1.943636e-05, 2.002619e-05, 
    1.996291e-05, 1.984827e-05, 1.958461e-05, 1.97271e-05, 1.956044e-05, 
    1.992793e-05, 2.011776e-05, 2.016681e-05, 2.025817e-05, 2.016471e-05, 
    2.017232e-05, 2.008278e-05, 2.011157e-05, 1.989614e-05, 2.001195e-05, 
    1.968243e-05, 1.956176e-05, 1.921982e-05, 1.900934e-05, 1.879447e-05, 
    1.869939e-05, 1.867042e-05, 1.865831e-05,
  1.394619e-05, 1.376974e-05, 1.380408e-05, 1.366155e-05, 1.374065e-05, 
    1.364727e-05, 1.391046e-05, 1.376272e-05, 1.385707e-05, 1.393034e-05, 
    1.33843e-05, 1.365519e-05, 1.310226e-05, 1.327557e-05, 1.283974e-05, 
    1.312923e-05, 1.278128e-05, 1.284813e-05, 1.26469e-05, 1.270458e-05, 
    1.244679e-05, 1.262027e-05, 1.231302e-05, 1.248826e-05, 1.246085e-05, 
    1.262598e-05, 1.360076e-05, 1.341805e-05, 1.361157e-05, 1.358554e-05, 
    1.359722e-05, 1.373901e-05, 1.381036e-05, 1.395969e-05, 1.39326e-05, 
    1.382292e-05, 1.357383e-05, 1.365848e-05, 1.344506e-05, 1.344989e-05, 
    1.321174e-05, 1.331918e-05, 1.291814e-05, 1.303228e-05, 1.270218e-05, 
    1.278527e-05, 1.270608e-05, 1.27301e-05, 1.270576e-05, 1.282762e-05, 
    1.277542e-05, 1.28826e-05, 1.329907e-05, 1.317682e-05, 1.354096e-05, 
    1.375922e-05, 1.390398e-05, 1.400654e-05, 1.399205e-05, 1.396441e-05, 
    1.382228e-05, 1.368847e-05, 1.358636e-05, 1.351799e-05, 1.345058e-05, 
    1.324619e-05, 1.313791e-05, 1.289503e-05, 1.293893e-05, 1.286458e-05, 
    1.279354e-05, 1.267415e-05, 1.269381e-05, 1.264117e-05, 1.286656e-05, 
    1.27168e-05, 1.296392e-05, 1.289638e-05, 1.343215e-05, 1.363565e-05, 
    1.372194e-05, 1.379747e-05, 1.39809e-05, 1.385427e-05, 1.390421e-05, 
    1.378537e-05, 1.370976e-05, 1.374717e-05, 1.351612e-05, 1.360601e-05, 
    1.313149e-05, 1.333615e-05, 1.280183e-05, 1.292992e-05, 1.277111e-05, 
    1.285218e-05, 1.271323e-05, 1.283829e-05, 1.262159e-05, 1.257434e-05, 
    1.260663e-05, 1.248259e-05, 1.284522e-05, 1.270607e-05, 1.374821e-05, 
    1.374211e-05, 1.37137e-05, 1.383853e-05, 1.384616e-05, 1.396042e-05, 
    1.385877e-05, 1.381544e-05, 1.370539e-05, 1.364021e-05, 1.357822e-05, 
    1.344179e-05, 1.328918e-05, 1.307543e-05, 1.292162e-05, 1.281841e-05, 
    1.288171e-05, 1.282582e-05, 1.28883e-05, 1.291757e-05, 1.259204e-05, 
    1.277493e-05, 1.250044e-05, 1.251565e-05, 1.263992e-05, 1.251393e-05, 
    1.373783e-05, 1.377293e-05, 1.389464e-05, 1.37994e-05, 1.397286e-05, 
    1.38758e-05, 1.381993e-05, 1.360411e-05, 1.355665e-05, 1.351259e-05, 
    1.342553e-05, 1.331369e-05, 1.311719e-05, 1.294594e-05, 1.278941e-05, 
    1.280089e-05, 1.279685e-05, 1.276184e-05, 1.284852e-05, 1.274761e-05, 
    1.273065e-05, 1.277496e-05, 1.251768e-05, 1.259124e-05, 1.251597e-05, 
    1.256387e-05, 1.376152e-05, 1.370246e-05, 1.373438e-05, 1.367434e-05, 
    1.371663e-05, 1.352841e-05, 1.34719e-05, 1.32071e-05, 1.331588e-05, 
    1.314273e-05, 1.329832e-05, 1.327076e-05, 1.313704e-05, 1.328992e-05, 
    1.295537e-05, 1.318226e-05, 1.276048e-05, 1.29874e-05, 1.274624e-05, 
    1.279009e-05, 1.27175e-05, 1.265244e-05, 1.257057e-05, 1.241934e-05, 
    1.245438e-05, 1.232783e-05, 1.361435e-05, 1.35376e-05, 1.354438e-05, 
    1.346402e-05, 1.340455e-05, 1.327554e-05, 1.306827e-05, 1.314627e-05, 
    1.300306e-05, 1.297428e-05, 1.319184e-05, 1.30583e-05, 1.348622e-05, 
    1.341719e-05, 1.345831e-05, 1.360829e-05, 1.312827e-05, 1.337489e-05, 
    1.291907e-05, 1.3053e-05, 1.266172e-05, 1.285645e-05, 1.247366e-05, 
    1.230963e-05, 1.215518e-05, 1.19744e-05, 1.349571e-05, 1.354789e-05, 
    1.345447e-05, 1.332504e-05, 1.320485e-05, 1.304484e-05, 1.302846e-05, 
    1.299845e-05, 1.292069e-05, 1.285526e-05, 1.298894e-05, 1.283886e-05, 
    1.340113e-05, 1.310685e-05, 1.356759e-05, 1.342904e-05, 1.333268e-05, 
    1.337498e-05, 1.315518e-05, 1.31033e-05, 1.289224e-05, 1.300141e-05, 
    1.235012e-05, 1.263867e-05, 1.183668e-05, 1.20612e-05, 1.35661e-05, 
    1.34959e-05, 1.325116e-05, 1.336769e-05, 1.303416e-05, 1.295189e-05, 
    1.288499e-05, 1.279939e-05, 1.279016e-05, 1.273941e-05, 1.282255e-05, 
    1.27427e-05, 1.30445e-05, 1.290973e-05, 1.327919e-05, 1.318937e-05, 
    1.323071e-05, 1.327601e-05, 1.313611e-05, 1.298683e-05, 1.298367e-05, 
    1.293575e-05, 1.280057e-05, 1.30328e-05, 1.231278e-05, 1.275788e-05, 
    1.341929e-05, 1.328379e-05, 1.326445e-05, 1.331697e-05, 1.296014e-05, 
    1.308956e-05, 1.274065e-05, 1.283505e-05, 1.268034e-05, 1.275724e-05, 
    1.276855e-05, 1.286725e-05, 1.292865e-05, 1.308363e-05, 1.320958e-05, 
    1.330936e-05, 1.328617e-05, 1.317653e-05, 1.29777e-05, 1.278931e-05, 
    1.28306e-05, 1.26921e-05, 1.305837e-05, 1.290491e-05, 1.296424e-05, 
    1.280949e-05, 1.314833e-05, 1.285976e-05, 1.322196e-05, 1.319026e-05, 
    1.309213e-05, 1.289448e-05, 1.285074e-05, 1.280398e-05, 1.283284e-05, 
    1.297265e-05, 1.299556e-05, 1.309452e-05, 1.312182e-05, 1.319716e-05, 
    1.325949e-05, 1.320254e-05, 1.314269e-05, 1.297261e-05, 1.281909e-05, 
    1.265151e-05, 1.261048e-05, 1.241427e-05, 1.257397e-05, 1.231029e-05, 
    1.253444e-05, 1.214624e-05, 1.284306e-05, 1.254109e-05, 1.308767e-05, 
    1.302892e-05, 1.292253e-05, 1.267824e-05, 1.281022e-05, 1.265587e-05, 
    1.299645e-05, 1.317273e-05, 1.321833e-05, 1.330329e-05, 1.321639e-05, 
    1.322346e-05, 1.314024e-05, 1.316699e-05, 1.296696e-05, 1.307445e-05, 
    1.276883e-05, 1.26571e-05, 1.234109e-05, 1.2147e-05, 1.194924e-05, 
    1.186185e-05, 1.183524e-05, 1.182412e-05,
  5.604382e-06, 5.5068e-06, 5.525749e-06, 5.44722e-06, 5.490761e-06, 
    5.439374e-06, 5.584579e-06, 5.502927e-06, 5.55503e-06, 5.595593e-06, 
    5.295431e-06, 5.443723e-06, 5.142336e-06, 5.236251e-06, 5.001041e-06, 
    5.156919e-06, 4.96974e-06, 5.005538e-06, 4.898003e-06, 4.928757e-06, 
    4.791762e-06, 4.883823e-06, 4.721124e-06, 4.813719e-06, 4.7992e-06, 
    4.886865e-06, 5.41383e-06, 5.313844e-06, 5.419762e-06, 5.405479e-06, 
    5.41189e-06, 5.489856e-06, 5.529216e-06, 5.611863e-06, 5.596845e-06, 
    5.536156e-06, 5.39906e-06, 5.445534e-06, 5.328587e-06, 5.331222e-06, 
    5.201604e-06, 5.259966e-06, 5.043116e-06, 5.104555e-06, 4.927473e-06, 
    4.971875e-06, 4.929554e-06, 4.94238e-06, 4.929387e-06, 4.994545e-06, 
    4.966604e-06, 5.024029e-06, 5.249023e-06, 5.182679e-06, 5.381044e-06, 
    5.501001e-06, 5.580991e-06, 5.63787e-06, 5.629823e-06, 5.614484e-06, 
    5.535801e-06, 5.462026e-06, 5.405928e-06, 5.368463e-06, 5.331601e-06, 
    5.220297e-06, 5.161614e-06, 5.030705e-06, 5.054289e-06, 5.01436e-06, 
    4.976298e-06, 4.912523e-06, 4.923009e-06, 4.894954e-06, 5.015422e-06, 
    4.935281e-06, 5.06773e-06, 5.031426e-06, 5.321538e-06, 5.432991e-06, 
    5.480455e-06, 5.522103e-06, 5.623635e-06, 5.55348e-06, 5.581116e-06, 
    5.515422e-06, 5.473749e-06, 5.494354e-06, 5.367439e-06, 5.41671e-06, 
    5.15814e-06, 5.269201e-06, 4.980735e-06, 5.049448e-06, 4.964297e-06, 
    5.00771e-06, 4.933372e-06, 5.000265e-06, 4.884526e-06, 4.859399e-06, 
    4.876566e-06, 4.810716e-06, 5.003978e-06, 4.92955e-06, 5.49493e-06, 
    5.491568e-06, 5.475916e-06, 5.54478e-06, 5.549e-06, 5.612273e-06, 
    5.555971e-06, 5.532024e-06, 5.471339e-06, 5.435495e-06, 5.401467e-06, 
    5.326799e-06, 5.243646e-06, 5.127839e-06, 5.044987e-06, 4.989612e-06, 
    5.023554e-06, 4.993584e-06, 5.027088e-06, 5.04281e-06, 4.868808e-06, 
    4.96634e-06, 4.820175e-06, 4.828239e-06, 4.894285e-06, 4.82733e-06, 
    5.489208e-06, 5.508557e-06, 5.575819e-06, 5.523168e-06, 5.619172e-06, 
    5.565389e-06, 5.534504e-06, 5.415669e-06, 5.389638e-06, 5.365508e-06, 
    5.317924e-06, 5.256975e-06, 5.150403e-06, 5.058061e-06, 4.974088e-06, 
    4.980231e-06, 4.978067e-06, 4.959342e-06, 5.005747e-06, 4.951734e-06, 
    4.942677e-06, 4.966358e-06, 4.829319e-06, 4.868381e-06, 4.82841e-06, 
    4.853836e-06, 5.502267e-06, 5.469727e-06, 5.487305e-06, 5.454256e-06, 
    5.477531e-06, 5.374169e-06, 5.343254e-06, 5.19909e-06, 5.258171e-06, 
    5.164222e-06, 5.248615e-06, 5.233638e-06, 5.161142e-06, 5.244051e-06, 
    5.063133e-06, 5.185625e-06, 4.958615e-06, 5.080371e-06, 4.951006e-06, 
    4.97445e-06, 4.935652e-06, 4.900956e-06, 4.857395e-06, 4.77724e-06, 
    4.795775e-06, 4.728929e-06, 5.421289e-06, 5.379205e-06, 5.382917e-06, 
    5.338947e-06, 5.306472e-06, 5.236234e-06, 5.123976e-06, 5.166133e-06, 
    5.088806e-06, 5.073309e-06, 5.190815e-06, 5.118591e-06, 5.351084e-06, 
    5.313369e-06, 5.335825e-06, 5.417961e-06, 5.156399e-06, 5.290301e-06, 
    5.043618e-06, 5.115734e-06, 4.905899e-06, 5.010003e-06, 4.805984e-06, 
    4.719342e-06, 4.638185e-06, 4.543729e-06, 5.356275e-06, 5.384838e-06, 
    5.333725e-06, 5.263151e-06, 5.197869e-06, 5.111327e-06, 5.102496e-06, 
    5.08632e-06, 5.044486e-06, 5.009365e-06, 5.0812e-06, 5.000571e-06, 
    5.304611e-06, 5.144814e-06, 5.395636e-06, 5.319841e-06, 5.26731e-06, 
    5.290351e-06, 5.170958e-06, 5.142898e-06, 5.029205e-06, 5.087915e-06, 
    4.740683e-06, 4.893622e-06, 4.472164e-06, 4.58901e-06, 5.394822e-06, 
    5.356378e-06, 5.222995e-06, 5.286375e-06, 5.105566e-06, 5.061261e-06, 
    5.025313e-06, 4.979428e-06, 4.974487e-06, 4.947351e-06, 4.991834e-06, 
    4.94911e-06, 5.111144e-06, 5.038595e-06, 5.238218e-06, 5.189475e-06, 
    5.21189e-06, 5.236493e-06, 5.160638e-06, 5.080065e-06, 5.078361e-06, 
    5.052582e-06, 4.980066e-06, 5.104837e-06, 4.720999e-06, 4.957226e-06, 
    5.314518e-06, 5.240718e-06, 5.230213e-06, 5.258761e-06, 5.065699e-06, 
    5.135474e-06, 4.948015e-06, 4.998531e-06, 4.915825e-06, 4.956883e-06, 
    4.96293e-06, 5.015792e-06, 5.048762e-06, 5.132267e-06, 5.200429e-06, 
    5.25462e-06, 5.242011e-06, 5.182519e-06, 5.075148e-06, 4.974032e-06, 
    4.996142e-06, 4.9221e-06, 5.118632e-06, 5.036009e-06, 5.067904e-06, 
    4.984836e-06, 5.16725e-06, 5.011778e-06, 5.207146e-06, 5.189957e-06, 
    5.136862e-06, 5.030406e-06, 5.006942e-06, 4.981887e-06, 4.997347e-06, 
    5.072432e-06, 5.084763e-06, 5.138154e-06, 5.152909e-06, 5.1937e-06, 
    5.227514e-06, 5.196614e-06, 5.164201e-06, 5.072406e-06, 4.98998e-06, 
    4.900461e-06, 4.878615e-06, 4.774558e-06, 4.859205e-06, 4.719687e-06, 
    4.838212e-06, 4.633499e-06, 5.002822e-06, 4.841738e-06, 5.134453e-06, 
    5.102742e-06, 5.045477e-06, 4.914705e-06, 4.985226e-06, 4.902782e-06, 
    5.085247e-06, 5.180461e-06, 5.205176e-06, 5.25132e-06, 5.204122e-06, 
    5.207958e-06, 5.16287e-06, 5.177351e-06, 5.069365e-06, 5.12731e-06, 
    4.963078e-06, 4.903436e-06, 4.735919e-06, 4.633899e-06, 4.53063e-06, 
    4.485216e-06, 4.471417e-06, 4.465651e-06,
  1.104549e-06, 1.075706e-06, 1.081285e-06, 1.058232e-06, 1.070992e-06, 
    1.055939e-06, 1.098673e-06, 1.074567e-06, 1.089927e-06, 1.10194e-06, 
    1.014189e-06, 1.05721e-06, 9.704585e-07, 9.97201e-07, 9.307226e-07, 
    9.745937e-07, 9.220014e-07, 9.319777e-07, 9.021263e-07, 9.106276e-07, 
    8.729814e-07, 8.982164e-07, 8.537949e-07, 8.789762e-07, 8.750106e-07, 
    8.990546e-07, 1.048485e-06, 1.019496e-06, 1.050214e-06, 1.046053e-06, 
    1.04792e-06, 1.070726e-06, 1.082307e-06, 1.106772e-06, 1.102311e-06, 
    1.084354e-06, 1.044184e-06, 1.057739e-06, 1.02375e-06, 1.024512e-06, 
    9.873045e-07, 1.003996e-06, 9.424919e-07, 9.597741e-07, 9.102721e-07, 
    9.225952e-07, 9.108484e-07, 9.144027e-07, 9.108022e-07, 9.289099e-07, 
    9.211292e-07, 9.37146e-07, 1.000858e-06, 9.819137e-07, 1.038946e-06, 
    1.074001e-06, 1.09761e-06, 1.114511e-06, 1.112114e-06, 1.107551e-06, 
    1.084249e-06, 1.062565e-06, 1.046183e-06, 1.035294e-06, 1.024621e-06, 
    9.926401e-07, 9.759264e-07, 9.390149e-07, 9.456261e-07, 9.344424e-07, 
    9.23826e-07, 9.061366e-07, 9.090366e-07, 9.012853e-07, 9.34739e-07, 
    9.12435e-07, 9.494018e-07, 9.392164e-07, 1.021716e-06, 1.054074e-06, 
    1.067967e-06, 1.080211e-06, 1.110273e-06, 1.089469e-06, 1.097647e-06, 
    1.078243e-06, 1.066e-06, 1.072047e-06, 1.034998e-06, 1.049325e-06, 
    9.749402e-07, 1.006646e-06, 9.25061e-07, 9.442675e-07, 9.204878e-07, 
    9.325841e-07, 9.119059e-07, 9.305055e-07, 8.984101e-07, 8.914964e-07, 
    8.962177e-07, 8.781554e-07, 9.315419e-07, 9.108472e-07, 1.072216e-06, 
    1.071229e-06, 1.066635e-06, 1.086899e-06, 1.088145e-06, 1.106893e-06, 
    1.090205e-06, 1.083135e-06, 1.065293e-06, 1.054806e-06, 1.044885e-06, 
    1.023234e-06, 9.993182e-07, 9.663535e-07, 9.430163e-07, 9.275342e-07, 
    9.370131e-07, 9.286419e-07, 9.380018e-07, 9.424058e-07, 8.940829e-07, 
    9.21056e-07, 8.807417e-07, 8.829487e-07, 9.011008e-07, 8.826999e-07, 
    1.070536e-06, 1.076223e-06, 1.096078e-06, 1.080524e-06, 1.108945e-06, 
    1.09299e-06, 1.083867e-06, 1.049021e-06, 1.041444e-06, 1.034437e-06, 
    1.020672e-06, 1.003138e-06, 9.727451e-07, 9.466854e-07, 9.232107e-07, 
    9.249208e-07, 9.243184e-07, 9.191108e-07, 9.32036e-07, 9.169979e-07, 
    9.14485e-07, 9.210607e-07, 8.832444e-07, 8.939654e-07, 8.829956e-07, 
    8.899679e-07, 1.074373e-06, 1.064821e-06, 1.069977e-06, 1.06029e-06, 
    1.067109e-06, 1.03695e-06, 1.027992e-06, 9.865879e-07, 1.003481e-06, 
    9.766668e-07, 1.000741e-06, 9.964534e-07, 9.757928e-07, 9.994337e-07, 
    9.481104e-07, 9.827528e-07, 9.189088e-07, 9.529585e-07, 9.167957e-07, 
    9.233116e-07, 9.125375e-07, 9.029416e-07, 8.909456e-07, 8.690241e-07, 
    8.740758e-07, 8.559072e-07, 1.05066e-06, 1.038413e-06, 1.03949e-06, 
    1.026745e-06, 1.017369e-06, 9.971959e-07, 9.652606e-07, 9.772092e-07, 
    9.55333e-07, 9.509706e-07, 9.842296e-07, 9.637384e-07, 1.030258e-06, 
    1.019358e-06, 1.025843e-06, 1.049689e-06, 9.744459e-07, 1.012712e-06, 
    9.426326e-07, 9.629309e-07, 9.043063e-07, 9.332249e-07, 8.768625e-07, 
    8.533131e-07, 8.314643e-07, 8.062941e-07, 1.031761e-06, 1.040048e-06, 
    1.025235e-06, 1.00491e-06, 9.862395e-07, 9.616862e-07, 9.591929e-07, 
    9.54633e-07, 9.428758e-07, 9.330464e-07, 9.531912e-07, 9.305908e-07, 
    1.016833e-06, 9.711604e-07, 1.043188e-06, 1.021226e-06, 1.006103e-06, 
    1.012726e-06, 9.785801e-07, 9.706171e-07, 9.385946e-07, 9.55082e-07, 
    8.590924e-07, 9.00918e-07, 7.874093e-07, 8.183256e-07, 1.042951e-06, 
    1.031791e-06, 9.934104e-07, 1.011582e-06, 9.600594e-07, 9.47584e-07, 
    9.375053e-07, 9.246975e-07, 9.233219e-07, 9.157817e-07, 9.281538e-07, 
    9.162697e-07, 9.616342e-07, 9.412246e-07, 9.977637e-07, 9.838483e-07, 
    9.902386e-07, 9.9727e-07, 9.756486e-07, 9.528717e-07, 9.52392e-07, 
    9.451472e-07, 9.248761e-07, 9.598535e-07, 8.537621e-07, 9.185242e-07, 
    1.019689e-06, 9.9848e-07, 9.954737e-07, 1.00365e-06, 9.488309e-07, 
    9.685143e-07, 9.159656e-07, 9.300217e-07, 9.070492e-07, 9.184277e-07, 
    9.201077e-07, 9.348424e-07, 9.440752e-07, 9.676066e-07, 9.869694e-07, 
    1.002462e-06, 9.988495e-07, 9.818682e-07, 9.514882e-07, 9.231956e-07, 
    9.293556e-07, 9.087849e-07, 9.637496e-07, 9.405002e-07, 9.494509e-07, 
    9.262035e-07, 9.775268e-07, 9.337217e-07, 9.888848e-07, 9.839854e-07, 
    9.689072e-07, 9.389311e-07, 9.323695e-07, 9.253822e-07, 9.296914e-07, 
    9.50724e-07, 9.541943e-07, 9.692732e-07, 9.734556e-07, 9.850513e-07, 
    9.947017e-07, 9.858817e-07, 9.766605e-07, 9.507167e-07, 9.276371e-07, 
    9.028048e-07, 8.967817e-07, 8.682948e-07, 8.914433e-07, 8.534075e-07, 
    8.856826e-07, 8.302098e-07, 9.312201e-07, 8.866489e-07, 9.682252e-07, 
    9.592625e-07, 9.431541e-07, 9.067402e-07, 9.263122e-07, 9.034459e-07, 
    9.543307e-07, 9.812829e-07, 9.883228e-07, 1.001516e-06, 9.880222e-07, 
    9.891164e-07, 9.762824e-07, 9.803977e-07, 9.498614e-07, 9.662037e-07, 
    9.201489e-07, 9.036263e-07, 8.578007e-07, 8.303164e-07, 8.028252e-07, 
    7.908413e-07, 7.87213e-07, 7.856985e-07,
  8.152712e-08, 7.847502e-08, 7.906245e-08, 7.664418e-08, 7.797968e-08, 
    7.640492e-08, 8.090232e-08, 7.835528e-08, 7.997516e-08, 8.124945e-08, 
    7.209113e-08, 7.653749e-08, 6.765902e-08, 7.035874e-08, 6.371003e-08, 
    6.807431e-08, 6.285342e-08, 6.383357e-08, 6.091499e-08, 6.174177e-08, 
    5.810753e-08, 6.053593e-08, 5.628225e-08, 5.868156e-08, 5.830163e-08, 
    6.061714e-08, 7.562888e-08, 7.2635e-08, 7.580869e-08, 7.537621e-08, 
    7.557014e-08, 7.79518e-08, 7.917028e-08, 8.176382e-08, 8.128895e-08, 
    7.93862e-08, 7.518228e-08, 7.659267e-08, 7.307192e-08, 7.315023e-08, 
    6.935574e-08, 7.104997e-08, 6.48718e-08, 6.658978e-08, 6.170712e-08, 
    6.29116e-08, 6.176329e-08, 6.211003e-08, 6.175878e-08, 6.353165e-08, 
    6.276792e-08, 6.434325e-08, 7.073054e-08, 6.881134e-08, 7.463951e-08, 
    7.829583e-08, 8.078941e-08, 8.258987e-08, 8.233375e-08, 8.184687e-08, 
    7.937514e-08, 7.709681e-08, 7.538971e-08, 7.426181e-08, 7.316149e-08, 
    6.989598e-08, 6.820829e-08, 6.452788e-08, 6.51823e-08, 6.407649e-08, 
    6.30323e-08, 6.130458e-08, 6.158677e-08, 6.08334e-08, 6.410572e-08, 
    6.191801e-08, 6.555697e-08, 6.454779e-08, 7.286297e-08, 7.621053e-08, 
    7.766248e-08, 7.894926e-08, 8.213716e-08, 7.992673e-08, 8.079334e-08, 
    7.874197e-08, 7.745629e-08, 7.809048e-08, 7.423112e-08, 7.571614e-08, 
    6.810912e-08, 7.132027e-08, 6.315349e-08, 6.504764e-08, 6.270509e-08, 
    6.38933e-08, 6.18664e-08, 6.368862e-08, 6.05547e-08, 5.98862e-08, 
    6.034247e-08, 5.860285e-08, 6.379065e-08, 6.176319e-08, 7.810824e-08, 
    7.800455e-08, 7.752283e-08, 7.9655e-08, 7.978675e-08, 8.17768e-08, 
    8.00046e-08, 7.925755e-08, 7.73823e-08, 7.628675e-08, 7.525493e-08, 
    7.301885e-08, 7.057392e-08, 6.724758e-08, 6.492371e-08, 6.33964e-08, 
    6.433012e-08, 6.350529e-08, 6.442777e-08, 6.486326e-08, 6.013602e-08, 
    6.276076e-08, 5.885095e-08, 5.906292e-08, 6.081552e-08, 5.903901e-08, 
    7.793182e-08, 7.852933e-08, 8.062682e-08, 7.898225e-08, 8.199547e-08, 
    8.029951e-08, 7.933478e-08, 7.568463e-08, 7.489812e-08, 7.417326e-08, 
    7.275562e-08, 7.096259e-08, 6.788853e-08, 6.528736e-08, 6.297195e-08, 
    6.313972e-08, 6.308061e-08, 6.257029e-08, 6.383932e-08, 6.23636e-08, 
    6.211808e-08, 6.276122e-08, 5.909135e-08, 6.012466e-08, 5.906744e-08, 
    5.97387e-08, 7.833481e-08, 7.733284e-08, 7.787319e-08, 7.685907e-08, 
    7.757251e-08, 7.443303e-08, 7.35084e-08, 6.928332e-08, 7.099754e-08, 
    6.828276e-08, 7.071865e-08, 7.028281e-08, 6.819488e-08, 7.058564e-08, 
    6.542879e-08, 6.889601e-08, 6.255051e-08, 6.591061e-08, 6.234384e-08, 
    6.298184e-08, 6.192799e-08, 6.099414e-08, 5.983303e-08, 5.772954e-08, 
    5.821216e-08, 5.648228e-08, 7.585499e-08, 7.458426e-08, 7.469581e-08, 
    7.338001e-08, 7.241678e-08, 7.035821e-08, 6.713817e-08, 6.833733e-08, 
    6.614694e-08, 6.571286e-08, 6.904503e-08, 6.698589e-08, 7.374192e-08, 
    7.262083e-08, 7.328713e-08, 7.575409e-08, 6.805943e-08, 7.19399e-08, 
    6.488572e-08, 6.690514e-08, 6.112668e-08, 6.395647e-08, 5.847895e-08, 
    5.623668e-08, 5.418112e-08, 5.184324e-08, 7.389698e-08, 7.475359e-08, 
    7.322463e-08, 7.114318e-08, 6.924807e-08, 6.678074e-08, 6.653178e-08, 
    6.607723e-08, 6.490979e-08, 6.393886e-08, 6.593373e-08, 6.369702e-08, 
    7.236198e-08, 6.772944e-08, 7.507893e-08, 7.281254e-08, 7.126488e-08, 
    7.194132e-08, 6.847534e-08, 6.76749e-08, 6.448635e-08, 6.612193e-08, 
    5.678441e-08, 6.079781e-08, 5.011053e-08, 5.295673e-08, 7.505437e-08, 
    7.390003e-08, 6.997404e-08, 7.182432e-08, 6.661826e-08, 6.537651e-08, 
    6.437872e-08, 6.311782e-08, 6.298285e-08, 6.224474e-08, 6.345731e-08, 
    6.229241e-08, 6.677554e-08, 6.474637e-08, 7.041588e-08, 6.900654e-08, 
    6.965261e-08, 7.036573e-08, 6.818032e-08, 6.590195e-08, 6.585419e-08, 
    6.513483e-08, 6.313545e-08, 6.659771e-08, 5.627922e-08, 6.251296e-08, 
    7.265474e-08, 7.048871e-08, 7.018333e-08, 7.101475e-08, 6.550029e-08, 
    6.746404e-08, 6.226271e-08, 6.364102e-08, 6.139334e-08, 6.250344e-08, 
    6.266787e-08, 6.411592e-08, 6.502859e-08, 6.737308e-08, 6.932187e-08, 
    7.08938e-08, 7.052623e-08, 6.880674e-08, 6.576434e-08, 6.297048e-08, 
    6.357549e-08, 6.156226e-08, 6.698699e-08, 6.467473e-08, 6.556187e-08, 
    6.326567e-08, 6.83693e-08, 6.40055e-08, 6.951559e-08, 6.902037e-08, 
    6.750341e-08, 6.451962e-08, 6.387216e-08, 6.318503e-08, 6.360851e-08, 
    6.568837e-08, 6.603356e-08, 6.754011e-08, 6.795989e-08, 6.912802e-08, 
    7.0105e-08, 6.921191e-08, 6.828213e-08, 6.568763e-08, 6.340653e-08, 
    6.098086e-08, 6.039703e-08, 5.766001e-08, 5.988111e-08, 5.624567e-08, 
    5.932596e-08, 5.40639e-08, 6.375902e-08, 5.941892e-08, 6.743505e-08, 
    6.653871e-08, 6.493738e-08, 6.136331e-08, 6.327634e-08, 6.104313e-08, 
    6.604713e-08, 6.874774e-08, 6.945872e-08, 7.07975e-08, 6.942831e-08, 
    6.953903e-08, 6.824406e-08, 6.865846e-08, 6.560264e-08, 6.723256e-08, 
    6.267192e-08, 6.106064e-08, 5.666181e-08, 5.407382e-08, 5.152355e-08, 
    5.042403e-08, 5.00926e-08, 4.995447e-08,
  1.725312e-09, 1.635417e-09, 1.652616e-09, 1.582135e-09, 1.620953e-09, 
    1.575208e-09, 1.706802e-09, 1.631918e-09, 1.679436e-09, 1.717079e-09, 
    1.45177e-09, 1.579045e-09, 1.327893e-09, 1.402987e-09, 1.220138e-09, 
    1.339371e-09, 1.197099e-09, 1.22347e-09, 1.145415e-09, 1.167382e-09, 
    1.071694e-09, 1.135382e-09, 1.024499e-09, 1.086657e-09, 1.076747e-09, 
    1.13753e-09, 1.552797e-09, 1.467179e-09, 1.557982e-09, 1.54552e-09, 
    1.551104e-09, 1.620141e-09, 1.655779e-09, 1.732338e-09, 1.718249e-09, 
    1.662116e-09, 1.539941e-09, 1.580642e-09, 1.479589e-09, 1.481816e-09, 
    1.374955e-09, 1.422396e-09, 1.251576e-09, 1.298469e-09, 1.166459e-09, 
    1.198659e-09, 1.167955e-09, 1.177203e-09, 1.167835e-09, 1.21533e-09, 
    1.194806e-09, 1.237246e-09, 1.413417e-09, 1.359806e-09, 1.524355e-09, 
    1.630182e-09, 1.703463e-09, 1.756922e-09, 1.74929e-09, 1.734806e-09, 
    1.661791e-09, 1.595262e-09, 1.545908e-09, 1.513535e-09, 1.482137e-09, 
    1.390035e-09, 1.343079e-09, 1.242247e-09, 1.260016e-09, 1.230031e-09, 
    1.201899e-09, 1.155752e-09, 1.163255e-09, 1.143254e-09, 1.23082e-09, 
    1.172079e-09, 1.270221e-09, 1.242786e-09, 1.473652e-09, 1.569585e-09, 
    1.611711e-09, 1.649298e-09, 1.743438e-09, 1.67801e-09, 1.703579e-09, 
    1.643226e-09, 1.605709e-09, 1.624185e-09, 1.512657e-09, 1.555313e-09, 
    1.340334e-09, 1.430006e-09, 1.205155e-09, 1.256354e-09, 1.193121e-09, 
    1.225082e-09, 1.170703e-09, 1.21956e-09, 1.135879e-09, 1.118243e-09, 
    1.130271e-09, 1.084601e-09, 1.222312e-09, 1.167953e-09, 1.624704e-09, 
    1.621679e-09, 1.607645e-09, 1.670015e-09, 1.67389e-09, 1.732724e-09, 
    1.680303e-09, 1.658339e-09, 1.603557e-09, 1.571789e-09, 1.54203e-09, 
    1.47808e-09, 1.409021e-09, 1.316549e-09, 1.252986e-09, 1.211688e-09, 
    1.23689e-09, 1.21462e-09, 1.239534e-09, 1.251344e-09, 1.124825e-09, 
    1.194614e-09, 1.091083e-09, 1.096629e-09, 1.14278e-09, 1.096003e-09, 
    1.619558e-09, 1.637005e-09, 1.698657e-09, 1.650265e-09, 1.739223e-09, 
    1.688996e-09, 1.660606e-09, 1.554404e-09, 1.531775e-09, 1.511002e-09, 
    1.470601e-09, 1.419938e-09, 1.334232e-09, 1.262875e-09, 1.200279e-09, 
    1.204785e-09, 1.203197e-09, 1.18951e-09, 1.223625e-09, 1.183979e-09, 
    1.177418e-09, 1.194626e-09, 1.097373e-09, 1.124525e-09, 1.096747e-09, 
    1.114362e-09, 1.631319e-09, 1.602119e-09, 1.617848e-09, 1.588363e-09, 
    1.609091e-09, 1.518438e-09, 1.492017e-09, 1.372937e-09, 1.420921e-09, 
    1.345141e-09, 1.413083e-09, 1.400859e-09, 1.342708e-09, 1.40935e-09, 
    1.266728e-09, 1.362159e-09, 1.188981e-09, 1.279875e-09, 1.183451e-09, 
    1.200544e-09, 1.172345e-09, 1.147513e-09, 1.116843e-09, 1.061872e-09, 
    1.074417e-09, 1.029642e-09, 1.559317e-09, 1.522771e-09, 1.525969e-09, 
    1.488358e-09, 1.46099e-09, 1.402972e-09, 1.313537e-09, 1.346653e-09, 
    1.286336e-09, 1.274474e-09, 1.366303e-09, 1.309348e-09, 1.498677e-09, 
    1.466776e-09, 1.485713e-09, 1.556407e-09, 1.338958e-09, 1.447492e-09, 
    1.251954e-09, 1.307128e-09, 1.151028e-09, 1.226788e-09, 1.081369e-09, 
    1.023329e-09, 9.709089e-10, 9.122301e-10, 1.503105e-09, 1.527627e-09, 
    1.483934e-09, 1.425019e-09, 1.371955e-09, 1.30371e-09, 1.296878e-09, 
    1.284429e-09, 1.252608e-09, 1.226312e-09, 1.280506e-09, 1.219786e-09, 
    1.459438e-09, 1.329837e-09, 1.536969e-09, 1.472218e-09, 1.428445e-09, 
    1.447532e-09, 1.350479e-09, 1.328331e-09, 1.241121e-09, 1.285651e-09, 
    1.037425e-09, 1.142311e-09, 8.694015e-10, 9.400514e-10, 1.536263e-09, 
    1.503192e-09, 1.392217e-09, 1.444226e-09, 1.29925e-09, 1.265303e-09, 
    1.238206e-09, 1.204197e-09, 1.200572e-09, 1.180802e-09, 1.213327e-09, 
    1.182076e-09, 1.303568e-09, 1.248171e-09, 1.404588e-09, 1.365232e-09, 
    1.383236e-09, 1.403182e-09, 1.342304e-09, 1.279638e-09, 1.278333e-09, 
    1.258725e-09, 1.204672e-09, 1.298686e-09, 1.024423e-09, 1.187977e-09, 
    1.467737e-09, 1.406631e-09, 1.398073e-09, 1.421405e-09, 1.268676e-09, 
    1.322514e-09, 1.181282e-09, 1.218276e-09, 1.15811e-09, 1.18772e-09, 
    1.192124e-09, 1.231096e-09, 1.255836e-09, 1.320006e-09, 1.374011e-09, 
    1.418004e-09, 1.407683e-09, 1.359678e-09, 1.275879e-09, 1.20024e-09, 
    1.216511e-09, 1.162602e-09, 1.309378e-09, 1.246228e-09, 1.270355e-09, 
    1.208171e-09, 1.347539e-09, 1.228113e-09, 1.379412e-09, 1.365617e-09, 
    1.323599e-09, 1.242023e-09, 1.224511e-09, 1.206003e-09, 1.2174e-09, 
    1.273805e-09, 1.283235e-09, 1.324611e-09, 1.336205e-09, 1.368612e-09, 
    1.39588e-09, 1.370948e-09, 1.345124e-09, 1.273785e-09, 1.211961e-09, 
    1.147161e-09, 1.131712e-09, 1.060069e-09, 1.118109e-09, 1.023561e-09, 
    1.103523e-09, 9.679438e-10, 1.221459e-09, 1.105961e-09, 1.321714e-09, 
    1.297068e-09, 1.253358e-09, 1.157313e-09, 1.208458e-09, 1.148812e-09, 
    1.283606e-09, 1.358039e-09, 1.377826e-09, 1.415298e-09, 1.376978e-09, 
    1.380066e-09, 1.344069e-09, 1.355559e-09, 1.271466e-09, 1.316135e-09, 
    1.192232e-09, 1.149277e-09, 1.034265e-09, 9.68194e-10, 9.042847e-10, 
    8.771079e-10, 8.689612e-10, 8.655722e-10,
  1.149871e-11, 1.066712e-11, 1.082501e-11, 1.018166e-11, 1.053478e-11, 
    1.011897e-11, 1.132621e-11, 1.063506e-11, 1.107238e-11, 1.14219e-11, 
    9.018357e-12, 1.015368e-11, 7.946855e-12, 8.592312e-12, 7.043585e-12, 
    8.04468e-12, 6.854115e-12, 7.071096e-12, 6.433948e-12, 6.611695e-12, 
    5.846705e-12, 6.353184e-12, 5.478518e-12, 5.964714e-12, 5.886487e-12, 
    6.370447e-12, 9.916794e-12, 9.154002e-12, 9.963475e-12, 9.851369e-12, 
    9.901569e-12, 1.052736e-11, 1.085412e-11, 1.156436e-11, 1.143281e-11, 
    1.091247e-11, 9.801282e-12, 1.016814e-11, 9.263598e-12, 9.283307e-12, 
    8.349878e-12, 8.761191e-12, 7.30424e-12, 7.697458e-12, 6.604202e-12, 
    6.866905e-12, 6.616352e-12, 6.691566e-12, 6.615376e-12, 7.003934e-12, 
    6.835328e-12, 7.185123e-12, 8.682965e-12, 8.219593e-12, 9.6617e-12, 
    1.061917e-11, 1.129516e-11, 1.179478e-11, 1.172312e-11, 1.158744e-11, 
    1.090948e-11, 1.030074e-11, 9.854855e-12, 9.565093e-12, 9.286143e-12, 
    8.480088e-12, 8.07635e-12, 7.226638e-12, 7.374623e-12, 7.125344e-12, 
    6.893482e-12, 6.517433e-12, 6.578208e-12, 6.416527e-12, 7.131879e-12, 
    6.649868e-12, 7.459955e-12, 7.231115e-12, 9.211129e-12, 1.006815e-11, 
    1.045044e-11, 1.079451e-11, 1.166825e-11, 1.10592e-11, 1.129625e-11, 
    1.073874e-11, 1.039575e-11, 1.056431e-11, 9.557264e-12, 9.939437e-12, 
    8.0529e-12, 8.82763e-12, 6.920218e-12, 7.344063e-12, 6.821537e-12, 
    7.084415e-12, 6.63868e-12, 7.038814e-12, 6.357172e-12, 6.215819e-12, 
    6.312141e-12, 5.948464e-12, 7.061528e-12, 6.616331e-12, 1.056905e-11, 
    1.054141e-11, 1.041338e-11, 1.098533e-11, 1.102111e-11, 1.156796e-11, 
    1.10804e-11, 1.087768e-11, 1.037616e-11, 1.008806e-11, 9.820028e-12, 
    9.250255e-12, 8.644729e-12, 7.850466e-12, 7.315985e-12, 6.973938e-12, 
    7.182173e-12, 6.998081e-12, 7.204112e-12, 7.302306e-12, 6.268478e-12, 
    6.833758e-12, 5.999737e-12, 6.0437e-12, 6.412712e-12, 6.038734e-12, 
    1.052203e-11, 1.068167e-11, 1.125052e-11, 1.080339e-11, 1.162877e-11, 
    1.116089e-11, 1.089857e-11, 9.931264e-12, 9.728089e-12, 9.542511e-12, 
    9.184179e-12, 8.739761e-12, 8.000845e-12, 7.398509e-12, 6.880187e-12, 
    6.917175e-12, 6.904134e-12, 6.791997e-12, 7.072374e-12, 6.746812e-12, 
    6.693319e-12, 6.833854e-12, 6.049606e-12, 6.266074e-12, 6.044637e-12, 
    6.18482e-12, 1.062958e-11, 1.036308e-11, 1.050642e-11, 1.023812e-11, 
    1.042655e-11, 9.608842e-12, 9.373705e-12, 8.3325e-12, 8.748328e-12, 
    8.093974e-12, 8.680058e-12, 8.573849e-12, 8.073184e-12, 8.647581e-12, 
    7.43072e-12, 8.239806e-12, 6.787667e-12, 7.540918e-12, 6.7425e-12, 
    6.882365e-12, 6.652029e-12, 6.450871e-12, 6.204634e-12, 5.769568e-12, 
    5.868129e-12, 5.518338e-12, 9.975511e-12, 9.647544e-12, 9.676131e-12, 
    9.341249e-12, 9.099443e-12, 8.592179e-12, 7.82492e-12, 8.106897e-12, 
    7.595214e-12, 7.495591e-12, 8.275403e-12, 7.789436e-12, 9.432836e-12, 
    9.150438e-12, 9.31781e-12, 9.949294e-12, 8.041159e-12, 8.980783e-12, 
    7.307389e-12, 7.770643e-12, 6.479252e-12, 7.098521e-12, 5.922936e-12, 
    5.469469e-12, 5.068108e-12, 4.628499e-12, 9.472196e-12, 9.690958e-12, 
    9.30205e-12, 8.784083e-12, 8.324039e-12, 7.741737e-12, 7.684031e-12, 
    7.579179e-12, 7.312833e-12, 7.094582e-12, 7.546215e-12, 7.040682e-12, 
    9.085791e-12, 7.9634e-12, 9.774632e-12, 9.19846e-12, 8.813999e-12, 
    8.981127e-12, 8.139636e-12, 7.950575e-12, 7.217291e-12, 7.589459e-12, 
    5.578741e-12, 6.408939e-12, 4.314361e-12, 4.835629e-12, 9.768301e-12, 
    9.472969e-12, 8.49896e-12, 8.952121e-12, 7.704056e-12, 7.418802e-12, 
    7.193089e-12, 6.912346e-12, 6.882589e-12, 6.720891e-12, 6.987437e-12, 
    6.731283e-12, 7.740533e-12, 7.275892e-12, 8.606211e-12, 8.266202e-12, 
    8.421307e-12, 8.594008e-12, 8.069722e-12, 7.538923e-12, 7.527963e-12, 
    7.363847e-12, 6.916259e-12, 7.699294e-12, 5.477935e-12, 6.779473e-12, 
    9.158911e-12, 8.62396e-12, 8.549689e-12, 8.752546e-12, 7.447019e-12, 
    7.901106e-12, 6.724806e-12, 7.028226e-12, 6.53652e-12, 6.777367e-12, 
    6.813375e-12, 7.134162e-12, 7.339742e-12, 7.879809e-12, 8.341745e-12, 
    8.722904e-12, 8.633093e-12, 8.218497e-12, 7.507381e-12, 6.879866e-12, 
    7.013671e-12, 6.572917e-12, 7.789687e-12, 7.259727e-12, 7.461079e-12, 
    6.945002e-12, 8.11448e-12, 7.10949e-12, 8.388301e-12, 8.269506e-12, 
    7.910334e-12, 7.224781e-12, 7.079698e-12, 6.927183e-12, 7.021001e-12, 
    7.489991e-12, 7.569138e-12, 7.918935e-12, 8.017665e-12, 8.295264e-12, 
    8.530681e-12, 8.315367e-12, 8.093824e-12, 7.48982e-12, 6.976186e-12, 
    6.448032e-12, 6.323704e-12, 5.755441e-12, 6.214757e-12, 5.471268e-12, 
    6.098481e-12, 5.045653e-12, 7.054497e-12, 6.117872e-12, 7.894311e-12, 
    7.685636e-12, 7.319086e-12, 6.530069e-12, 6.947362e-12, 6.46136e-12, 
    7.572258e-12, 8.204435e-12, 8.374622e-12, 8.699335e-12, 8.367311e-12, 
    8.393944e-12, 8.084805e-12, 8.183165e-12, 7.47039e-12, 7.846952e-12, 
    6.814263e-12, 6.465108e-12, 5.554189e-12, 5.047543e-12, 4.569782e-12, 
    4.370454e-12, 4.31116e-12, 4.286558e-12,
  1.443577e-14, 1.260062e-14, 1.29434e-14, 1.156402e-14, 1.231542e-14, 
    1.143208e-14, 1.404913e-14, 1.253137e-14, 1.348582e-14, 1.426323e-14, 
    9.192573e-15, 1.150508e-14, 7.162965e-15, 8.366721e-15, 5.582379e-15, 
    7.341595e-15, 5.267456e-15, 5.628598e-15, 4.591195e-15, 4.873476e-15, 
    3.700426e-15, 4.464822e-15, 3.176846e-15, 3.874085e-15, 3.758657e-15, 
    4.491735e-15, 1.100975e-14, 9.460484e-15, 1.110684e-14, 1.08741e-14, 
    1.097814e-14, 1.229949e-14, 1.300689e-14, 1.458369e-14, 1.42877e-14, 
    1.313444e-14, 1.07706e-14, 1.153552e-14, 9.678632e-15, 9.718028e-15, 
    7.907718e-15, 8.691187e-15, 6.025312e-15, 6.713956e-15, 4.861461e-15, 
    5.288517e-15, 4.880947e-15, 5.002149e-15, 4.879382e-15, 5.51597e-15, 
    5.236557e-15, 5.82152e-15, 8.540416e-15, 7.664426e-15, 1.048374e-14, 
    1.249709e-14, 1.397987e-14, 1.510637e-14, 1.494326e-14, 1.463581e-14, 
    1.312789e-14, 1.181582e-14, 1.088131e-14, 1.028657e-14, 9.7237e-15, 
    8.153255e-15, 7.399721e-15, 5.892291e-15, 6.146796e-15, 5.720117e-15, 
    5.332385e-15, 4.723074e-15, 4.819862e-15, 4.563838e-15, 5.731171e-15, 
    4.934837e-15, 6.295132e-15, 5.899935e-15, 9.57402e-15, 1.132547e-14, 
    1.213469e-14, 1.287697e-14, 1.48187e-14, 1.345675e-14, 1.398229e-14, 
    1.275576e-14, 1.20179e-14, 1.23789e-14, 1.027065e-14, 1.105681e-14, 
    7.356667e-15, 8.819887e-15, 5.376634e-15, 6.093951e-15, 5.213914e-15, 
    5.65102e-15, 4.916826e-15, 5.574367e-15, 4.471037e-15, 4.252664e-15, 
    4.401067e-15, 3.850004e-15, 5.612506e-15, 4.880916e-15, 1.23891e-14, 
    1.232966e-14, 1.20555e-14, 1.32942e-14, 1.337287e-14, 1.459183e-14, 
    1.350351e-14, 1.305834e-14, 1.197614e-14, 1.13672e-14, 1.08093e-14, 
    9.651992e-15, 8.467024e-15, 6.988329e-15, 6.045531e-15, 5.465907e-15, 
    5.816501e-15, 5.506187e-15, 5.853853e-15, 6.021984e-15, 4.333581e-15, 
    5.233978e-15, 3.926152e-15, 3.991852e-15, 4.557855e-15, 3.984412e-15, 
    1.228805e-14, 1.263209e-14, 1.388045e-14, 1.28963e-14, 1.472927e-14, 
    1.368148e-14, 1.310401e-14, 1.103982e-14, 1.061988e-14, 1.024065e-14, 
    9.520381e-15, 8.649801e-15, 7.261372e-15, 6.188205e-15, 5.310423e-15, 
    5.37159e-15, 5.349998e-15, 5.165528e-15, 5.630748e-15, 5.091806e-15, 
    5.004989e-15, 5.234133e-15, 4.000707e-15, 4.329872e-15, 3.993257e-15, 
    4.20527e-15, 1.251952e-14, 1.194829e-14, 1.225456e-14, 1.168319e-14, 
    1.208363e-14, 1.037573e-14, 9.899358e-15, 7.875134e-15, 8.666341e-15, 
    7.432127e-15, 8.534826e-15, 8.331482e-15, 7.39391e-15, 8.472483e-15, 
    6.24419e-15, 7.702021e-15, 5.158448e-15, 6.436941e-15, 5.084789e-15, 
    5.31402e-15, 4.938314e-15, 4.617826e-15, 4.235541e-15, 3.588414e-15, 
    3.731742e-15, 3.2321e-15, 1.113191e-14, 1.045478e-14, 1.051329e-14, 
    9.834131e-15, 9.352419e-15, 8.366465e-15, 6.942275e-15, 7.455914e-15, 
    6.53259e-15, 6.357419e-15, 7.768347e-15, 6.87847e-15, 1.001851e-14, 
    9.453399e-15, 9.787116e-15, 1.107732e-14, 7.335137e-15, 9.118765e-15, 
    6.030732e-15, 6.844751e-15, 4.662604e-15, 5.674808e-15, 3.812286e-15, 
    3.164342e-15, 2.62767e-15, 2.083062e-15, 1.009806e-14, 1.054367e-14, 
    9.755538e-15, 8.735471e-15, 7.859275e-15, 6.792996e-15, 6.690047e-15, 
    6.504292e-15, 6.0401e-15, 5.668158e-15, 6.446246e-15, 5.5775e-15, 
    9.325463e-15, 7.193073e-15, 1.071565e-14, 9.548789e-15, 8.793434e-15, 
    9.119435e-15, 7.516298e-15, 7.169722e-15, 5.876332e-15, 6.522429e-15, 
    3.31657e-15, 4.551942e-15, 1.723894e-15, 2.333792e-15, 1.070261e-14, 
    1.009962e-14, 8.189023e-15, 9.062592e-15, 6.725715e-15, 6.22345e-15, 
    5.835076e-15, 5.363595e-15, 5.314389e-15, 5.049675e-15, 5.488416e-15, 
    5.06655e-15, 6.790842e-15, 5.976604e-15, 8.393276e-15, 7.751186e-15, 
    8.042109e-15, 8.369956e-15, 7.387533e-15, 6.433428e-15, 6.414171e-15, 
    6.128148e-15, 5.370096e-15, 6.717228e-15, 3.176053e-15, 5.145078e-15, 
    9.470199e-15, 8.427241e-15, 8.285435e-15, 8.674482e-15, 6.272572e-15, 
    7.0799e-15, 5.05603e-15, 5.556617e-15, 4.753399e-15, 5.141619e-15, 
    5.20053e-15, 5.735034e-15, 6.086491e-15, 7.041343e-15, 7.892461e-15, 
    8.617289e-15, 8.444718e-15, 7.662388e-15, 6.378075e-15, 5.309898e-15, 
    5.532254e-15, 4.811409e-15, 6.878918e-15, 5.948891e-15, 6.297099e-15, 
    5.417761e-15, 7.469888e-15, 5.693337e-15, 7.97992e-15, 7.757345e-15, 
    7.096629e-15, 5.889122e-15, 5.643075e-15, 5.388183e-15, 5.544517e-15, 
    6.347622e-15, 6.486594e-15, 7.112231e-15, 7.292117e-15, 7.805436e-15, 
    8.249266e-15, 7.843036e-15, 7.431848e-15, 6.347318e-15, 5.469658e-15, 
    4.613356e-15, 4.418995e-15, 3.568039e-15, 4.251044e-15, 3.166839e-15, 
    4.074267e-15, 2.598736e-15, 5.600703e-15, 4.10356e-15, 7.067589e-15, 
    6.692904e-15, 6.050878e-15, 4.743149e-15, 5.421683e-15, 4.634363e-15, 
    6.492091e-15, 7.636279e-15, 7.95419e-15, 8.571897e-15, 7.940449e-15, 
    7.99054e-15, 7.415252e-15, 7.596823e-15, 6.31335e-15, 6.981983e-15, 
    5.201987e-15, 4.640274e-15, 3.28214e-15, 2.601161e-15, 2.013953e-15, 
    1.786095e-15, 1.72037e-15, 1.693382e-15,
  5.467507e-20, 4.780206e-20, 4.908677e-20, 4.391401e-20, 4.673277e-20, 
    4.341885e-20, 5.322804e-20, 4.754245e-20, 5.111884e-20, 5.402939e-20, 
    3.500145e-20, 4.369284e-20, 2.734996e-20, 3.189098e-20, 2.137217e-20, 
    2.802441e-20, 2.017882e-20, 2.154725e-20, 1.761317e-20, 1.868465e-20, 
    1.42262e-20, 1.713321e-20, 1.223071e-20, 1.488725e-20, 1.44479e-20, 
    1.723544e-20, 4.183324e-20, 3.600971e-20, 4.219783e-20, 4.132383e-20, 
    4.171454e-20, 4.667302e-20, 4.932468e-20, 5.522854e-20, 5.412099e-20, 
    4.980258e-20, 4.093507e-20, 4.380708e-20, 3.683041e-20, 3.69786e-20, 
    3.016051e-20, 3.311349e-20, 2.304929e-20, 2.56537e-20, 1.863907e-20, 
    2.025865e-20, 1.8713e-20, 1.917281e-20, 1.870706e-20, 2.112057e-20, 
    2.006168e-20, 2.227786e-20, 3.25455e-20, 2.924277e-20, 3.985733e-20, 
    4.741393e-20, 5.296879e-20, 5.718369e-20, 5.657363e-20, 5.542354e-20, 
    4.977806e-20, 4.485886e-20, 4.13509e-20, 3.911633e-20, 3.699993e-20, 
    3.108636e-20, 2.824382e-20, 2.254579e-20, 2.3509e-20, 2.189388e-20, 
    2.042491e-20, 1.811386e-20, 1.848121e-20, 1.750929e-20, 2.193574e-20, 
    1.891746e-20, 2.407017e-20, 2.257473e-20, 3.643688e-20, 4.301867e-20, 
    4.6055e-20, 4.883783e-20, 5.610773e-20, 5.100997e-20, 5.297783e-20, 
    4.838357e-20, 4.561695e-20, 4.69708e-20, 3.905647e-20, 4.200997e-20, 
    2.80813e-20, 3.359824e-20, 2.059261e-20, 2.330905e-20, 1.997584e-20, 
    2.163218e-20, 1.884913e-20, 2.134182e-20, 1.715682e-20, 1.632706e-20, 
    1.689101e-20, 1.479561e-20, 2.148629e-20, 1.871289e-20, 4.700903e-20, 
    4.678614e-20, 4.5758e-20, 5.04011e-20, 5.069581e-20, 5.5259e-20, 
    5.118511e-20, 4.951747e-20, 4.546032e-20, 4.317531e-20, 4.108043e-20, 
    3.67302e-20, 3.226897e-20, 2.669039e-20, 2.312581e-20, 2.093089e-20, 
    2.225885e-20, 2.108351e-20, 2.240027e-20, 2.30367e-20, 1.663458e-20, 
    2.005191e-20, 1.508537e-20, 1.533532e-20, 1.748656e-20, 1.530702e-20, 
    4.663013e-20, 4.792e-20, 5.259658e-20, 4.891026e-20, 5.57732e-20, 
    5.18516e-20, 4.968857e-20, 4.194618e-20, 4.036886e-20, 3.894373e-20, 
    3.623507e-20, 3.29576e-20, 2.772154e-20, 2.366567e-20, 2.034168e-20, 
    2.05735e-20, 2.049167e-20, 1.97924e-20, 2.155539e-20, 1.951285e-20, 
    1.918358e-20, 2.00525e-20, 1.536901e-20, 1.662049e-20, 1.534067e-20, 
    1.61469e-20, 4.749802e-20, 4.535583e-20, 4.650456e-20, 4.436124e-20, 
    4.586349e-20, 3.945142e-20, 3.766057e-20, 3.003762e-20, 3.30199e-20, 
    2.836614e-20, 3.252444e-20, 3.175817e-20, 2.822188e-20, 3.228954e-20, 
    2.387747e-20, 2.938461e-20, 1.976556e-20, 2.460648e-20, 1.948624e-20, 
    2.035531e-20, 1.893066e-20, 1.771429e-20, 1.626197e-20, 1.379962e-20, 
    1.434544e-20, 1.244148e-20, 4.229197e-20, 3.974849e-20, 3.996834e-20, 
    3.741528e-20, 3.560306e-20, 3.189002e-20, 2.651642e-20, 2.845592e-20, 
    2.496813e-20, 2.430575e-20, 2.963482e-20, 2.627536e-20, 3.81086e-20, 
    3.598305e-20, 3.723846e-20, 4.208699e-20, 2.800002e-20, 3.472361e-20, 
    2.306981e-20, 2.614796e-20, 1.78843e-20, 2.172228e-20, 1.465205e-20, 
    1.218301e-20, 1.01332e-20, 8.047706e-21, 3.840769e-20, 4.008251e-20, 
    3.711968e-20, 3.32803e-20, 2.997781e-20, 2.59524e-20, 2.556334e-20, 
    2.486114e-20, 2.310526e-20, 2.169709e-20, 2.464166e-20, 2.135368e-20, 
    3.550161e-20, 2.746365e-20, 4.072864e-20, 3.634195e-20, 3.349862e-20, 
    3.472613e-20, 2.868382e-20, 2.737548e-20, 2.248537e-20, 2.492971e-20, 
    1.276361e-20, 1.746411e-20, 6.668734e-21, 9.00858e-21, 4.067963e-20, 
    3.841356e-20, 3.12212e-20, 3.451214e-20, 2.569814e-20, 2.379901e-20, 
    2.232918e-20, 2.05432e-20, 2.035671e-20, 1.935307e-20, 2.101617e-20, 
    1.941707e-20, 2.594426e-20, 2.286495e-20, 3.199106e-20, 2.957008e-20, 
    3.066731e-20, 3.190318e-20, 2.819781e-20, 2.45932e-20, 2.452037e-20, 
    2.343844e-20, 2.056783e-20, 2.566607e-20, 1.222769e-20, 1.971486e-20, 
    3.604626e-20, 3.211905e-20, 3.158462e-20, 3.305057e-20, 2.398483e-20, 
    2.703627e-20, 1.937717e-20, 2.127457e-20, 1.822897e-20, 1.970174e-20, 
    1.992511e-20, 2.195037e-20, 2.328082e-20, 2.689064e-20, 3.010297e-20, 
    3.283512e-20, 3.218491e-20, 2.923508e-20, 2.438387e-20, 2.033969e-20, 
    2.118227e-20, 1.844913e-20, 2.627706e-20, 2.276005e-20, 2.407761e-20, 
    2.074846e-20, 2.850866e-20, 2.179245e-20, 3.043281e-20, 2.959332e-20, 
    2.709945e-20, 2.253379e-20, 2.160209e-20, 2.063638e-20, 2.122873e-20, 
    2.42687e-20, 2.479423e-20, 2.715837e-20, 2.783762e-20, 2.977473e-20, 
    3.144829e-20, 2.991656e-20, 2.836509e-20, 2.426755e-20, 2.09451e-20, 
    1.769732e-20, 1.695912e-20, 1.3722e-20, 1.63209e-20, 1.219253e-20, 
    1.564879e-20, 1.002254e-20, 2.144158e-20, 1.576019e-20, 2.698977e-20, 
    2.557414e-20, 2.314605e-20, 1.819006e-20, 2.076332e-20, 1.777708e-20, 
    2.481501e-20, 2.913657e-20, 3.033578e-20, 3.266411e-20, 3.028395e-20, 
    3.047285e-20, 2.830245e-20, 2.898769e-20, 2.413908e-20, 2.666642e-20, 
    1.993063e-20, 1.779952e-20, 1.263233e-20, 1.003182e-20, 7.782614e-21, 
    6.907777e-21, 6.655187e-21, 6.551434e-21,
  4.403182e-26, 3.851916e-26, 3.954979e-26, 3.539946e-26, 3.766128e-26, 
    3.500208e-26, 4.28714e-26, 3.831089e-26, 4.117978e-26, 4.351404e-26, 
    2.824416e-26, 3.522196e-26, 2.209567e-26, 2.574541e-26, 1.728716e-26, 
    2.263788e-26, 1.632652e-26, 1.742807e-26, 1.426024e-26, 1.512333e-26, 
    1.153032e-26, 1.387355e-26, 9.920511e-27, 1.206335e-26, 1.17091e-26, 
    1.395592e-26, 3.372948e-26, 2.905394e-26, 3.402211e-26, 3.332059e-26, 
    3.36342e-26, 3.761334e-26, 3.974064e-26, 4.447563e-26, 4.358749e-26, 
    4.0124e-26, 3.300853e-26, 3.531364e-26, 2.971302e-26, 2.983202e-26, 
    2.435485e-26, 2.672761e-26, 1.863676e-26, 2.073171e-26, 1.508661e-26, 
    1.639079e-26, 1.514616e-26, 1.551647e-26, 1.514138e-26, 1.708466e-26, 
    1.623221e-26, 1.801603e-26, 2.627129e-26, 2.361725e-26, 3.214337e-26, 
    3.820778e-26, 4.266349e-26, 4.604329e-26, 4.555416e-26, 4.463199e-26, 
    4.010432e-26, 3.615767e-26, 3.334232e-26, 3.154848e-26, 2.984916e-26, 
    2.509888e-26, 2.281427e-26, 1.823163e-26, 1.900661e-26, 1.770703e-26, 
    1.652465e-26, 1.466357e-26, 1.495947e-26, 1.417654e-26, 1.774072e-26, 
    1.531083e-26, 1.945805e-26, 1.825492e-26, 2.939699e-26, 3.468091e-26, 
    3.711747e-26, 3.935009e-26, 4.51806e-26, 4.109245e-26, 4.267074e-26, 
    3.898568e-26, 3.676598e-26, 3.785225e-26, 3.150042e-26, 3.387133e-26, 
    2.268362e-26, 2.711703e-26, 1.665966e-26, 1.884575e-26, 1.61631e-26, 
    1.749642e-26, 1.52558e-26, 1.726273e-26, 1.389257e-26, 1.322394e-26, 
    1.36784e-26, 1.198946e-26, 1.737901e-26, 1.514607e-26, 3.788292e-26, 
    3.77041e-26, 3.687916e-26, 4.060409e-26, 4.084047e-26, 4.450005e-26, 
    4.123293e-26, 3.989529e-26, 3.664031e-26, 3.480662e-26, 3.312521e-26, 
    2.963255e-26, 2.604911e-26, 2.156535e-26, 1.869832e-26, 1.693198e-26, 
    1.800074e-26, 1.705483e-26, 1.811454e-26, 1.862663e-26, 1.347177e-26, 
    1.622434e-26, 1.222308e-26, 1.242458e-26, 1.415824e-26, 1.240177e-26, 
    3.757893e-26, 3.861378e-26, 4.236498e-26, 3.94082e-26, 4.491236e-26, 
    4.176749e-26, 4.003254e-26, 3.382013e-26, 3.255401e-26, 3.140991e-26, 
    2.923493e-26, 2.660236e-26, 2.23944e-26, 1.913265e-26, 1.645764e-26, 
    1.664427e-26, 1.657839e-26, 1.601539e-26, 1.743463e-26, 1.579029e-26, 
    1.552514e-26, 1.622482e-26, 1.245174e-26, 1.346041e-26, 1.242889e-26, 
    1.307875e-26, 3.827524e-26, 3.655647e-26, 3.747818e-26, 3.575836e-26, 
    3.696381e-26, 3.18175e-26, 3.037964e-26, 2.425609e-26, 2.665242e-26, 
    2.29126e-26, 2.625437e-26, 2.563871e-26, 2.279663e-26, 2.606564e-26, 
    1.930304e-26, 2.373125e-26, 1.599378e-26, 1.988945e-26, 1.576887e-26, 
    1.646861e-26, 1.532145e-26, 1.43417e-26, 1.317149e-26, 1.118628e-26, 
    1.162647e-26, 1.00906e-26, 3.409767e-26, 3.2056e-26, 3.223249e-26, 
    3.018267e-26, 2.872735e-26, 2.574464e-26, 2.142546e-26, 2.298477e-26, 
    2.018034e-26, 1.964756e-26, 2.393236e-26, 2.123163e-26, 3.073939e-26, 
    2.903253e-26, 3.004069e-26, 3.393314e-26, 2.261828e-26, 2.8021e-26, 
    1.865326e-26, 2.112918e-26, 1.447866e-26, 1.756894e-26, 1.187371e-26, 
    9.88201e-27, 8.226951e-27, 6.541249e-27, 3.097953e-26, 3.232415e-26, 
    2.994532e-26, 2.686161e-26, 2.420802e-26, 2.097192e-26, 2.065904e-26, 
    2.009429e-26, 1.868179e-26, 1.754866e-26, 1.991775e-26, 1.727229e-26, 
    2.864588e-26, 2.218707e-26, 3.284283e-26, 2.932076e-26, 2.7037e-26, 
    2.802303e-26, 2.316797e-26, 2.211618e-26, 1.818302e-26, 2.014944e-26, 
    1.035053e-26, 1.414015e-26, 5.425323e-27, 7.318186e-27, 3.280348e-26, 
    3.098424e-26, 2.520723e-26, 2.785114e-26, 2.076745e-26, 1.923992e-26, 
    1.805733e-26, 1.661988e-26, 1.646974e-26, 1.566163e-26, 1.700063e-26, 
    1.571317e-26, 2.096537e-26, 1.848843e-26, 2.582582e-26, 2.388033e-26, 
    2.476213e-26, 2.575521e-26, 2.277729e-26, 1.987877e-26, 1.982019e-26, 
    1.894985e-26, 1.663971e-26, 2.074166e-26, 9.918069e-27, 1.595295e-26, 
    2.90833e-26, 2.592866e-26, 2.549925e-26, 2.667706e-26, 1.93894e-26, 
    2.184345e-26, 1.568104e-26, 1.720861e-26, 1.475629e-26, 1.594239e-26, 
    1.612224e-26, 1.775249e-26, 1.882303e-26, 2.172636e-26, 2.430861e-26, 
    2.650397e-26, 2.598158e-26, 2.361107e-26, 1.971039e-26, 1.645604e-26, 
    1.713432e-26, 1.493363e-26, 2.123299e-26, 1.840403e-26, 1.946404e-26, 
    1.678513e-26, 2.302717e-26, 1.762541e-26, 2.457368e-26, 2.3899e-26, 
    2.189425e-26, 1.822198e-26, 1.747221e-26, 1.669489e-26, 1.717172e-26, 
    1.961775e-26, 2.004046e-26, 2.194163e-26, 2.248772e-26, 2.404481e-26, 
    2.538971e-26, 2.415879e-26, 2.291175e-26, 1.961683e-26, 1.694342e-26, 
    1.432803e-26, 1.373328e-26, 1.112368e-26, 1.321898e-26, 9.889698e-27, 
    1.267727e-26, 8.137562e-27, 1.734303e-26, 1.276706e-26, 2.180607e-26, 
    2.066772e-26, 1.87146e-26, 1.472496e-26, 1.679709e-26, 1.439228e-26, 
    2.005718e-26, 2.353189e-26, 2.44957e-26, 2.636658e-26, 2.445406e-26, 
    2.460586e-26, 2.28614e-26, 2.341222e-26, 1.951348e-26, 2.154608e-26, 
    1.612669e-26, 1.441036e-26, 1.02446e-26, 8.145055e-27, 6.326815e-27, 
    5.618854e-27, 5.414353e-27, 5.33034e-27,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_SAT =
  0.00476377, 0.004763827, 0.004763817, 0.004763857, 0.004763837, 
    0.004763862, 0.004763784, 0.004763827, 0.004763802, 0.004763779, 
    0.004763919, 0.00476386, 0.004764045, 0.004764012, 0.004764092, 
    0.004764037, 0.004764103, 0.004764096, 0.004764127, 0.004764119, 
    0.00476414, 0.00476413, 0.004764156, 0.004764141, 0.004764142, 
    0.004764129, 0.004763877, 0.004763911, 0.004763874, 0.004763879, 
    0.004763878, 0.004763836, 0.00476381, 0.004763769, 0.004763778, 
    0.00476381, 0.004763882, 0.004763862, 0.00476392, 0.004763919, 
    0.004764027, 0.00476395, 0.004764084, 0.004764065, 0.004764119, 
    0.004764107, 0.004764118, 0.004764115, 0.004764118, 0.004764099, 
    0.004764107, 0.004764091, 0.004763953, 0.004764033, 0.004763892, 
    0.004763823, 0.004763785, 0.004763753, 0.004763757, 0.004763765, 
    0.00476381, 0.004763853, 0.004763883, 0.004763901, 0.004763919, 
    0.00476401, 0.004764038, 0.004764086, 0.004764082, 0.004764091, 
    0.004764105, 0.004764121, 0.00476412, 0.004764125, 0.004764094, 
    0.004764114, 0.004764079, 0.004764089, 0.004763906, 0.004763868, 
    0.004763835, 0.004763818, 0.004763761, 0.0047638, 0.004763784, 
    0.004763825, 0.004763847, 0.004763837, 0.004763902, 0.004763877, 
    0.00476404, 0.004763943, 0.004764104, 0.004764083, 0.004764109, 
    0.004764097, 0.004764115, 0.004764099, 0.004764129, 0.004764132, 
    0.004764129, 0.004764145, 0.004764098, 0.004764116, 0.004763836, 
    0.004763837, 0.004763846, 0.004763805, 0.004763803, 0.004763768, 
    0.004763801, 0.004763813, 0.00476385, 0.004763867, 0.004763884, 
    0.004763919, 0.004763953, 0.004764053, 0.004764084, 0.004764102, 
    0.004764093, 0.004764101, 0.004764091, 0.004764087, 0.00476413, 
    0.004764106, 0.004764143, 0.004764142, 0.004764125, 0.004764142, 
    0.004763839, 0.004763829, 0.004763789, 0.004763821, 0.004763764, 
    0.004763794, 0.004763809, 0.004763874, 0.004763891, 0.004763901, 
    0.004763925, 0.004763951, 0.004764045, 0.004764078, 0.004764107, 
    0.004764105, 0.004764106, 0.00476411, 0.004764097, 0.004764112, 
    0.004764113, 0.004764108, 0.004764142, 0.004764133, 0.004764142, 
    0.004764137, 0.004763833, 0.00476385, 0.00476384, 0.004763857, 
    0.004763843, 0.004763893, 0.004763907, 0.004764024, 0.004763949, 
    0.00476404, 0.004763954, 0.004764013, 0.004764033, 0.004764012, 
    0.004764073, 0.004764027, 0.00476411, 0.004764063, 0.004764112, 
    0.004764107, 0.004764117, 0.004764124, 0.004764135, 0.004764148, 
    0.004764146, 0.004764157, 0.004763875, 0.004763893, 0.004763894, 
    0.004763915, 0.004763928, 0.004764014, 0.004764056, 0.004764043, 
    0.004764071, 0.004764075, 0.004764033, 0.004764057, 0.004763907, 
    0.004763921, 0.004763915, 0.004763874, 0.004764041, 0.004763932, 
    0.004764084, 0.00476406, 0.004764123, 0.004764091, 0.004764144, 
    0.004764151, 0.004764169, 0.004764169, 0.004763906, 0.004763894, 
    0.004763918, 0.004763944, 0.004764029, 0.004764061, 0.004764066, 
    0.004764071, 0.004764086, 0.004764096, 0.004764069, 0.004764099, 
    0.004763918, 0.004764047, 0.004763886, 0.004763917, 0.004763944, 
    0.004763936, 0.004764042, 0.004764052, 0.004764087, 0.004764072, 
    0.004764147, 0.004764121, 0.004764176, 0.004764168, 0.004763888, 
    0.004763907, 0.004764017, 0.004763938, 0.004764065, 0.004764079, 
    0.004764092, 0.004764103, 0.004764106, 0.004764112, 0.004764102, 
    0.004764113, 0.004764061, 0.004764087, 0.004764015, 0.004764032, 
    0.004764026, 0.004764015, 0.004764045, 0.004764068, 0.004764074, 
    0.00476408, 0.004764085, 0.004764065, 0.00476414, 0.004764094, 
    0.004763927, 0.004764006, 0.004764016, 0.004763952, 0.004764077, 
    0.004764053, 0.004764113, 0.0047641, 0.004764122, 0.004764111, 
    0.004764109, 0.004764094, 0.004764083, 0.004764053, 0.004764027, 
    0.004763953, 0.004764013, 0.004764034, 0.004764071, 0.004764104, 
    0.004764097, 0.004764121, 0.00476406, 0.004764085, 0.004764074, 
    0.004764103, 0.004764041, 0.004764079, 0.004764027, 0.004764034, 
    0.004764053, 0.004764083, 0.004764097, 0.004764102, 0.0047641, 
    0.004764073, 0.004764071, 0.004764054, 0.004764046, 0.004764033, 
    0.004764019, 0.00476403, 0.00476404, 0.004764075, 0.004764099, 
    0.004764124, 0.004764131, 0.004764139, 0.004764126, 0.004764139, 
    0.004764117, 0.004764155, 0.004764088, 0.004764127, 0.004764055, 
    0.004764067, 0.00476408, 0.004764115, 0.004764103, 0.00476412, 
    0.004764071, 0.004764032, 0.004764028, 0.004763954, 0.004764028, 
    0.004764027, 0.004764045, 0.00476404, 0.004764076, 0.004764058, 
    0.004764108, 0.004764121, 0.004764155, 0.004764164, 0.004764177, 
    0.004764178, 0.004764178, 0.004764178,
  9.944767e-06, 9.956249e-06, 9.954025e-06, 9.963253e-06, 9.958147e-06, 
    9.964177e-06, 9.94711e-06, 9.956692e-06, 9.950585e-06, 9.945818e-06, 
    9.981065e-06, 9.963666e-06, 9.999262e-06, 9.988205e-06, 1.001596e-05, 
    9.997527e-06, 1.001967e-05, 1.001546e-05, 1.00282e-05, 1.002455e-05, 
    1.004074e-05, 1.002988e-05, 1.004915e-05, 1.003817e-05, 1.003988e-05, 
    1.002951e-05, 9.967201e-06, 9.978894e-06, 9.9665e-06, 9.968172e-06, 
    9.967429e-06, 9.958243e-06, 9.953587e-06, 9.943908e-06, 9.945672e-06, 
    9.952792e-06, 9.968924e-06, 9.963473e-06, 9.977251e-06, 9.976941e-06, 
    9.992295e-06, 9.985332e-06, 1.001101e-05, 1.000376e-05, 1.002471e-05, 
    1.001945e-05, 1.002445e-05, 1.002294e-05, 1.002447e-05, 1.001676e-05, 
    1.002006e-05, 1.001328e-05, 9.986616e-06, 9.99452e-06, 9.971054e-06, 
    9.95689e-06, 9.947526e-06, 9.940846e-06, 9.941791e-06, 9.943586e-06, 
    9.952832e-06, 9.961532e-06, 9.96814e-06, 9.972551e-06, 9.976897e-06, 
    9.990034e-06, 9.996987e-06, 1.001247e-05, 1.00097e-05, 1.00144e-05, 
    1.001892e-05, 1.002647e-05, 1.002523e-05, 1.002855e-05, 1.00143e-05, 
    1.002376e-05, 1.000812e-05, 1.00124e-05, 9.977982e-06, 9.964949e-06, 
    9.959314e-06, 9.954449e-06, 9.942515e-06, 9.950755e-06, 9.947506e-06, 
    9.955251e-06, 9.96015e-06, 9.957732e-06, 9.972672e-06, 9.966866e-06, 
    9.997398e-06, 9.984227e-06, 1.00184e-05, 1.001027e-05, 1.002034e-05, 
    1.001521e-05, 1.002399e-05, 1.001609e-05, 1.002979e-05, 1.003275e-05, 
    1.003072e-05, 1.003854e-05, 1.001565e-05, 1.002445e-05, 9.957659e-06, 
    9.958054e-06, 9.9599e-06, 9.951777e-06, 9.951284e-06, 9.943854e-06, 
    9.950475e-06, 9.953284e-06, 9.960442e-06, 9.964652e-06, 9.968658e-06, 
    9.977452e-06, 9.987235e-06, 1.000099e-05, 1.00108e-05, 1.001735e-05, 
    1.001334e-05, 1.001688e-05, 1.001292e-05, 1.001106e-05, 1.003164e-05, 
    1.002009e-05, 1.003742e-05, 1.003646e-05, 1.002862e-05, 1.003657e-05, 
    9.958332e-06, 9.956061e-06, 9.948137e-06, 9.954339e-06, 9.943045e-06, 
    9.949359e-06, 9.952978e-06, 9.966967e-06, 9.970057e-06, 9.97289e-06, 
    9.978503e-06, 9.985683e-06, 9.998328e-06, 1.000924e-05, 1.001919e-05, 
    1.001846e-05, 1.001872e-05, 1.002093e-05, 1.001544e-05, 1.002183e-05, 
    1.002289e-05, 1.00201e-05, 1.003634e-05, 1.003171e-05, 1.003644e-05, 
    1.003343e-05, 9.956801e-06, 9.960626e-06, 9.958559e-06, 9.962439e-06, 
    9.959698e-06, 9.971848e-06, 9.975483e-06, 9.992566e-06, 9.985537e-06, 
    9.996693e-06, 9.986671e-06, 9.988513e-06, 9.997013e-06, 9.9873e-06, 
    1.000862e-05, 9.994142e-06, 1.002101e-05, 1.000656e-05, 1.002192e-05, 
    1.001915e-05, 1.002374e-05, 1.002784e-05, 1.003301e-05, 1.004249e-05, 
    1.00403e-05, 1.004824e-05, 9.966328e-06, 9.971268e-06, 9.97085e-06, 
    9.976026e-06, 9.979845e-06, 9.988219e-06, 1.000146e-05, 9.99649e-06, 
    1.000562e-05, 1.000745e-05, 9.993581e-06, 1.000208e-05, 9.974583e-06, 
    9.979007e-06, 9.976387e-06, 9.966708e-06, 9.997611e-06, 9.981728e-06, 
    1.001095e-05, 1.000244e-05, 1.002725e-05, 1.001491e-05, 1.003909e-05, 
    1.004934e-05, 1.005904e-05, 1.007025e-05, 9.97398e-06, 9.970625e-06, 
    9.976647e-06, 9.98493e-06, 9.992737e-06, 1.000295e-05, 1.000401e-05, 
    1.000591e-05, 1.001086e-05, 1.001501e-05, 1.00065e-05, 1.001606e-05, 
    9.979995e-06, 9.998987e-06, 9.969339e-06, 9.978239e-06, 9.98445e-06, 
    9.981745e-06, 9.995927e-06, 9.999236e-06, 1.001265e-05, 1.000573e-05, 
    1.00468e-05, 1.002868e-05, 1.007882e-05, 1.006486e-05, 9.969447e-06, 
    9.973977e-06, 9.989761e-06, 9.982216e-06, 1.000364e-05, 1.000887e-05, 
    1.001313e-05, 1.001854e-05, 1.001914e-05, 1.002234e-05, 1.001709e-05, 
    1.002214e-05, 1.000297e-05, 1.001155e-05, 9.987991e-06, 9.993728e-06, 
    9.991096e-06, 9.988194e-06, 9.997142e-06, 1.000663e-05, 1.000686e-05, 
    1.000989e-05, 1.001836e-05, 1.000373e-05, 1.004907e-05, 1.002108e-05, 
    9.978909e-06, 9.987653e-06, 9.988924e-06, 9.985481e-06, 1.000835e-05, 
    1.00001e-05, 1.002227e-05, 1.00163e-05, 1.002608e-05, 1.002122e-05, 
    1.00205e-05, 1.001425e-05, 1.001035e-05, 1.000048e-05, 9.992433e-06, 
    9.985973e-06, 9.987542e-06, 9.994544e-06, 1.000721e-05, 1.001918e-05, 
    1.001656e-05, 1.002534e-05, 1.00021e-05, 1.001185e-05, 1.000807e-05, 
    1.001791e-05, 9.996352e-06, 1.001463e-05, 9.991656e-06, 9.993681e-06, 
    9.99994e-06, 1.001249e-05, 1.00153e-05, 1.001825e-05, 1.001644e-05, 
    1.000754e-05, 1.000609e-05, 9.999795e-06, 9.998041e-06, 9.993243e-06, 
    9.989253e-06, 9.992891e-06, 9.996703e-06, 1.000755e-05, 1.001729e-05, 
    1.002789e-05, 1.003049e-05, 1.004276e-05, 1.003274e-05, 1.004922e-05, 
    1.003515e-05, 1.005951e-05, 1.001573e-05, 1.00348e-05, 1.000023e-05, 
    1.000398e-05, 1.001071e-05, 1.002618e-05, 1.001787e-05, 1.00276e-05, 
    1.000604e-05, 9.99477e-06, 9.991886e-06, 9.986355e-06, 9.992011e-06, 
    9.991559e-06, 9.996881e-06, 9.995173e-06, 1.000791e-05, 1.000108e-05, 
    1.002048e-05, 1.002753e-05, 1.00474e-05, 1.005951e-05, 1.007185e-05, 
    1.007727e-05, 1.007892e-05, 1.007961e-05,
  2.18823e-10, 2.192973e-10, 2.192053e-10, 2.195874e-10, 2.193758e-10, 
    2.196257e-10, 2.189196e-10, 2.193158e-10, 2.190631e-10, 2.188663e-10, 
    2.203273e-10, 2.196045e-10, 2.210832e-10, 2.206218e-10, 2.21782e-10, 
    2.210109e-10, 2.219376e-10, 2.217607e-10, 2.222954e-10, 2.221423e-10, 
    2.228238e-10, 2.22366e-10, 2.231786e-10, 2.22715e-10, 2.227872e-10, 
    2.223508e-10, 2.197509e-10, 2.20237e-10, 2.197219e-10, 2.197913e-10, 
    2.197604e-10, 2.193799e-10, 2.191874e-10, 2.187874e-10, 2.188602e-10, 
    2.191544e-10, 2.198225e-10, 2.195964e-10, 2.201681e-10, 2.201553e-10, 
    2.207923e-10, 2.205043e-10, 2.215745e-10, 2.21271e-10, 2.221487e-10, 
    2.219279e-10, 2.221381e-10, 2.220745e-10, 2.22139e-10, 2.218151e-10, 
    2.219538e-10, 2.216692e-10, 2.205578e-10, 2.208852e-10, 2.199109e-10, 
    2.193242e-10, 2.189368e-10, 2.186611e-10, 2.187001e-10, 2.187742e-10, 
    2.191561e-10, 2.195159e-10, 2.197898e-10, 2.199729e-10, 2.201534e-10, 
    2.206984e-10, 2.209882e-10, 2.216354e-10, 2.215195e-10, 2.217165e-10, 
    2.219059e-10, 2.222228e-10, 2.221708e-10, 2.223101e-10, 2.217119e-10, 
    2.221092e-10, 2.214532e-10, 2.216325e-10, 2.201991e-10, 2.196575e-10, 
    2.194245e-10, 2.192229e-10, 2.1873e-10, 2.190702e-10, 2.18936e-10, 
    2.19256e-10, 2.194588e-10, 2.193586e-10, 2.199779e-10, 2.19737e-10, 
    2.210054e-10, 2.204584e-10, 2.218838e-10, 2.215433e-10, 2.219656e-10, 
    2.217503e-10, 2.221189e-10, 2.217872e-10, 2.223623e-10, 2.224871e-10, 
    2.224017e-10, 2.227307e-10, 2.217687e-10, 2.221378e-10, 2.193556e-10, 
    2.19372e-10, 2.194483e-10, 2.191125e-10, 2.190921e-10, 2.187852e-10, 
    2.190586e-10, 2.191747e-10, 2.194708e-10, 2.196453e-10, 2.198114e-10, 
    2.201765e-10, 2.205837e-10, 2.211553e-10, 2.215654e-10, 2.2184e-10, 
    2.216718e-10, 2.218203e-10, 2.216542e-10, 2.215765e-10, 2.224401e-10, 
    2.219549e-10, 2.226834e-10, 2.226432e-10, 2.223133e-10, 2.226478e-10, 
    2.193835e-10, 2.192895e-10, 2.18962e-10, 2.192183e-10, 2.187518e-10, 
    2.190125e-10, 2.191622e-10, 2.197414e-10, 2.198694e-10, 2.19987e-10, 
    2.202202e-10, 2.20519e-10, 2.210441e-10, 2.215003e-10, 2.219171e-10, 
    2.218866e-10, 2.218973e-10, 2.219901e-10, 2.217598e-10, 2.220279e-10, 
    2.220726e-10, 2.219553e-10, 2.226378e-10, 2.224429e-10, 2.226424e-10, 
    2.225155e-10, 2.193201e-10, 2.194784e-10, 2.193928e-10, 2.195536e-10, 
    2.194401e-10, 2.199439e-10, 2.200949e-10, 2.208038e-10, 2.205129e-10, 
    2.209759e-10, 2.205601e-10, 2.206347e-10, 2.209895e-10, 2.20584e-10, 
    2.214745e-10, 2.208696e-10, 2.219937e-10, 2.213885e-10, 2.220315e-10, 
    2.219153e-10, 2.221081e-10, 2.222803e-10, 2.224976e-10, 2.228975e-10, 
    2.228051e-10, 2.2314e-10, 2.197147e-10, 2.199197e-10, 2.199023e-10, 
    2.201172e-10, 2.202761e-10, 2.206224e-10, 2.211748e-10, 2.209673e-10, 
    2.213489e-10, 2.214253e-10, 2.208459e-10, 2.21201e-10, 2.200574e-10, 
    2.202413e-10, 2.201323e-10, 2.197305e-10, 2.210142e-10, 2.203545e-10, 
    2.21572e-10, 2.212156e-10, 2.222557e-10, 2.217379e-10, 2.22754e-10, 
    2.231866e-10, 2.235964e-10, 2.240718e-10, 2.200323e-10, 2.198929e-10, 
    2.20143e-10, 2.204878e-10, 2.208107e-10, 2.212373e-10, 2.212812e-10, 
    2.213609e-10, 2.215681e-10, 2.21742e-10, 2.213855e-10, 2.217857e-10, 
    2.202828e-10, 2.210717e-10, 2.198397e-10, 2.202095e-10, 2.204677e-10, 
    2.203551e-10, 2.209437e-10, 2.210819e-10, 2.21643e-10, 2.213533e-10, 
    2.230793e-10, 2.223158e-10, 2.244358e-10, 2.238433e-10, 2.198441e-10, 
    2.200321e-10, 2.206867e-10, 2.203747e-10, 2.21266e-10, 2.214848e-10, 
    2.216631e-10, 2.2189e-10, 2.21915e-10, 2.220495e-10, 2.21829e-10, 
    2.22041e-10, 2.212382e-10, 2.215971e-10, 2.206128e-10, 2.208521e-10, 
    2.207422e-10, 2.206213e-10, 2.209945e-10, 2.21391e-10, 2.214005e-10, 
    2.215274e-10, 2.218833e-10, 2.212697e-10, 2.231759e-10, 2.219972e-10, 
    2.20237e-10, 2.205991e-10, 2.206518e-10, 2.205105e-10, 2.214628e-10, 
    2.211182e-10, 2.220464e-10, 2.217958e-10, 2.222066e-10, 2.220024e-10, 
    2.219723e-10, 2.217102e-10, 2.215467e-10, 2.211338e-10, 2.20798e-10, 
    2.205309e-10, 2.205942e-10, 2.208861e-10, 2.214155e-10, 2.219168e-10, 
    2.218069e-10, 2.221754e-10, 2.212015e-10, 2.216094e-10, 2.214514e-10, 
    2.218635e-10, 2.209615e-10, 2.217266e-10, 2.207656e-10, 2.208501e-10, 
    2.211114e-10, 2.216364e-10, 2.21754e-10, 2.218778e-10, 2.218017e-10, 
    2.214291e-10, 2.213685e-10, 2.211052e-10, 2.210321e-10, 2.208317e-10, 
    2.206654e-10, 2.208171e-10, 2.209762e-10, 2.214297e-10, 2.218376e-10, 
    2.222826e-10, 2.223919e-10, 2.229091e-10, 2.224867e-10, 2.231823e-10, 
    2.225888e-10, 2.23617e-10, 2.217724e-10, 2.225734e-10, 2.211236e-10, 
    2.212801e-10, 2.21562e-10, 2.222107e-10, 2.218616e-10, 2.222703e-10, 
    2.213662e-10, 2.208957e-10, 2.207752e-10, 2.205469e-10, 2.207804e-10, 
    2.207615e-10, 2.209836e-10, 2.209123e-10, 2.214447e-10, 2.211588e-10, 
    2.219712e-10, 2.222674e-10, 2.231045e-10, 2.236168e-10, 2.241397e-10, 
    2.2437e-10, 2.244401e-10, 2.244694e-10,
  4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13,
  4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13,
  3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13,
  3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13,
  3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_UNSAT =
  2.496702, 2.473692, 2.478171, 2.459572, 2.469896, 2.457708, 2.492044, 
    2.472776, 2.485082, 2.494635, 2.42335, 2.458741, 2.386434, 2.409123, 
    2.352012, 2.389967, 2.344339, 2.353112, 2.326687, 2.334266, 2.300375, 
    2.323187, 2.28276, 2.305829, 2.302223, 2.323939, 2.451634, 2.427763, 
    2.453045, 2.449646, 2.451172, 2.469682, 2.478991, 2.49846, 2.49493, 
    2.480629, 2.448118, 2.459171, 2.43129, 2.431921, 2.40077, 2.41483, 
    2.362298, 2.377262, 2.33395, 2.344862, 2.334462, 2.337618, 2.334421, 
    2.35042, 2.343569, 2.357635, 2.412198, 2.396198, 2.443823, 2.472322, 
    2.491199, 2.504566, 2.502678, 2.499076, 2.480546, 2.463085, 2.449752, 
    2.440821, 2.432012, 2.405281, 2.391104, 2.359267, 2.365024, 2.355271, 
    2.345948, 2.330268, 2.332851, 2.325936, 2.355531, 2.335872, 2.3683, 
    2.359443, 2.429606, 2.456191, 2.467456, 2.47731, 2.501225, 2.484717, 
    2.491229, 2.47573, 2.465865, 2.470746, 2.440577, 2.452319, 2.390262, 
    2.41705, 2.347036, 2.363843, 2.343003, 2.353643, 2.335402, 2.351821, 
    2.323361, 2.317151, 2.321395, 2.305083, 2.35273, 2.334461, 2.470882, 
    2.470087, 2.466378, 2.482665, 2.48366, 2.498556, 2.485304, 2.479653, 
    2.465293, 2.456786, 2.44869, 2.430863, 2.410904, 2.382917, 2.362754, 
    2.349211, 2.357519, 2.350185, 2.358382, 2.362222, 2.319478, 2.343505, 
    2.307431, 2.309432, 2.325771, 2.309206, 2.469528, 2.474107, 2.489981, 
    2.477561, 2.500177, 2.487525, 2.48024, 2.452072, 2.445872, 2.440116, 
    2.428737, 2.414111, 2.388388, 2.365944, 2.345405, 2.346912, 2.346381, 
    2.341786, 2.353163, 2.339917, 2.337691, 2.343508, 2.309699, 2.319372, 
    2.309474, 2.315773, 2.472619, 2.464911, 2.469077, 2.461241, 2.466762, 
    2.442184, 2.4348, 2.400163, 2.414398, 2.391734, 2.4121, 2.408494, 
    2.39099, 2.411001, 2.367182, 2.396912, 2.341607, 2.371382, 2.339738, 
    2.345494, 2.335963, 2.327416, 2.316654, 2.29676, 2.301371, 2.28471, 
    2.453408, 2.443385, 2.444269, 2.433769, 2.425994, 2.409119, 2.381979, 
    2.392196, 2.373432, 2.36966, 2.398164, 2.380673, 2.436671, 2.427648, 
    2.433022, 2.452617, 2.389841, 2.422117, 2.36242, 2.379978, 2.328635, 
    2.354206, 2.303908, 2.282315, 2.261954, 2.238093, 2.437911, 2.444727, 
    2.43252, 2.415596, 2.399868, 2.378908, 2.376762, 2.372828, 2.362632, 
    2.354048, 2.371582, 2.351896, 2.42555, 2.387034, 2.447302, 2.429198, 
    2.416596, 2.422128, 2.393363, 2.386569, 2.358901, 2.373215, 2.287648, 
    2.325608, 2.219891, 2.249555, 2.447107, 2.437935, 2.40593, 2.421174, 
    2.377508, 2.366724, 2.357949, 2.346716, 2.345503, 2.33884, 2.349756, 
    2.339272, 2.378864, 2.361194, 2.409596, 2.39784, 2.403251, 2.409181, 
    2.390866, 2.371306, 2.37089, 2.364608, 2.346875, 2.377331, 2.282732, 
    2.341269, 2.427922, 2.4102, 2.407669, 2.41454, 2.367806, 2.384769, 
    2.339003, 2.351396, 2.331081, 2.341182, 2.342667, 2.355621, 2.363675, 
    2.383991, 2.400486, 2.413544, 2.41051, 2.39616, 2.370109, 2.345392, 
    2.350812, 2.332627, 2.380682, 2.360563, 2.368344, 2.348041, 2.392467, 
    2.354642, 2.402107, 2.397956, 2.385105, 2.359195, 2.353456, 2.347318, 
    2.351106, 2.369447, 2.372449, 2.385419, 2.388995, 2.39886, 2.407018, 
    2.399564, 2.391729, 2.36944, 2.349302, 2.327294, 2.321901, 2.296094, 
    2.317104, 2.282404, 2.311908, 2.260777, 2.352449, 2.31278, 2.384521, 
    2.376822, 2.362875, 2.330807, 2.348137, 2.327867, 2.372567, 2.395663, 
    2.401631, 2.41275, 2.401377, 2.402303, 2.391406, 2.394909, 2.368699, 
    2.382788, 2.342703, 2.328028, 2.286457, 2.260876, 2.234768, 2.223218, 
    2.2197, 2.218229,
  1.658949, 1.637626, 1.641774, 1.624554, 1.634111, 1.62283, 1.65463, 
    1.636777, 1.648178, 1.657033, 1.591069, 1.623785, 1.557021, 1.577941, 
    1.525343, 1.560276, 1.518292, 1.526355, 1.502084, 1.50904, 1.477956, 
    1.498872, 1.46183, 1.482954, 1.47965, 1.499561, 1.617211, 1.595145, 
    1.618516, 1.615372, 1.616784, 1.633912, 1.642533, 1.660579, 1.657306, 
    1.644051, 1.613958, 1.624183, 1.598406, 1.598989, 1.570236, 1.583207, 
    1.534802, 1.548575, 1.50875, 1.518773, 1.50922, 1.512118, 1.509183, 
    1.523881, 1.517585, 1.530514, 1.580778, 1.566021, 1.609988, 1.636355, 
    1.653847, 1.666243, 1.664491, 1.66115, 1.643974, 1.627806, 1.615471, 
    1.607213, 1.599073, 1.574394, 1.561324, 1.532015, 1.537311, 1.52834, 
    1.51977, 1.50537, 1.507741, 1.501393, 1.528579, 1.510514, 1.540326, 
    1.532177, 1.596847, 1.621426, 1.63185, 1.640977, 1.663144, 1.647839, 
    1.653874, 1.639514, 1.630379, 1.634898, 1.606987, 1.617845, 1.560549, 
    1.585256, 1.52077, 1.536224, 1.517064, 1.526844, 1.510083, 1.525169, 
    1.499031, 1.493334, 1.497227, 1.482271, 1.526004, 1.509219, 1.635024, 
    1.634287, 1.630855, 1.645937, 1.64686, 1.660669, 1.648383, 1.643147, 
    1.629851, 1.621977, 1.614489, 1.598011, 1.579584, 1.553782, 1.535222, 
    1.52277, 1.530407, 1.523665, 1.531202, 1.534734, 1.495468, 1.517525, 
    1.484423, 1.486257, 1.501242, 1.48605, 1.63377, 1.638011, 1.652718, 
    1.64121, 1.662172, 1.650441, 1.64369, 1.617616, 1.611883, 1.606561, 
    1.596048, 1.582543, 1.558822, 1.538157, 1.519272, 1.520657, 1.520169, 
    1.515947, 1.526402, 1.51423, 1.512185, 1.517529, 1.486502, 1.495371, 
    1.486296, 1.492071, 1.636633, 1.629497, 1.633353, 1.6261, 1.631209, 
    1.608472, 1.601648, 1.569676, 1.582808, 1.561906, 1.580687, 1.57736, 
    1.561219, 1.579674, 1.539295, 1.566677, 1.515783, 1.543159, 1.514065, 
    1.519354, 1.510598, 1.502752, 1.492879, 1.474646, 1.47887, 1.463615, 
    1.618852, 1.609583, 1.610401, 1.600696, 1.593514, 1.577937, 1.552919, 
    1.562332, 1.545049, 1.541577, 1.567833, 1.551715, 1.603377, 1.59504, 
    1.600006, 1.61812, 1.56016, 1.589933, 1.534915, 1.551076, 1.503871, 
    1.52736, 1.481194, 1.461422, 1.442809, 1.42103, 1.604523, 1.610825, 
    1.599542, 1.583913, 1.569404, 1.55009, 1.548114, 1.544492, 1.53511, 
    1.527217, 1.543345, 1.525237, 1.593102, 1.557575, 1.613204, 1.596472, 
    1.584836, 1.589944, 1.563408, 1.557147, 1.531677, 1.54485, 1.466302, 
    1.501091, 1.404444, 1.431486, 1.613025, 1.604546, 1.574994, 1.589063, 
    1.548801, 1.538875, 1.530803, 1.520476, 1.519362, 1.51324, 1.52327, 
    1.513638, 1.550049, 1.533787, 1.578378, 1.567535, 1.572525, 1.577995, 
    1.561106, 1.543091, 1.542709, 1.536927, 1.520619, 1.548638, 1.461801, 
    1.515469, 1.595294, 1.578933, 1.576599, 1.582939, 1.53987, 1.555488, 
    1.51339, 1.524778, 1.506116, 1.515392, 1.516756, 1.528662, 1.53607, 
    1.554772, 1.569974, 1.58202, 1.57922, 1.565985, 1.541989, 1.51926, 
    1.52424, 1.507535, 1.551724, 1.533206, 1.540365, 1.521694, 1.562581, 
    1.527759, 1.571469, 1.567642, 1.555798, 1.531947, 1.526671, 1.52103, 
    1.524512, 1.54138, 1.544143, 1.556087, 1.559382, 1.568476, 1.575999, 
    1.569125, 1.561901, 1.541374, 1.522853, 1.50264, 1.497692, 1.474034, 
    1.493289, 1.461501, 1.488523, 1.441732, 1.525744, 1.489324, 1.55526, 
    1.548169, 1.535332, 1.505863, 1.521782, 1.503165, 1.544252, 1.565526, 
    1.571031, 1.581288, 1.570796, 1.57165, 1.561604, 1.564833, 1.540692, 
    1.553664, 1.516789, 1.503313, 1.465213, 1.441824, 1.418, 1.407474, 
    1.40427, 1.402931,
  0.6537312, 0.6421599, 0.6444065, 0.635097, 0.6402584, 0.6341671, 0.6513826, 
    0.6417007, 0.6478785, 0.6526888, 0.617111, 0.6346825, 0.5989814, 
    0.6101015, 0.5822594, 0.6007078, 0.5785563, 0.5827914, 0.5700713, 
    0.5737086, 0.5575102, 0.5683945, 0.5491617, 0.5601057, 0.5583894, 
    0.5687542, 0.6311395, 0.6192923, 0.6318426, 0.6301499, 0.6309097, 
    0.640151, 0.6448176, 0.6546185, 0.6528373, 0.6456405, 0.6293892, 
    0.6348971, 0.6210387, 0.621351, 0.6059986, 0.6129102, 0.5872379, 
    0.5945091, 0.5735567, 0.5788089, 0.5738029, 0.5753199, 0.5737831, 
    0.5814908, 0.5781853, 0.5849793, 0.611614, 0.6037577, 0.6272542, 
    0.6414724, 0.650957, 0.6577032, 0.6567487, 0.6549293, 0.6455984, 
    0.6368521, 0.6302031, 0.6257634, 0.6213959, 0.6082122, 0.6012637, 
    0.5857693, 0.58856, 0.5838353, 0.5793321, 0.5717886, 0.5730288, 
    0.5697108, 0.5839609, 0.5744803, 0.5901507, 0.5858546, 0.6202038, 
    0.6334105, 0.6390367, 0.6439743, 0.6560148, 0.6476947, 0.6509718, 
    0.6431822, 0.6382416, 0.6406844, 0.6256421, 0.6314809, 0.6008524, 
    0.614004, 0.5798569, 0.5879871, 0.5779124, 0.5830485, 0.5742545, 
    0.5821676, 0.5684776, 0.5655065, 0.5675363, 0.5597508, 0.5826068, 
    0.5738024, 0.6407526, 0.640354, 0.6384985, 0.646663, 0.6471635, 
    0.6546671, 0.64799, 0.6451505, 0.637956, 0.6337073, 0.6296744, 0.620827, 
    0.6109774, 0.5972652, 0.5874592, 0.5809072, 0.5849231, 0.5813771, 
    0.5853412, 0.5872016, 0.5666189, 0.5781542, 0.560869, 0.5618222, 
    0.5696318, 0.5617148, 0.6400743, 0.6423682, 0.6503437, 0.6441004, 
    0.6554853, 0.6491069, 0.6454446, 0.6313575, 0.6282727, 0.6254132, 
    0.6197755, 0.6125559, 0.5999364, 0.5890064, 0.5790706, 0.5797974, 
    0.5795414, 0.5773264, 0.5828162, 0.5764263, 0.575355, 0.5781562, 
    0.5619499, 0.5665686, 0.5618425, 0.5648487, 0.6416225, 0.6377649, 
    0.6398487, 0.635931, 0.6386901, 0.6264396, 0.6227765, 0.6057009, 
    0.6126975, 0.6015724, 0.6115658, 0.609792, 0.6012078, 0.6110252, 
    0.5896067, 0.6041066, 0.5772403, 0.5916468, 0.5763402, 0.5791135, 
    0.5745241, 0.5704206, 0.5652695, 0.5557936, 0.5579846, 0.5500841, 
    0.6320236, 0.6270363, 0.6274762, 0.6222662, 0.6184188, 0.6100994, 
    0.5968079, 0.6017987, 0.592645, 0.5908109, 0.604721, 0.5961705, 
    0.6237042, 0.619236, 0.6218963, 0.6316292, 0.6006462, 0.6165033, 
    0.5872972, 0.5958323, 0.5710051, 0.5833197, 0.5591913, 0.5489511, 
    0.5393628, 0.5282077, 0.6243193, 0.6277038, 0.6216475, 0.6132874, 
    0.6055562, 0.5953107, 0.5942653, 0.5923509, 0.5874, 0.5832443, 0.5917448, 
    0.5822037, 0.6181985, 0.5992748, 0.6289834, 0.6200027, 0.61378, 
    0.6165092, 0.6023699, 0.5990479, 0.5855917, 0.5925395, 0.5514731, 
    0.5695533, 0.5197591, 0.5335546, 0.628887, 0.6243315, 0.6085317, 
    0.6160383, 0.5946288, 0.5893851, 0.5851313, 0.5797024, 0.5791179, 
    0.5759079, 0.5811701, 0.576116, 0.595289, 0.5867029, 0.6103344, 
    0.6045624, 0.6072166, 0.6101301, 0.601148, 0.5916104, 0.5914088, 
    0.588358, 0.5797779, 0.5945424, 0.549147, 0.5770761, 0.619372, 0.6106305, 
    0.6093864, 0.6127674, 0.5899103, 0.598169, 0.5759864, 0.5819624, 
    0.5721791, 0.5770354, 0.5777507, 0.5840047, 0.5879059, 0.5977895, 
    0.6058595, 0.612277, 0.6107836, 0.6037388, 0.5910286, 0.5790641, 
    0.5816798, 0.5729212, 0.5961753, 0.5863969, 0.5901712, 0.5803422, 
    0.601931, 0.5835298, 0.6066548, 0.6046194, 0.5983333, 0.5857338, 
    0.5829575, 0.5799933, 0.5818223, 0.5907071, 0.5921665, 0.5984863, 
    0.6002331, 0.6050626, 0.6090668, 0.6054077, 0.6015699, 0.5907041, 
    0.5809507, 0.570362, 0.5677786, 0.5554767, 0.5654835, 0.548992, 
    0.5630015, 0.5388092, 0.5824702, 0.5634184, 0.5980482, 0.5942945, 
    0.5875172, 0.5720467, 0.5803883, 0.5706366, 0.5922238, 0.6034951, 
    0.6064215, 0.6118861, 0.6062967, 0.606751, 0.6014123, 0.6031268, 
    0.5903441, 0.5972027, 0.5777682, 0.5707139, 0.5509101, 0.5388565, 
    0.5266611, 0.5212998, 0.519671, 0.5189905,
  0.1245632, 0.1212687, 0.1219058, 0.1192736, 0.1207304, 0.1190118, 
    0.1238919, 0.1211387, 0.1228928, 0.1242651, 0.1142472, 0.1191569, 
    0.1092601, 0.1123095, 0.1047318, 0.1097316, 0.1037383, 0.1048747, 
    0.1014748, 0.1024429, 0.09815709, 0.1010296, 0.09597393, 0.09883936, 
    0.09838802, 0.1011251, 0.1181609, 0.1148527, 0.1183583, 0.1178833, 
    0.1180964, 0.1207, 0.1220226, 0.1248171, 0.1243075, 0.1222563, 0.11767, 
    0.1192173, 0.1153381, 0.115425, 0.1111808, 0.1130844, 0.1060727, 
    0.1080422, 0.1024024, 0.1038059, 0.102468, 0.1028728, 0.1024628, 
    0.1045253, 0.1036389, 0.1054636, 0.1127266, 0.1105661, 0.1170722, 
    0.1210741, 0.1237704, 0.1257014, 0.1254275, 0.1249061, 0.1222444, 
    0.1197682, 0.1178981, 0.1166554, 0.1154375, 0.1117893, 0.1098835, 
    0.1056765, 0.1064298, 0.1051555, 0.1039461, 0.1019315, 0.1022617, 
    0.101379, 0.1051893, 0.1026487, 0.1068601, 0.1056995, 0.115106, 
    0.1187989, 0.120385, 0.1217832, 0.1252171, 0.1228405, 0.1237747, 
    0.1215585, 0.1201604, 0.1208509, 0.1166215, 0.1182567, 0.1097711, 
    0.1133868, 0.1040868, 0.106275, 0.1035659, 0.1049438, 0.1025885, 
    0.104707, 0.1010517, 0.1002645, 0.1008021, 0.09874594, 0.1048251, 
    0.1024679, 0.1208702, 0.1207574, 0.1202329, 0.122547, 0.1226894, 
    0.124831, 0.1229246, 0.1221171, 0.1200797, 0.1188824, 0.1177499, 
    0.1152792, 0.1125509, 0.1087922, 0.1061324, 0.1043685, 0.1054484, 
    0.1044947, 0.1055611, 0.1060629, 0.100559, 0.1036306, 0.09904031, 
    0.09929151, 0.101358, 0.09926319, 0.1206783, 0.1213277, 0.1235954, 
    0.121819, 0.1250654, 0.1232428, 0.1222007, 0.1182221, 0.1173572, 
    0.1165576, 0.1149868, 0.1129866, 0.1095208, 0.1065505, 0.103876, 
    0.1040708, 0.1040022, 0.1034091, 0.1048814, 0.1031684, 0.1028822, 
    0.1036311, 0.09932517, 0.1005456, 0.09929685, 0.1000905, 0.1211165, 
    0.1200258, 0.1206145, 0.1195085, 0.1202871, 0.1168444, 0.115822, 
    0.1110991, 0.1130257, 0.1099679, 0.1127133, 0.1122242, 0.1098683, 
    0.1125641, 0.1067129, 0.1106618, 0.103386, 0.1072654, 0.1031454, 
    0.1038875, 0.1026604, 0.1015676, 0.1002018, 0.09770674, 0.09828162, 
    0.09621423, 0.1184091, 0.1170113, 0.1171343, 0.1156798, 0.11461, 
    0.1123089, 0.1086676, 0.1100298, 0.107536, 0.1070389, 0.1108302, 
    0.1084941, 0.1160806, 0.114837, 0.1155768, 0.1182984, 0.1097147, 
    0.1140787, 0.1060887, 0.108402, 0.101723, 0.1050168, 0.09859879, 
    0.09591912, 0.09343401, 0.09057239, 0.1162522, 0.117198, 0.1155075, 
    0.1131887, 0.1110594, 0.1082602, 0.107976, 0.1074563, 0.1061164, 
    0.1049965, 0.1072919, 0.1047167, 0.1145489, 0.1093401, 0.1175563, 
    0.11505, 0.1133249, 0.1140803, 0.1101861, 0.1092782, 0.1056286, 
    0.1075074, 0.09657665, 0.1013372, 0.08842628, 0.09194009, 0.1175293, 
    0.1162556, 0.1118772, 0.1139498, 0.1080747, 0.1066529, 0.1055045, 
    0.1040454, 0.1038887, 0.1030299, 0.1044391, 0.1030855, 0.1082542, 
    0.1059283, 0.1123736, 0.1107867, 0.1115154, 0.1123173, 0.1098518, 
    0.1072555, 0.1072009, 0.1063753, 0.1040658, 0.1080513, 0.09597021, 
    0.1033422, 0.1148747, 0.1124553, 0.1121125, 0.113045, 0.106795, 
    0.1090385, 0.1030508, 0.1046519, 0.1020354, 0.1033312, 0.1035226, 
    0.1052011, 0.1062531, 0.108935, 0.1111426, 0.1129095, 0.1124975, 
    0.110561, 0.1070979, 0.1038743, 0.104576, 0.102233, 0.1084954, 0.1058457, 
    0.1068657, 0.1042169, 0.110066, 0.1050734, 0.1113611, 0.1108024, 
    0.1090833, 0.105667, 0.1049194, 0.1041234, 0.1046143, 0.1070108, 
    0.1074063, 0.109125, 0.1096018, 0.1109239, 0.1120244, 0.1110186, 
    0.1099672, 0.1070099, 0.1043803, 0.1015521, 0.1008663, 0.09762375, 
    0.1002585, 0.09592988, 0.09960273, 0.09329136, 0.1047884, 0.09971271, 
    0.1090055, 0.1079839, 0.1061481, 0.1020002, 0.1042293, 0.1016251, 
    0.1074218, 0.1104942, 0.111297, 0.1128016, 0.1112627, 0.1113875, 
    0.1099241, 0.1103933, 0.1069125, 0.1087751, 0.1035273, 0.1016456, 
    0.09642966, 0.09330347, 0.09017811, 0.08881623, 0.08840396, 0.0882319,
  0.008816758, 0.008484081, 0.0085481, 0.008284585, 0.008430102, 0.008258518, 
    0.008748644, 0.008471033, 0.008647579, 0.008786486, 0.007788677, 
    0.008272961, 0.007306243, 0.00760007, 0.00687666, 0.007351434, 
    0.006783509, 0.006890095, 0.006572763, 0.006662642, 0.00626765, 
    0.006531558, 0.006069354, 0.006330024, 0.006288739, 0.006540385, 
    0.008173973, 0.007847899, 0.008193562, 0.008146449, 0.008167575, 
    0.008427064, 0.008559853, 0.008842562, 0.008790793, 0.008583385, 
    0.008125324, 0.008278972, 0.007895476, 0.007904003, 0.007490894, 
    0.00767532, 0.007003014, 0.007189902, 0.006658875, 0.006789835, 
    0.006664982, 0.006702679, 0.006664491, 0.006857261, 0.006774212, 
    0.006945525, 0.007640543, 0.007431643, 0.008066203, 0.008464553, 
    0.008736336, 0.008932628, 0.008904701, 0.008851619, 0.00858218, 
    0.008333901, 0.00814792, 0.008025063, 0.00790523, 0.007549698, 
    0.007366015, 0.006965607, 0.007036788, 0.006916513, 0.006802959, 
    0.006615113, 0.006645791, 0.006563894, 0.006919692, 0.006681802, 
    0.007077544, 0.006967772, 0.007872723, 0.008237339, 0.008395539, 
    0.008535764, 0.008883267, 0.0086423, 0.008736765, 0.008513173, 
    0.008373071, 0.008442176, 0.008021721, 0.00818348, 0.007355223, 
    0.007704746, 0.006816138, 0.007022141, 0.00676738, 0.006896591, 
    0.006676192, 0.006874332, 0.006533598, 0.006460938, 0.006510529, 
    0.00632147, 0.006885427, 0.00666497, 0.008444111, 0.008432812, 
    0.008380321, 0.008612683, 0.008627042, 0.008843978, 0.008650787, 
    0.008569364, 0.008365007, 0.008245642, 0.008133238, 0.007889697, 
    0.007623494, 0.007261473, 0.00700866, 0.006842553, 0.006944097, 
    0.006854394, 0.006954719, 0.007002085, 0.006488091, 0.006773434, 
    0.00634843, 0.006371465, 0.006561949, 0.006368867, 0.008424887, 
    0.008489999, 0.008718612, 0.00853936, 0.00886782, 0.008682934, 
    0.008577781, 0.008180047, 0.00809437, 0.008015418, 0.007861031, 
    0.007665806, 0.007331217, 0.007048215, 0.006796397, 0.00681464, 
    0.006808213, 0.006752722, 0.006890719, 0.006730249, 0.006703555, 
    0.006773483, 0.006374554, 0.006486855, 0.006371955, 0.006444907, 
    0.008468801, 0.008359618, 0.008418498, 0.008307998, 0.008385734, 
    0.008043713, 0.00794301, 0.007483012, 0.00766961, 0.007374118, 
    0.007639249, 0.007591804, 0.007364555, 0.00762477, 0.0070636, 
    0.007440858, 0.006750572, 0.007116015, 0.0067281, 0.006797472, 
    0.006682888, 0.006581366, 0.006455158, 0.00622658, 0.006279018, 
    0.006091082, 0.008198606, 0.008060184, 0.008072334, 0.007929027, 
    0.007824135, 0.007600012, 0.007249568, 0.007380057, 0.007141724, 
    0.007094502, 0.007457077, 0.007232999, 0.007968441, 0.007846355, 
    0.007918911, 0.008187614, 0.007349814, 0.00777221, 0.007004528, 
    0.007224213, 0.006595774, 0.006903461, 0.006308007, 0.006064404, 
    0.005841166, 0.005587362, 0.007985328, 0.008078628, 0.007912106, 
    0.007685468, 0.007479176, 0.007210678, 0.007183591, 0.00713414, 
    0.007007146, 0.006901545, 0.007118529, 0.006875245, 0.007818169, 
    0.007313905, 0.008114066, 0.00786723, 0.007698717, 0.007772364, 
    0.007395076, 0.00730797, 0.00696109, 0.007139003, 0.006123902, 
    0.006560024, 0.005399325, 0.005708231, 0.00811139, 0.007985661, 
    0.007558193, 0.007759626, 0.007193001, 0.007057913, 0.006949384, 
    0.006812259, 0.006797582, 0.006717325, 0.006849176, 0.006722509, 
    0.007210114, 0.006989371, 0.00760629, 0.007452888, 0.007523207, 
    0.007600831, 0.00736297, 0.007115072, 0.007109877, 0.007031625, 
    0.006814176, 0.007190765, 0.006069025, 0.00674649, 0.007850046, 
    0.007614219, 0.007580976, 0.007671484, 0.007071377, 0.007285026, 
    0.006719279, 0.006869154, 0.006624762, 0.006745453, 0.006763333, 
    0.006920801, 0.007020068, 0.007275129, 0.007487208, 0.007658318, 
    0.007618302, 0.007431143, 0.007100102, 0.006796237, 0.006862029, 
    0.006643126, 0.007233119, 0.006981579, 0.007078077, 0.006828336, 
    0.007383537, 0.006908793, 0.007508292, 0.007454393, 0.007289311, 
    0.006964708, 0.006894291, 0.006819567, 0.006865619, 0.007091837, 
    0.007129389, 0.007293303, 0.007338983, 0.007466109, 0.007572448, 
    0.00747524, 0.00737405, 0.007091757, 0.006843654, 0.006579923, 
    0.006516461, 0.006219026, 0.006460385, 0.006065381, 0.006400051, 
    0.005828438, 0.006881988, 0.006410153, 0.007281872, 0.007184347, 
    0.007010147, 0.006621498, 0.006829496, 0.006586691, 0.007130866, 
    0.007424721, 0.007502102, 0.007647833, 0.007498793, 0.007510843, 
    0.007369907, 0.007415004, 0.007082512, 0.007259839, 0.006763772, 
    0.006588595, 0.006110583, 0.005829515, 0.005552664, 0.005433342, 
    0.005397379, 0.005382393,
  0.0001783912, 0.0001690617, 0.0001708464, 0.0001635332, 0.0001675609, 
    0.0001628146, 0.0001764699, 0.0001686986, 0.0001736297, 0.0001775366, 
    0.0001500111, 0.0001632127, 0.0001371677, 0.0001449526, 0.0001260006, 
    0.0001383574, 0.0001236136, 0.0001263459, 0.0001182596, 0.000120535, 
    0.0001106247, 0.0001172204, 0.0001057383, 0.0001121741, 0.0001111479, 
    0.0001174428, 0.0001604896, 0.0001516092, 0.0001610275, 0.0001597347, 
    0.0001603141, 0.0001674765, 0.0001711746, 0.0001791204, 0.0001776581, 
    0.0001718322, 0.000159156, 0.0001633784, 0.0001528961, 0.0001531271, 
    0.0001420463, 0.0001469651, 0.0001292582, 0.0001341179, 0.0001204394, 
    0.0001237752, 0.0001205944, 0.0001215524, 0.000120582, 0.0001255024, 
    0.000123376, 0.0001277732, 0.0001460341, 0.0001404758, 0.0001575393, 
    0.0001685185, 0.0001761233, 0.0001816723, 0.00018088, 0.0001793766, 
    0.0001717986, 0.0001648952, 0.000159775, 0.000156417, 0.0001531604, 
    0.0001436098, 0.0001387418, 0.0001282914, 0.0001301328, 0.0001270256, 
    0.0001241109, 0.0001193303, 0.0001201075, 0.0001180357, 0.0001271074, 
    0.0001210216, 0.0001311903, 0.0001283473, 0.0001522804, 0.0001622313, 
    0.0001666019, 0.0001705021, 0.0001802726, 0.0001734817, 0.0001761354, 
    0.000169872, 0.0001659791, 0.0001678962, 0.0001563259, 0.0001607506, 
    0.0001384573, 0.0001477542, 0.0001244483, 0.0001297533, 0.0001232015, 
    0.0001265129, 0.0001208791, 0.0001259407, 0.0001172718, 0.0001154452, 
    0.000116691, 0.0001119612, 0.0001262258, 0.0001205941, 0.00016795, 
    0.0001676361, 0.00016618, 0.000172652, 0.0001730541, 0.0001791605, 
    0.0001737197, 0.0001714403, 0.0001657558, 0.0001624599, 0.0001593727, 
    0.0001527397, 0.0001455783, 0.0001359919, 0.0001294043, 0.0001251251, 
    0.0001277364, 0.0001254288, 0.0001280104, 0.0001292342, 0.0001161269, 
    0.0001233561, 0.0001126324, 0.0001132068, 0.0001179866, 0.000113142, 
    0.000167416, 0.0001692264, 0.0001756246, 0.0001706024, 0.0001798351, 
    0.0001746218, 0.0001716756, 0.0001606564, 0.0001583089, 0.0001561542, 
    0.000151964, 0.0001467103, 0.0001378248, 0.0001304291, 0.000123943, 
    0.0001244099, 0.0001242454, 0.0001228274, 0.0001263619, 0.0001222544, 
    0.0001215747, 0.0001233574, 0.0001132839, 0.0001160958, 0.000113219, 
    0.0001150433, 0.0001686365, 0.0001656067, 0.0001672387, 0.0001641794, 
    0.00016633, 0.0001569255, 0.0001541851, 0.0001418372, 0.0001468122, 
    0.0001389556, 0.0001459995, 0.000144732, 0.0001387034, 0.0001456123, 
    0.0001308283, 0.0001407198, 0.0001227725, 0.0001321908, 0.0001221996, 
    0.0001239706, 0.0001210492, 0.0001184769, 0.0001153002, 0.0001096077, 
    0.0001109066, 0.0001062707, 0.0001611661, 0.000157375, 0.0001577067, 
    0.0001538056, 0.0001509672, 0.0001449511, 0.0001356796, 0.0001391123, 
    0.0001328604, 0.000131631, 0.0001411493, 0.0001352455, 0.0001548759, 
    0.0001515673, 0.0001535313, 0.0001608641, 0.0001383147, 0.0001495675, 
    0.0001292974, 0.0001350154, 0.000118841, 0.0001266897, 0.0001116265, 
    0.0001056171, 0.0001001909, 9.411835e-05, 0.0001553351, 0.0001578786, 
    0.0001533467, 0.0001472371, 0.0001417353, 0.0001346611, 0.000133953, 
    0.0001326628, 0.0001293651, 0.0001266403, 0.0001322562, 0.0001259642, 
    0.0001508063, 0.0001373692, 0.0001588478, 0.0001521317, 0.0001475924, 
    0.0001495716, 0.0001395089, 0.0001372131, 0.0001281748, 0.0001327895, 
    0.0001070765, 0.0001179381, 8.968722e-05, 9.69973e-05, 0.0001587745, 
    0.0001553441, 0.000143836, 0.0001492288, 0.0001341989, 0.0001306807, 
    0.0001278727, 0.000124349, 0.0001239734, 0.0001219252, 0.000125295, 
    0.0001220572, 0.0001346464, 0.0001289053, 0.0001451187, 0.0001410384, 
    0.0001429048, 0.0001449729, 0.0001386615, 0.0001321662, 0.000132031, 
    0.000129999, 0.0001243982, 0.0001341404, 0.0001057304, 0.0001226686, 
    0.000151667, 0.0001453305, 0.0001444432, 0.0001468623, 0.0001310302, 
    0.0001366101, 0.0001219749, 0.0001258077, 0.0001195746, 0.000122642, 
    0.0001230982, 0.000127136, 0.0001296996, 0.0001363502, 0.0001419485, 
    0.0001465097, 0.0001454395, 0.0001404626, 0.0001317767, 0.000123939, 
    0.0001256248, 0.0001200399, 0.0001352486, 0.000128704, 0.0001312042, 
    0.0001247607, 0.0001392042, 0.000126827, 0.0001425084, 0.0001410782, 
    0.0001367226, 0.0001282683, 0.0001264537, 0.0001245361, 0.000125717, 
    0.0001315618, 0.000132539, 0.0001368275, 0.0001380293, 0.0001413888, 
    0.0001442158, 0.0001416309, 0.0001389538, 0.0001315597, 0.0001251534, 
    0.0001184404, 0.0001168403, 0.000109421, 0.0001154314, 0.0001056411, 
    0.0001139208, 9.9884e-05, 0.0001261375, 0.0001141733, 0.0001365272, 
    0.0001339727, 0.0001294428, 0.000119492, 0.0001247904, 0.0001186115, 
    0.0001325775, 0.0001402927, 0.0001423439, 0.0001462291, 0.000142256, 
    0.0001425762, 0.0001388445, 0.0001400356, 0.0001313194, 0.000135949, 
    0.0001231094, 0.0001186596, 0.0001067493, 9.990989e-05, 9.329624e-05, 
    9.048446e-05, 8.964166e-05, 8.929107e-05,
  1.13769e-06, 1.055365e-06, 1.070995e-06, 1.007312e-06, 1.042265e-06, 
    1.001106e-06, 1.120612e-06, 1.052192e-06, 1.095483e-06, 1.130085e-06, 
    8.92176e-07, 1.004542e-06, 7.861449e-07, 8.500142e-07, 6.967758e-07, 
    7.958245e-07, 6.780314e-07, 6.994975e-07, 6.36466e-07, 6.540494e-07, 
    5.783774e-07, 6.284766e-07, 5.4196e-07, 5.900501e-07, 5.823123e-07, 
    6.301843e-07, 9.810952e-07, 9.056001e-07, 9.857157e-07, 9.746196e-07, 
    9.795883e-07, 1.04153e-06, 1.073876e-06, 1.144188e-06, 1.131166e-06, 
    1.079653e-06, 9.696622e-07, 1.005974e-06, 9.164464e-07, 9.183969e-07, 
    8.260241e-07, 8.667262e-07, 7.225634e-07, 7.614684e-07, 6.533081e-07, 
    6.792966e-07, 6.5451e-07, 6.619507e-07, 6.544135e-07, 6.92853e-07, 
    6.761728e-07, 7.107786e-07, 8.58985e-07, 8.131321e-07, 9.558471e-07, 
    1.050619e-06, 1.117538e-06, 1.167001e-06, 1.159907e-06, 1.146474e-06, 
    1.079357e-06, 1.019098e-06, 9.749647e-07, 9.462854e-07, 9.186776e-07, 
    8.38909e-07, 7.989582e-07, 7.148859e-07, 7.29527e-07, 7.048644e-07, 
    6.819259e-07, 6.447246e-07, 6.507366e-07, 6.347427e-07, 7.05511e-07, 
    6.578257e-07, 7.379696e-07, 7.153288e-07, 9.112538e-07, 9.960761e-07, 
    1.033917e-06, 1.067976e-06, 1.154474e-06, 1.094178e-06, 1.117645e-06, 
    1.062455e-06, 1.028503e-06, 1.045189e-06, 9.455106e-07, 9.833365e-07, 
    7.966379e-07, 8.733012e-07, 6.845709e-07, 7.265035e-07, 6.748084e-07, 
    7.008151e-07, 6.56719e-07, 6.963037e-07, 6.288712e-07, 6.148886e-07, 
    6.244167e-07, 5.884427e-07, 6.985509e-07, 6.54508e-07, 1.045658e-06, 
    1.042921e-06, 1.030248e-06, 1.086866e-06, 1.090408e-06, 1.144545e-06, 
    1.096277e-06, 1.076209e-06, 1.026564e-06, 9.980467e-07, 9.715176e-07, 
    9.15126e-07, 8.552013e-07, 7.766076e-07, 7.237256e-07, 6.898854e-07, 
    7.104867e-07, 6.922739e-07, 7.126573e-07, 7.223722e-07, 6.200975e-07, 
    6.760174e-07, 5.935144e-07, 5.97863e-07, 6.343653e-07, 5.973718e-07, 
    1.041003e-06, 1.056805e-06, 1.113118e-06, 1.068855e-06, 1.150566e-06, 
    1.104245e-06, 1.078276e-06, 9.825275e-07, 9.624179e-07, 9.440504e-07, 
    9.085866e-07, 8.646055e-07, 7.91487e-07, 7.318902e-07, 6.806105e-07, 
    6.842698e-07, 6.829796e-07, 6.71886e-07, 6.99624e-07, 6.67416e-07, 
    6.621241e-07, 6.760269e-07, 5.984472e-07, 6.198597e-07, 5.979557e-07, 
    6.118221e-07, 1.051649e-06, 1.025269e-06, 1.039458e-06, 1.0129e-06, 
    1.031552e-06, 9.506155e-07, 9.273436e-07, 8.243044e-07, 8.654534e-07, 
    8.007021e-07, 8.586973e-07, 8.481872e-07, 7.986449e-07, 8.554835e-07, 
    7.350771e-07, 8.151321e-07, 6.714578e-07, 7.459801e-07, 6.669894e-07, 
    6.808261e-07, 6.580395e-07, 6.3814e-07, 6.137821e-07, 5.707476e-07, 
    5.804965e-07, 5.458984e-07, 9.869069e-07, 9.544459e-07, 9.572753e-07, 
    9.241314e-07, 9.002006e-07, 8.500011e-07, 7.7408e-07, 8.019808e-07, 
    7.513521e-07, 7.414953e-07, 8.186545e-07, 7.705689e-07, 9.331958e-07, 
    9.052474e-07, 9.218117e-07, 9.84312e-07, 7.954761e-07, 8.884575e-07, 
    7.228751e-07, 7.687095e-07, 6.409476e-07, 7.022107e-07, 5.859176e-07, 
    5.41065e-07, 5.01369e-07, 4.578929e-07, 9.370913e-07, 9.587428e-07, 
    9.202519e-07, 8.689917e-07, 8.234672e-07, 7.658495e-07, 7.601398e-07, 
    7.497655e-07, 7.234137e-07, 7.01821e-07, 7.46504e-07, 6.964885e-07, 
    8.988496e-07, 7.87782e-07, 9.670244e-07, 9.099999e-07, 8.719522e-07, 
    8.884916e-07, 8.052203e-07, 7.865129e-07, 7.139611e-07, 7.507827e-07, 
    5.518729e-07, 6.33992e-07, 4.268272e-07, 4.783771e-07, 9.663978e-07, 
    9.371678e-07, 8.407765e-07, 8.85621e-07, 7.621211e-07, 7.338979e-07, 
    7.115667e-07, 6.837921e-07, 6.808482e-07, 6.648517e-07, 6.912209e-07, 
    6.658797e-07, 7.657303e-07, 7.197588e-07, 8.513896e-07, 8.177441e-07, 
    8.330923e-07, 8.50182e-07, 7.983023e-07, 7.457826e-07, 7.446982e-07, 
    7.284609e-07, 6.841793e-07, 7.6165e-07, 5.419024e-07, 6.706471e-07, 
    9.06086e-07, 8.531461e-07, 8.457963e-07, 8.658707e-07, 7.366897e-07, 
    7.816182e-07, 6.65239e-07, 6.952562e-07, 6.466128e-07, 6.704387e-07, 
    6.74001e-07, 7.057367e-07, 7.260759e-07, 7.795109e-07, 8.252193e-07, 
    8.629374e-07, 8.540497e-07, 8.130236e-07, 7.426619e-07, 6.805789e-07, 
    6.938163e-07, 6.502133e-07, 7.705938e-07, 7.181595e-07, 7.380809e-07, 
    6.870228e-07, 8.027311e-07, 7.032959e-07, 8.298262e-07, 8.18071e-07, 
    7.825312e-07, 7.147021e-07, 7.003484e-07, 6.852599e-07, 6.945415e-07, 
    7.409413e-07, 7.487722e-07, 7.833823e-07, 7.931513e-07, 8.206198e-07, 
    8.439154e-07, 8.22609e-07, 8.006872e-07, 7.409243e-07, 6.901079e-07, 
    6.378592e-07, 6.255605e-07, 5.693503e-07, 6.147835e-07, 5.412431e-07, 
    6.032818e-07, 4.991481e-07, 6.978553e-07, 6.051999e-07, 7.809459e-07, 
    7.602986e-07, 7.240324e-07, 6.459746e-07, 6.872563e-07, 6.391777e-07, 
    7.490808e-07, 8.116322e-07, 8.284726e-07, 8.60605e-07, 8.277491e-07, 
    8.303845e-07, 7.997947e-07, 8.095274e-07, 7.390019e-07, 7.762599e-07, 
    6.740888e-07, 6.395484e-07, 5.494445e-07, 4.993351e-07, 4.520861e-07, 
    4.323743e-07, 4.265108e-07, 4.240779e-07,
  1.369036e-09, 1.195348e-09, 1.227792e-09, 1.097223e-09, 1.168352e-09, 
    1.084733e-09, 1.332445e-09, 1.188793e-09, 1.279132e-09, 1.352708e-09, 
    8.726922e-10, 1.091644e-09, 6.804559e-10, 7.944799e-10, 5.306861e-10, 
    6.973783e-10, 5.008369e-10, 5.350666e-10, 4.367275e-10, 4.634897e-10, 
    3.522546e-10, 4.247456e-10, 3.025842e-10, 3.687258e-10, 3.577778e-10, 
    4.272973e-10, 1.04475e-09, 8.980622e-10, 1.053942e-09, 1.031909e-09, 
    1.041758e-09, 1.166844e-09, 1.233802e-09, 1.383035e-09, 1.355024e-09, 
    1.245874e-09, 1.02211e-09, 1.094525e-09, 9.18719e-10, 9.224494e-10, 
    7.51005e-10, 8.252098e-10, 5.726633e-10, 6.379162e-10, 4.623507e-10, 
    5.028332e-10, 4.64198e-10, 4.756879e-10, 4.640496e-10, 5.243919e-10, 
    4.97908e-10, 5.533505e-10, 8.109307e-10, 7.279596e-10, 9.949508e-10, 
    1.185548e-09, 1.325891e-09, 1.432499e-09, 1.417063e-09, 1.387968e-09, 
    1.245255e-09, 1.121059e-09, 1.032591e-09, 9.762826e-10, 9.229865e-10, 
    7.742618e-10, 7.028846e-10, 5.600574e-10, 5.841755e-10, 5.437404e-10, 
    5.069912e-10, 4.492309e-10, 4.58407e-10, 4.341338e-10, 5.447879e-10, 
    4.693068e-10, 5.982317e-10, 5.607818e-10, 9.088133e-10, 1.07464e-09, 
    1.151244e-09, 1.221505e-09, 1.405276e-09, 1.27638e-09, 1.326119e-09, 
    1.210032e-09, 1.140188e-09, 1.17436e-09, 9.747746e-10, 1.049206e-09, 
    6.98806e-10, 8.373984e-10, 5.111854e-10, 5.791679e-10, 4.957617e-10, 
    5.371916e-10, 4.675994e-10, 5.299268e-10, 4.253348e-10, 4.046284e-10, 
    4.187004e-10, 3.664418e-10, 5.335415e-10, 4.641951e-10, 1.175326e-09, 
    1.169699e-09, 1.143748e-09, 1.260995e-09, 1.268442e-09, 1.383805e-09, 
    1.280806e-09, 1.238672e-09, 1.136236e-09, 1.078591e-09, 1.025774e-09, 
    9.161965e-10, 8.039798e-10, 6.639112e-10, 5.745794e-10, 5.19647e-10, 
    5.528748e-10, 5.234648e-10, 5.564147e-10, 5.72348e-10, 4.123012e-10, 
    4.976636e-10, 3.73664e-10, 3.79895e-10, 4.335665e-10, 3.791894e-10, 
    1.165761e-09, 1.198326e-09, 1.316481e-09, 1.223334e-09, 1.396813e-09, 
    1.29765e-09, 1.242994e-09, 1.047598e-09, 1.00784e-09, 9.719348e-10, 
    9.03734e-10, 8.212903e-10, 6.897785e-10, 5.880995e-10, 5.049096e-10, 
    5.107074e-10, 5.086607e-10, 4.911752e-10, 5.352704e-10, 4.841869e-10, 
    4.759571e-10, 4.976783e-10, 3.807347e-10, 4.119495e-10, 3.800282e-10, 
    4.001341e-10, 1.187671e-09, 1.133599e-09, 1.162591e-09, 1.108504e-09, 
    1.146411e-09, 9.847241e-10, 9.396193e-10, 7.479185e-10, 8.228568e-10, 
    7.059545e-10, 8.104013e-10, 7.911424e-10, 7.023341e-10, 8.044968e-10, 
    5.934046e-10, 7.315208e-10, 4.905041e-10, 6.11669e-10, 4.835217e-10, 
    5.052505e-10, 4.696364e-10, 4.392525e-10, 4.030046e-10, 3.416296e-10, 
    3.55225e-10, 3.078267e-10, 1.056316e-09, 9.922086e-10, 9.97748e-10, 
    9.334431e-10, 8.87829e-10, 7.944557e-10, 6.59548e-10, 7.082078e-10, 
    6.207319e-10, 6.041339e-10, 7.378034e-10, 6.53503e-10, 9.509011e-10, 
    8.973913e-10, 9.289913e-10, 1.051148e-09, 6.967664e-10, 8.657026e-10, 
    5.73177e-10, 6.503083e-10, 4.434979e-10, 5.394462e-10, 3.628645e-10, 
    3.013977e-10, 2.504669e-10, 1.987598e-10, 9.584334e-10, 1.000625e-09, 
    9.260012e-10, 8.294038e-10, 7.464164e-10, 6.454048e-10, 6.356508e-10, 
    6.180506e-10, 5.740648e-10, 5.388159e-10, 6.125506e-10, 5.302237e-10, 
    8.852764e-10, 6.833081e-10, 1.016907e-09, 9.06424e-10, 8.348933e-10, 
    8.65766e-10, 7.139279e-10, 6.81096e-10, 5.58545e-10, 6.197691e-10, 
    3.158409e-10, 4.330059e-10, 1.646426e-10, 2.225683e-10, 1.015672e-09, 
    9.585813e-10, 7.776496e-10, 8.60383e-10, 6.390302e-10, 5.914393e-10, 
    5.546352e-10, 5.099495e-10, 5.052855e-10, 4.801931e-10, 5.217805e-10, 
    4.817928e-10, 6.452008e-10, 5.680476e-10, 7.96995e-10, 7.361779e-10, 
    7.637344e-10, 7.947863e-10, 7.0173e-10, 6.113361e-10, 6.095114e-10, 
    5.824084e-10, 5.105658e-10, 6.382261e-10, 3.02509e-10, 4.892367e-10, 
    8.989821e-10, 8.00212e-10, 7.867812e-10, 8.236278e-10, 5.960941e-10, 
    6.725865e-10, 4.807955e-10, 5.282444e-10, 4.52106e-10, 4.889088e-10, 
    4.944931e-10, 5.45154e-10, 5.784609e-10, 6.689336e-10, 7.495597e-10, 
    8.182111e-10, 8.018671e-10, 7.277666e-10, 6.060911e-10, 5.048599e-10, 
    5.259354e-10, 4.576057e-10, 6.535454e-10, 5.654213e-10, 5.984181e-10, 
    5.150836e-10, 7.095314e-10, 5.412023e-10, 7.578439e-10, 7.367613e-10, 
    6.741713e-10, 5.597571e-10, 5.364387e-10, 5.122801e-10, 5.270976e-10, 
    6.032055e-10, 6.163736e-10, 6.756495e-10, 6.92691e-10, 7.413166e-10, 
    7.833554e-10, 7.448782e-10, 7.05928e-10, 6.031768e-10, 5.200025e-10, 
    4.388288e-10, 4.204004e-10, 3.396969e-10, 4.044747e-10, 3.016347e-10, 
    3.877109e-10, 2.477205e-10, 5.324228e-10, 3.904888e-10, 6.714202e-10, 
    6.359215e-10, 5.750861e-10, 4.511343e-10, 5.154553e-10, 4.408204e-10, 
    6.168945e-10, 7.252933e-10, 7.554068e-10, 8.139122e-10, 7.541053e-10, 
    7.588498e-10, 7.043559e-10, 7.215558e-10, 5.999581e-10, 6.6331e-10, 
    4.946312e-10, 4.413808e-10, 3.125744e-10, 2.479507e-10, 1.921962e-10, 
    1.705521e-10, 1.643077e-10, 1.617435e-10,
  4.068486e-13, 4.060852e-13, 4.062279e-13, 4.056536e-13, 4.059665e-13, 
    4.055986e-13, 4.066878e-13, 4.060564e-13, 4.064536e-13, 4.067769e-13, 
    4.046646e-13, 4.05629e-13, 4.038162e-13, 4.043196e-13, 4.03154e-13, 
    4.038909e-13, 4.030219e-13, 4.031733e-13, 4.027379e-13, 4.028565e-13, 
    4.023634e-13, 4.026848e-13, 4.021429e-13, 4.024364e-13, 4.023879e-13, 
    4.026961e-13, 4.054226e-13, 4.047764e-13, 4.054631e-13, 4.053661e-13, 
    4.054094e-13, 4.059599e-13, 4.062543e-13, 4.069101e-13, 4.06787e-13, 
    4.063074e-13, 4.053229e-13, 4.056417e-13, 4.048674e-13, 4.048839e-13, 
    4.041277e-13, 4.044551e-13, 4.033397e-13, 4.036282e-13, 4.028514e-13, 
    4.030307e-13, 4.028596e-13, 4.029105e-13, 4.02859e-13, 4.031261e-13, 
    4.030089e-13, 4.032543e-13, 4.043922e-13, 4.04026e-13, 4.052033e-13, 
    4.060421e-13, 4.06659e-13, 4.071273e-13, 4.070595e-13, 4.069317e-13, 
    4.063047e-13, 4.057585e-13, 4.053691e-13, 4.051211e-13, 4.048862e-13, 
    4.042304e-13, 4.039152e-13, 4.032839e-13, 4.033906e-13, 4.032117e-13, 
    4.030491e-13, 4.027933e-13, 4.02834e-13, 4.027264e-13, 4.032164e-13, 
    4.028822e-13, 4.034528e-13, 4.032871e-13, 4.048238e-13, 4.055542e-13, 
    4.058912e-13, 4.062002e-13, 4.070077e-13, 4.064415e-13, 4.066601e-13, 
    4.061498e-13, 4.058426e-13, 4.059929e-13, 4.051144e-13, 4.054422e-13, 
    4.038972e-13, 4.045089e-13, 4.030677e-13, 4.033685e-13, 4.029994e-13, 
    4.031827e-13, 4.028747e-13, 4.031506e-13, 4.026874e-13, 4.025957e-13, 
    4.02658e-13, 4.024263e-13, 4.031666e-13, 4.028596e-13, 4.059972e-13, 
    4.059724e-13, 4.058583e-13, 4.063739e-13, 4.064066e-13, 4.069134e-13, 
    4.064609e-13, 4.062757e-13, 4.058252e-13, 4.055716e-13, 4.05339e-13, 
    4.048563e-13, 4.043615e-13, 4.037431e-13, 4.033482e-13, 4.031051e-13, 
    4.032521e-13, 4.03122e-13, 4.032678e-13, 4.033383e-13, 4.026297e-13, 
    4.030078e-13, 4.024583e-13, 4.02486e-13, 4.027239e-13, 4.024828e-13, 
    4.059551e-13, 4.060983e-13, 4.066177e-13, 4.062083e-13, 4.069706e-13, 
    4.065349e-13, 4.062947e-13, 4.054351e-13, 4.052601e-13, 4.051019e-13, 
    4.048014e-13, 4.044378e-13, 4.038573e-13, 4.03408e-13, 4.030399e-13, 
    4.030655e-13, 4.030565e-13, 4.029791e-13, 4.031743e-13, 4.029481e-13, 
    4.029117e-13, 4.030079e-13, 4.024897e-13, 4.026281e-13, 4.024866e-13, 
    4.025757e-13, 4.060515e-13, 4.058136e-13, 4.059411e-13, 4.057032e-13, 
    4.0587e-13, 4.051582e-13, 4.049595e-13, 4.041141e-13, 4.044448e-13, 
    4.039288e-13, 4.043898e-13, 4.043048e-13, 4.039128e-13, 4.043638e-13, 
    4.034314e-13, 4.040417e-13, 4.029761e-13, 4.035122e-13, 4.029452e-13, 
    4.030414e-13, 4.028837e-13, 4.027491e-13, 4.025884e-13, 4.023162e-13, 
    4.023765e-13, 4.021661e-13, 4.054735e-13, 4.051912e-13, 4.052156e-13, 
    4.049323e-13, 4.047313e-13, 4.043195e-13, 4.037238e-13, 4.039387e-13, 
    4.035522e-13, 4.034789e-13, 4.040694e-13, 4.036971e-13, 4.050093e-13, 
    4.047734e-13, 4.049127e-13, 4.054508e-13, 4.038882e-13, 4.046337e-13, 
    4.03342e-13, 4.03683e-13, 4.027679e-13, 4.031927e-13, 4.024104e-13, 
    4.021376e-13, 4.019113e-13, 4.016812e-13, 4.050425e-13, 4.052283e-13, 
    4.048995e-13, 4.044737e-13, 4.041075e-13, 4.036613e-13, 4.036182e-13, 
    4.035404e-13, 4.033459e-13, 4.031899e-13, 4.035161e-13, 4.031519e-13, 
    4.0472e-13, 4.038288e-13, 4.053e-13, 4.048133e-13, 4.044979e-13, 
    4.04634e-13, 4.03964e-13, 4.03819e-13, 4.032772e-13, 4.03548e-13, 
    4.022017e-13, 4.027214e-13, 4.015293e-13, 4.017872e-13, 4.052946e-13, 
    4.050431e-13, 4.042453e-13, 4.046103e-13, 4.036331e-13, 4.034227e-13, 
    4.032599e-13, 4.030622e-13, 4.030415e-13, 4.029305e-13, 4.031146e-13, 
    4.029375e-13, 4.036604e-13, 4.033193e-13, 4.043307e-13, 4.040623e-13, 
    4.041839e-13, 4.043209e-13, 4.039101e-13, 4.035107e-13, 4.035026e-13, 
    4.033828e-13, 4.030649e-13, 4.036296e-13, 4.021425e-13, 4.029705e-13, 
    4.047805e-13, 4.043449e-13, 4.042856e-13, 4.044482e-13, 4.034433e-13, 
    4.037814e-13, 4.029331e-13, 4.031431e-13, 4.02806e-13, 4.029691e-13, 
    4.029938e-13, 4.03218e-13, 4.033653e-13, 4.037653e-13, 4.041213e-13, 
    4.044243e-13, 4.043522e-13, 4.040251e-13, 4.034875e-13, 4.030397e-13, 
    4.031329e-13, 4.028304e-13, 4.036973e-13, 4.033076e-13, 4.034536e-13, 
    4.030849e-13, 4.039446e-13, 4.032005e-13, 4.041579e-13, 4.040648e-13, 
    4.037884e-13, 4.032826e-13, 4.031794e-13, 4.030725e-13, 4.031381e-13, 
    4.034748e-13, 4.03533e-13, 4.037949e-13, 4.038702e-13, 4.040849e-13, 
    4.042705e-13, 4.041007e-13, 4.039287e-13, 4.034746e-13, 4.031067e-13, 
    4.027472e-13, 4.026656e-13, 4.023076e-13, 4.02595e-13, 4.021386e-13, 
    4.025206e-13, 4.018991e-13, 4.031617e-13, 4.02533e-13, 4.037762e-13, 
    4.036194e-13, 4.033504e-13, 4.028017e-13, 4.030866e-13, 4.027561e-13, 
    4.035353e-13, 4.040142e-13, 4.041471e-13, 4.044053e-13, 4.041414e-13, 
    4.041623e-13, 4.039217e-13, 4.039977e-13, 4.034604e-13, 4.037404e-13, 
    4.029944e-13, 4.027585e-13, 4.021872e-13, 4.019001e-13, 4.01652e-13, 
    4.015556e-13, 4.015278e-13, 4.015164e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC =
  8.94965e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 
    8.94965e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 
    8.949648e-07, 8.94965e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 
    8.949648e-07, 8.949647e-07, 8.949647e-07, 8.949646e-07, 8.949647e-07, 
    8.949646e-07, 8.949646e-07, 8.949646e-07, 8.949646e-07, 8.949646e-07, 
    8.949646e-07, 8.94965e-07, 8.949649e-07, 8.94965e-07, 8.949649e-07, 
    8.94965e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 
    8.94965e-07, 8.949649e-07, 8.94965e-07, 8.949649e-07, 8.949649e-07, 
    8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949648e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949648e-07, 8.949648e-07, 8.949649e-07, 
    8.94965e-07, 8.94965e-07, 8.949651e-07, 8.949651e-07, 8.949651e-07, 
    8.94965e-07, 8.94965e-07, 8.949649e-07, 8.949649e-07, 8.949649e-07, 
    8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949646e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949649e-07, 8.94965e-07, 
    8.94965e-07, 8.94965e-07, 8.949651e-07, 8.94965e-07, 8.94965e-07, 
    8.94965e-07, 8.94965e-07, 8.94965e-07, 8.949649e-07, 8.94965e-07, 
    8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949646e-07, 8.949646e-07, 
    8.949646e-07, 8.949646e-07, 8.949647e-07, 8.949647e-07, 8.94965e-07, 
    8.94965e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 8.949651e-07, 
    8.94965e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 8.949649e-07, 
    8.949649e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949646e-07, 
    8.949647e-07, 8.949646e-07, 8.949646e-07, 8.949646e-07, 8.949646e-07, 
    8.94965e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 8.949651e-07, 
    8.94965e-07, 8.94965e-07, 8.94965e-07, 8.949649e-07, 8.949649e-07, 
    8.949649e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949646e-07, 8.949646e-07, 8.949646e-07, 
    8.949646e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 8.94965e-07, 
    8.94965e-07, 8.949649e-07, 8.949649e-07, 8.949648e-07, 8.949648e-07, 
    8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949648e-07, 
    8.949647e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949646e-07, 8.949646e-07, 8.949646e-07, 
    8.949646e-07, 8.949646e-07, 8.94965e-07, 8.949649e-07, 8.949649e-07, 
    8.949649e-07, 8.949649e-07, 8.949648e-07, 8.949648e-07, 8.949648e-07, 
    8.949647e-07, 8.949647e-07, 8.949648e-07, 8.949648e-07, 8.949649e-07, 
    8.949649e-07, 8.949649e-07, 8.94965e-07, 8.949648e-07, 8.949648e-07, 
    8.949647e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 8.949646e-07, 
    8.949646e-07, 8.949645e-07, 8.949644e-07, 8.949649e-07, 8.949649e-07, 
    8.949649e-07, 8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949648e-07, 8.949648e-07, 8.949649e-07, 8.949649e-07, 8.949648e-07, 
    8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 
    8.949646e-07, 8.949646e-07, 8.949644e-07, 8.949644e-07, 8.949649e-07, 
    8.949649e-07, 8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949648e-07, 8.949647e-07, 8.949648e-07, 8.949648e-07, 
    8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949648e-07, 8.949646e-07, 8.949647e-07, 
    8.949649e-07, 8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 
    8.949648e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949648e-07, 8.949648e-07, 
    8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949648e-07, 8.949647e-07, 8.949648e-07, 8.949648e-07, 
    8.949648e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949647e-07, 8.949648e-07, 8.949648e-07, 8.949648e-07, 
    8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949647e-07, 
    8.949646e-07, 8.949646e-07, 8.949646e-07, 8.949646e-07, 8.949646e-07, 
    8.949646e-07, 8.949645e-07, 8.949647e-07, 8.949646e-07, 8.949648e-07, 
    8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 8.949647e-07, 
    8.949647e-07, 8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949648e-07, 
    8.949648e-07, 8.949648e-07, 8.949648e-07, 8.949647e-07, 8.949648e-07, 
    8.949647e-07, 8.949647e-07, 8.949646e-07, 8.949645e-07, 8.949644e-07, 
    8.949644e-07, 8.949644e-07, 8.949644e-07 ;

 CWDC_HR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC_LOSS =
  6.969069e-16, 6.986815e-16, 6.983368e-16, 6.997667e-16, 6.989739e-16, 
    6.999098e-16, 6.97267e-16, 6.987517e-16, 6.978043e-16, 6.970671e-16, 
    7.025372e-16, 6.998306e-16, 7.053463e-16, 7.036234e-16, 7.079484e-16, 
    7.050779e-16, 7.085266e-16, 7.078663e-16, 7.098544e-16, 7.092851e-16, 
    7.118236e-16, 7.10117e-16, 7.131388e-16, 7.114166e-16, 7.116859e-16, 
    7.100606e-16, 7.003763e-16, 7.022003e-16, 7.00268e-16, 7.005283e-16, 
    7.004116e-16, 6.989901e-16, 6.982728e-16, 6.967716e-16, 6.970444e-16, 
    6.981472e-16, 7.006453e-16, 6.997982e-16, 7.019336e-16, 7.018854e-16, 
    7.042588e-16, 7.031891e-16, 7.071732e-16, 7.060421e-16, 7.093089e-16, 
    7.08488e-16, 7.092702e-16, 7.090332e-16, 7.092733e-16, 7.080691e-16, 
    7.085851e-16, 7.075253e-16, 7.033894e-16, 7.046059e-16, 7.009745e-16, 
    6.987859e-16, 6.973321e-16, 6.962992e-16, 6.964453e-16, 6.967236e-16, 
    6.981536e-16, 6.994975e-16, 7.005208e-16, 7.012047e-16, 7.018784e-16, 
    7.039143e-16, 7.049921e-16, 7.074015e-16, 7.069676e-16, 7.077031e-16, 
    7.084063e-16, 7.095853e-16, 7.093914e-16, 7.099104e-16, 7.076841e-16, 
    7.091639e-16, 7.067201e-16, 7.073889e-16, 7.020594e-16, 7.000269e-16, 
    6.991603e-16, 6.98403e-16, 6.965575e-16, 6.978321e-16, 6.973297e-16, 
    6.985251e-16, 6.992839e-16, 6.989087e-16, 7.012234e-16, 7.003239e-16, 
    7.050559e-16, 7.030195e-16, 7.083243e-16, 7.070567e-16, 7.08628e-16, 
    7.078265e-16, 7.091994e-16, 7.079639e-16, 7.101038e-16, 7.105691e-16, 
    7.10251e-16, 7.114729e-16, 7.078953e-16, 7.0927e-16, 6.988981e-16, 
    6.989593e-16, 6.992445e-16, 6.979902e-16, 6.979136e-16, 6.96764e-16, 
    6.977872e-16, 6.982225e-16, 6.99328e-16, 6.999811e-16, 7.006019e-16, 
    7.019659e-16, 7.034875e-16, 7.056132e-16, 7.071388e-16, 7.081606e-16, 
    7.075343e-16, 7.080872e-16, 7.07469e-16, 7.071793e-16, 7.103946e-16, 
    7.085899e-16, 7.112972e-16, 7.111476e-16, 7.099227e-16, 7.111645e-16, 
    6.990023e-16, 6.986501e-16, 6.974262e-16, 6.983841e-16, 6.966388e-16, 
    6.976157e-16, 6.98177e-16, 7.003422e-16, 7.00818e-16, 7.012584e-16, 
    7.021284e-16, 7.032439e-16, 7.051986e-16, 7.068976e-16, 7.084472e-16, 
    7.083338e-16, 7.083737e-16, 7.087195e-16, 7.078626e-16, 7.088601e-16, 
    7.090272e-16, 7.085899e-16, 7.111276e-16, 7.104031e-16, 7.111445e-16, 
    7.106728e-16, 6.987646e-16, 6.993572e-16, 6.99037e-16, 6.996389e-16, 
    6.992147e-16, 7.010995e-16, 7.016642e-16, 7.043042e-16, 7.032218e-16, 
    7.049447e-16, 7.033971e-16, 7.036713e-16, 7.049999e-16, 7.034809e-16, 
    7.068036e-16, 7.045509e-16, 7.087329e-16, 7.064854e-16, 7.088736e-16, 
    7.084406e-16, 7.091576e-16, 7.097994e-16, 7.106067e-16, 7.120945e-16, 
    7.117502e-16, 7.129938e-16, 7.002403e-16, 7.01008e-16, 7.009408e-16, 
    7.01744e-16, 7.023376e-16, 7.036241e-16, 7.056846e-16, 7.049102e-16, 
    7.06332e-16, 7.066171e-16, 7.044572e-16, 7.057834e-16, 7.015218e-16, 
    7.022107e-16, 7.018008e-16, 7.003007e-16, 7.050882e-16, 7.026328e-16, 
    7.07164e-16, 7.058363e-16, 7.097078e-16, 7.077833e-16, 7.115605e-16, 
    7.131711e-16, 7.146872e-16, 7.164546e-16, 7.014271e-16, 7.009057e-16, 
    7.018396e-16, 7.0313e-16, 7.043274e-16, 7.059173e-16, 7.0608e-16, 
    7.063775e-16, 7.071484e-16, 7.077959e-16, 7.064712e-16, 7.079582e-16, 
    7.023696e-16, 7.053013e-16, 7.007082e-16, 7.020922e-16, 7.030541e-16, 
    7.026326e-16, 7.048218e-16, 7.053371e-16, 7.074294e-16, 7.063485e-16, 
    7.127734e-16, 7.099343e-16, 7.178002e-16, 7.156062e-16, 7.007234e-16, 
    7.014255e-16, 7.038662e-16, 7.027055e-16, 7.060235e-16, 7.068389e-16, 
    7.075018e-16, 7.083481e-16, 7.084398e-16, 7.08941e-16, 7.081195e-16, 
    7.089087e-16, 7.059206e-16, 7.072567e-16, 7.035879e-16, 7.044815e-16, 
    7.040706e-16, 7.036195e-16, 7.050113e-16, 7.064919e-16, 7.065242e-16, 
    7.069985e-16, 7.083333e-16, 7.06037e-16, 7.131382e-16, 7.087557e-16, 
    7.021908e-16, 7.035408e-16, 7.037343e-16, 7.032114e-16, 7.067572e-16, 
    7.054733e-16, 7.089288e-16, 7.079959e-16, 7.095244e-16, 7.08765e-16, 
    7.086532e-16, 7.076773e-16, 7.070693e-16, 7.055321e-16, 7.042804e-16, 
    7.032873e-16, 7.035184e-16, 7.04609e-16, 7.065826e-16, 7.084478e-16, 
    7.080393e-16, 7.094083e-16, 7.057832e-16, 7.07304e-16, 7.067162e-16, 
    7.082486e-16, 7.048895e-16, 7.077484e-16, 7.041577e-16, 7.04473e-16, 
    7.054478e-16, 7.074067e-16, 7.078407e-16, 7.083027e-16, 7.080177e-16, 
    7.066328e-16, 7.064061e-16, 7.054243e-16, 7.051528e-16, 7.044044e-16, 
    7.037841e-16, 7.043507e-16, 7.049452e-16, 7.066337e-16, 7.081533e-16, 
    7.098084e-16, 7.102135e-16, 7.121427e-16, 7.105715e-16, 7.131625e-16, 
    7.109586e-16, 7.147721e-16, 7.079149e-16, 7.108951e-16, 7.054924e-16, 
    7.060755e-16, 7.07129e-16, 7.095438e-16, 7.082414e-16, 7.097648e-16, 
    7.063973e-16, 7.046463e-16, 7.041937e-16, 7.033476e-16, 7.04213e-16, 
    7.041427e-16, 7.049703e-16, 7.047045e-16, 7.066897e-16, 7.056237e-16, 
    7.086502e-16, 7.097529e-16, 7.128634e-16, 7.147663e-16, 7.167018e-16, 
    7.175551e-16, 7.178147e-16, 7.179232e-16 ;

 CWDC_TO_LITR2C =
  5.296492e-16, 5.30998e-16, 5.30736e-16, 5.318227e-16, 5.312202e-16, 
    5.319315e-16, 5.29923e-16, 5.310513e-16, 5.303312e-16, 5.29771e-16, 
    5.339283e-16, 5.318713e-16, 5.360632e-16, 5.347538e-16, 5.380408e-16, 
    5.358592e-16, 5.384802e-16, 5.379784e-16, 5.394893e-16, 5.390567e-16, 
    5.40986e-16, 5.396889e-16, 5.419855e-16, 5.406766e-16, 5.408813e-16, 
    5.39646e-16, 5.32286e-16, 5.336722e-16, 5.322037e-16, 5.324015e-16, 
    5.323128e-16, 5.312325e-16, 5.306874e-16, 5.295464e-16, 5.297537e-16, 
    5.305919e-16, 5.324904e-16, 5.318466e-16, 5.334695e-16, 5.334329e-16, 
    5.352367e-16, 5.344237e-16, 5.374517e-16, 5.36592e-16, 5.390747e-16, 
    5.384509e-16, 5.390454e-16, 5.388652e-16, 5.390477e-16, 5.381325e-16, 
    5.385247e-16, 5.377192e-16, 5.345759e-16, 5.355005e-16, 5.327406e-16, 
    5.310773e-16, 5.299724e-16, 5.291874e-16, 5.292984e-16, 5.295099e-16, 
    5.305967e-16, 5.316181e-16, 5.323958e-16, 5.329156e-16, 5.334276e-16, 
    5.349748e-16, 5.35794e-16, 5.376252e-16, 5.372953e-16, 5.378544e-16, 
    5.383888e-16, 5.392848e-16, 5.391374e-16, 5.395319e-16, 5.378399e-16, 
    5.389646e-16, 5.371073e-16, 5.376156e-16, 5.335651e-16, 5.320204e-16, 
    5.313618e-16, 5.307863e-16, 5.293837e-16, 5.303524e-16, 5.299706e-16, 
    5.308791e-16, 5.314557e-16, 5.311707e-16, 5.329298e-16, 5.322461e-16, 
    5.358425e-16, 5.342948e-16, 5.383264e-16, 5.373631e-16, 5.385573e-16, 
    5.379481e-16, 5.389915e-16, 5.380525e-16, 5.396788e-16, 5.400325e-16, 
    5.397908e-16, 5.407194e-16, 5.380004e-16, 5.390452e-16, 5.311626e-16, 
    5.31209e-16, 5.314258e-16, 5.304726e-16, 5.304144e-16, 5.295406e-16, 
    5.303183e-16, 5.306491e-16, 5.314893e-16, 5.319857e-16, 5.324575e-16, 
    5.334941e-16, 5.346505e-16, 5.36266e-16, 5.374255e-16, 5.38202e-16, 
    5.377261e-16, 5.381463e-16, 5.376765e-16, 5.374563e-16, 5.398999e-16, 
    5.385283e-16, 5.405859e-16, 5.404722e-16, 5.395412e-16, 5.40485e-16, 
    5.312418e-16, 5.309741e-16, 5.300439e-16, 5.307719e-16, 5.294455e-16, 
    5.301879e-16, 5.306145e-16, 5.3226e-16, 5.326217e-16, 5.329564e-16, 
    5.336176e-16, 5.344653e-16, 5.359509e-16, 5.372422e-16, 5.384199e-16, 
    5.383337e-16, 5.38364e-16, 5.386268e-16, 5.379756e-16, 5.387337e-16, 
    5.388607e-16, 5.385283e-16, 5.404569e-16, 5.399063e-16, 5.404698e-16, 
    5.401114e-16, 5.310612e-16, 5.315115e-16, 5.312681e-16, 5.317256e-16, 
    5.314032e-16, 5.328357e-16, 5.332648e-16, 5.352712e-16, 5.344486e-16, 
    5.357579e-16, 5.345818e-16, 5.347902e-16, 5.357999e-16, 5.346455e-16, 
    5.371707e-16, 5.354587e-16, 5.38637e-16, 5.369289e-16, 5.387439e-16, 
    5.384148e-16, 5.389598e-16, 5.394475e-16, 5.400611e-16, 5.411918e-16, 
    5.409301e-16, 5.418754e-16, 5.321826e-16, 5.32766e-16, 5.32715e-16, 
    5.333255e-16, 5.337766e-16, 5.347543e-16, 5.363203e-16, 5.357318e-16, 
    5.368123e-16, 5.37029e-16, 5.353875e-16, 5.363954e-16, 5.331565e-16, 
    5.336801e-16, 5.333687e-16, 5.322285e-16, 5.35867e-16, 5.34001e-16, 
    5.374446e-16, 5.364356e-16, 5.39378e-16, 5.379153e-16, 5.40786e-16, 
    5.420101e-16, 5.431623e-16, 5.445055e-16, 5.330846e-16, 5.326884e-16, 
    5.333981e-16, 5.343788e-16, 5.352888e-16, 5.364971e-16, 5.366208e-16, 
    5.368469e-16, 5.374328e-16, 5.379249e-16, 5.369181e-16, 5.380483e-16, 
    5.338009e-16, 5.36029e-16, 5.325382e-16, 5.3359e-16, 5.343211e-16, 
    5.340008e-16, 5.356646e-16, 5.360562e-16, 5.376463e-16, 5.368248e-16, 
    5.417078e-16, 5.395501e-16, 5.455281e-16, 5.438607e-16, 5.325498e-16, 
    5.330834e-16, 5.349383e-16, 5.340562e-16, 5.365779e-16, 5.371976e-16, 
    5.377014e-16, 5.383446e-16, 5.384142e-16, 5.387951e-16, 5.381709e-16, 
    5.387706e-16, 5.364997e-16, 5.375151e-16, 5.347268e-16, 5.354059e-16, 
    5.350936e-16, 5.347508e-16, 5.358086e-16, 5.369339e-16, 5.369584e-16, 
    5.373189e-16, 5.383333e-16, 5.365881e-16, 5.41985e-16, 5.386543e-16, 
    5.33665e-16, 5.34691e-16, 5.348381e-16, 5.344407e-16, 5.371355e-16, 
    5.361597e-16, 5.387859e-16, 5.380769e-16, 5.392385e-16, 5.386614e-16, 
    5.385764e-16, 5.378348e-16, 5.373727e-16, 5.362044e-16, 5.352531e-16, 
    5.344984e-16, 5.34674e-16, 5.355028e-16, 5.370028e-16, 5.384203e-16, 
    5.381099e-16, 5.391503e-16, 5.363952e-16, 5.37551e-16, 5.371043e-16, 
    5.382689e-16, 5.35716e-16, 5.378888e-16, 5.351598e-16, 5.353994e-16, 
    5.361404e-16, 5.376291e-16, 5.379589e-16, 5.383101e-16, 5.380935e-16, 
    5.37041e-16, 5.368686e-16, 5.361225e-16, 5.359161e-16, 5.353473e-16, 
    5.348759e-16, 5.353065e-16, 5.357584e-16, 5.370416e-16, 5.381965e-16, 
    5.394544e-16, 5.397622e-16, 5.412285e-16, 5.400343e-16, 5.420035e-16, 
    5.403285e-16, 5.432268e-16, 5.380153e-16, 5.402802e-16, 5.361742e-16, 
    5.366174e-16, 5.374181e-16, 5.392533e-16, 5.382634e-16, 5.394212e-16, 
    5.368619e-16, 5.355312e-16, 5.351872e-16, 5.345442e-16, 5.352019e-16, 
    5.351484e-16, 5.357775e-16, 5.355754e-16, 5.370842e-16, 5.36274e-16, 
    5.385741e-16, 5.394122e-16, 5.417761e-16, 5.432224e-16, 5.446934e-16, 
    5.453418e-16, 5.455392e-16, 5.456216e-16 ;

 CWDC_TO_LITR3C =
  1.672577e-16, 1.676836e-16, 1.676008e-16, 1.67944e-16, 1.677538e-16, 
    1.679784e-16, 1.673441e-16, 1.677004e-16, 1.67473e-16, 1.672961e-16, 
    1.686089e-16, 1.679593e-16, 1.692831e-16, 1.688696e-16, 1.699076e-16, 
    1.692187e-16, 1.700464e-16, 1.698879e-16, 1.70365e-16, 1.702284e-16, 
    1.708377e-16, 1.704281e-16, 1.711533e-16, 1.7074e-16, 1.708046e-16, 
    1.704145e-16, 1.680903e-16, 1.685281e-16, 1.680643e-16, 1.681268e-16, 
    1.680988e-16, 1.677576e-16, 1.675855e-16, 1.672252e-16, 1.672906e-16, 
    1.675553e-16, 1.681549e-16, 1.679516e-16, 1.684641e-16, 1.684525e-16, 
    1.690221e-16, 1.687654e-16, 1.697216e-16, 1.694501e-16, 1.702341e-16, 
    1.700371e-16, 1.702249e-16, 1.70168e-16, 1.702256e-16, 1.699366e-16, 
    1.700604e-16, 1.698061e-16, 1.688135e-16, 1.691054e-16, 1.682339e-16, 
    1.677086e-16, 1.673597e-16, 1.671118e-16, 1.671469e-16, 1.672137e-16, 
    1.675569e-16, 1.678794e-16, 1.68125e-16, 1.682891e-16, 1.684508e-16, 
    1.689394e-16, 1.691981e-16, 1.697764e-16, 1.696722e-16, 1.698487e-16, 
    1.700175e-16, 1.703005e-16, 1.702539e-16, 1.703785e-16, 1.698442e-16, 
    1.701993e-16, 1.696128e-16, 1.697733e-16, 1.684943e-16, 1.680064e-16, 
    1.677985e-16, 1.676167e-16, 1.671738e-16, 1.674797e-16, 1.673591e-16, 
    1.67646e-16, 1.678281e-16, 1.677381e-16, 1.682936e-16, 1.680777e-16, 
    1.692134e-16, 1.687247e-16, 1.699978e-16, 1.696936e-16, 1.700707e-16, 
    1.698784e-16, 1.702079e-16, 1.699113e-16, 1.704249e-16, 1.705366e-16, 
    1.704603e-16, 1.707535e-16, 1.698949e-16, 1.702248e-16, 1.677356e-16, 
    1.677502e-16, 1.678187e-16, 1.675177e-16, 1.674993e-16, 1.672234e-16, 
    1.674689e-16, 1.675734e-16, 1.678387e-16, 1.679955e-16, 1.681445e-16, 
    1.684718e-16, 1.68837e-16, 1.693472e-16, 1.697133e-16, 1.699585e-16, 
    1.698082e-16, 1.699409e-16, 1.697926e-16, 1.69723e-16, 1.704947e-16, 
    1.700616e-16, 1.707113e-16, 1.706754e-16, 1.703814e-16, 1.706795e-16, 
    1.677606e-16, 1.67676e-16, 1.673823e-16, 1.676122e-16, 1.671933e-16, 
    1.674278e-16, 1.675625e-16, 1.680821e-16, 1.681963e-16, 1.68302e-16, 
    1.685108e-16, 1.687785e-16, 1.692477e-16, 1.696554e-16, 1.700273e-16, 
    1.700001e-16, 1.700097e-16, 1.700927e-16, 1.69887e-16, 1.701264e-16, 
    1.701665e-16, 1.700616e-16, 1.706706e-16, 1.704967e-16, 1.706747e-16, 
    1.705615e-16, 1.677035e-16, 1.678457e-16, 1.677689e-16, 1.679133e-16, 
    1.678115e-16, 1.682639e-16, 1.683994e-16, 1.69033e-16, 1.687732e-16, 
    1.691867e-16, 1.688153e-16, 1.688811e-16, 1.692e-16, 1.688354e-16, 
    1.696329e-16, 1.690922e-16, 1.700959e-16, 1.695565e-16, 1.701297e-16, 
    1.700257e-16, 1.701978e-16, 1.703519e-16, 1.705456e-16, 1.709027e-16, 
    1.7082e-16, 1.711185e-16, 1.680577e-16, 1.682419e-16, 1.682258e-16, 
    1.684186e-16, 1.68561e-16, 1.688698e-16, 1.693643e-16, 1.691785e-16, 
    1.695197e-16, 1.695881e-16, 1.690697e-16, 1.69388e-16, 1.683652e-16, 
    1.685306e-16, 1.684322e-16, 1.680722e-16, 1.692212e-16, 1.686319e-16, 
    1.697194e-16, 1.694007e-16, 1.703299e-16, 1.69868e-16, 1.707745e-16, 
    1.711611e-16, 1.715249e-16, 1.719491e-16, 1.683425e-16, 1.682174e-16, 
    1.684415e-16, 1.687512e-16, 1.690386e-16, 1.694201e-16, 1.694592e-16, 
    1.695306e-16, 1.697156e-16, 1.69871e-16, 1.695531e-16, 1.6991e-16, 
    1.685687e-16, 1.692723e-16, 1.6817e-16, 1.685021e-16, 1.68733e-16, 
    1.686318e-16, 1.691572e-16, 1.692809e-16, 1.697831e-16, 1.695236e-16, 
    1.710656e-16, 1.703842e-16, 1.72272e-16, 1.717455e-16, 1.681736e-16, 
    1.683421e-16, 1.689279e-16, 1.686493e-16, 1.694456e-16, 1.696413e-16, 
    1.698004e-16, 1.700035e-16, 1.700255e-16, 1.701458e-16, 1.699487e-16, 
    1.701381e-16, 1.694209e-16, 1.697416e-16, 1.688611e-16, 1.690755e-16, 
    1.689769e-16, 1.688687e-16, 1.692027e-16, 1.695581e-16, 1.695658e-16, 
    1.696797e-16, 1.7e-16, 1.694489e-16, 1.711532e-16, 1.701014e-16, 
    1.685258e-16, 1.688498e-16, 1.688962e-16, 1.687707e-16, 1.696217e-16, 
    1.693136e-16, 1.701429e-16, 1.69919e-16, 1.702858e-16, 1.701036e-16, 
    1.700768e-16, 1.698426e-16, 1.696966e-16, 1.693277e-16, 1.690273e-16, 
    1.68789e-16, 1.688444e-16, 1.691062e-16, 1.695798e-16, 1.700275e-16, 
    1.699294e-16, 1.70258e-16, 1.69388e-16, 1.69753e-16, 1.696119e-16, 
    1.699796e-16, 1.691735e-16, 1.698596e-16, 1.689978e-16, 1.690735e-16, 
    1.693075e-16, 1.697776e-16, 1.698818e-16, 1.699927e-16, 1.699243e-16, 
    1.695919e-16, 1.695375e-16, 1.693018e-16, 1.692367e-16, 1.69057e-16, 
    1.689082e-16, 1.690442e-16, 1.691869e-16, 1.695921e-16, 1.699568e-16, 
    1.70354e-16, 1.704512e-16, 1.709143e-16, 1.705372e-16, 1.71159e-16, 
    1.706301e-16, 1.715453e-16, 1.698996e-16, 1.706148e-16, 1.693182e-16, 
    1.694581e-16, 1.69711e-16, 1.702905e-16, 1.699779e-16, 1.703436e-16, 
    1.695353e-16, 1.691151e-16, 1.690065e-16, 1.688034e-16, 1.690111e-16, 
    1.689942e-16, 1.691929e-16, 1.691291e-16, 1.696055e-16, 1.693497e-16, 
    1.70076e-16, 1.703407e-16, 1.710872e-16, 1.715439e-16, 1.720084e-16, 
    1.722132e-16, 1.722755e-16, 1.723016e-16 ;

 CWDC_vr =
  5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110342e-05, 5.110341e-05, 
    5.110342e-05, 5.110341e-05, 5.110341e-05, 5.11034e-05, 5.11034e-05, 
    5.11034e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 
    5.11034e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 5.11034e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.11034e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.11034e-05, 5.11034e-05, 
    5.11034e-05, 5.11034e-05, 5.110341e-05, 5.110341e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 5.11034e-05, 
    5.110341e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 
    5.110342e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 5.110343e-05, 
    5.110343e-05, 5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 
    5.11034e-05, 5.110343e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110341e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 
    5.11034e-05, 5.11034e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110342e-05, 
    5.110341e-05, 5.110341e-05, 5.110342e-05, 5.110341e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110341e-05, 5.110341e-05, 5.11034e-05, 5.110341e-05, 5.11034e-05, 
    5.11034e-05, 5.11034e-05, 5.110339e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110342e-05, 5.110341e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.11034e-05, 5.11034e-05, 5.110339e-05, 5.110339e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.11034e-05, 5.110341e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.11034e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.11034e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110342e-05, 5.110341e-05, 5.110342e-05, 5.110342e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110341e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 
    5.11034e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 
    5.11034e-05, 5.11034e-05, 5.110341e-05, 5.11034e-05, 5.110341e-05, 
    5.110341e-05, 5.110341e-05, 5.11034e-05, 5.110341e-05, 5.11034e-05, 
    5.110341e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110342e-05, 
    5.110342e-05, 5.110342e-05, 5.110342e-05, 5.110341e-05, 5.110341e-05, 
    5.110341e-05, 5.11034e-05, 5.11034e-05, 5.11034e-05, 5.110339e-05, 
    5.110339e-05, 5.110339e-05, 5.110339e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDN =
  1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789929e-09, 
    1.78993e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789929e-09, 1.78993e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789929e-09, 1.78993e-09, 1.789929e-09, 1.78993e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789929e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789929e-09, 1.78993e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789929e-09, 1.789929e-09, 1.78993e-09, 1.789929e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789929e-09, 1.78993e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.78993e-09, 1.789929e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.789929e-09, 1.789929e-09, 1.78993e-09, 1.789929e-09, 1.789929e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789929e-09, 
    1.78993e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.78993e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.78993e-09, 1.789929e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.78993e-09, 
    1.78993e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09, 1.789929e-09, 1.78993e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 1.789929e-09, 
    1.789929e-09, 1.789929e-09, 1.789929e-09 ;

 CWDN_TO_LITR2N =
  1.059298e-18, 1.061996e-18, 1.061472e-18, 1.063645e-18, 1.06244e-18, 
    1.063863e-18, 1.059846e-18, 1.062103e-18, 1.060662e-18, 1.059542e-18, 
    1.067856e-18, 1.063742e-18, 1.072126e-18, 1.069508e-18, 1.076082e-18, 
    1.071718e-18, 1.07696e-18, 1.075957e-18, 1.078979e-18, 1.078113e-18, 
    1.081972e-18, 1.079378e-18, 1.083971e-18, 1.081353e-18, 1.081763e-18, 
    1.079292e-18, 1.064572e-18, 1.067344e-18, 1.064407e-18, 1.064803e-18, 
    1.064626e-18, 1.062465e-18, 1.061375e-18, 1.059093e-18, 1.059507e-18, 
    1.061184e-18, 1.064981e-18, 1.063693e-18, 1.066939e-18, 1.066866e-18, 
    1.070473e-18, 1.068847e-18, 1.074903e-18, 1.073184e-18, 1.078149e-18, 
    1.076902e-18, 1.078091e-18, 1.07773e-18, 1.078095e-18, 1.076265e-18, 
    1.077049e-18, 1.075438e-18, 1.069152e-18, 1.071001e-18, 1.065481e-18, 
    1.062155e-18, 1.059945e-18, 1.058375e-18, 1.058597e-18, 1.05902e-18, 
    1.061194e-18, 1.063236e-18, 1.064792e-18, 1.065831e-18, 1.066855e-18, 
    1.06995e-18, 1.071588e-18, 1.07525e-18, 1.074591e-18, 1.075709e-18, 
    1.076778e-18, 1.07857e-18, 1.078275e-18, 1.079064e-18, 1.07568e-18, 
    1.077929e-18, 1.074215e-18, 1.075231e-18, 1.06713e-18, 1.064041e-18, 
    1.062724e-18, 1.061573e-18, 1.058768e-18, 1.060705e-18, 1.059941e-18, 
    1.061758e-18, 1.062911e-18, 1.062341e-18, 1.06586e-18, 1.064492e-18, 
    1.071685e-18, 1.06859e-18, 1.076653e-18, 1.074726e-18, 1.077115e-18, 
    1.075896e-18, 1.077983e-18, 1.076105e-18, 1.079358e-18, 1.080065e-18, 
    1.079582e-18, 1.081439e-18, 1.076001e-18, 1.07809e-18, 1.062325e-18, 
    1.062418e-18, 1.062852e-18, 1.060945e-18, 1.060829e-18, 1.059081e-18, 
    1.060637e-18, 1.061298e-18, 1.062979e-18, 1.063971e-18, 1.064915e-18, 
    1.066988e-18, 1.069301e-18, 1.072532e-18, 1.074851e-18, 1.076404e-18, 
    1.075452e-18, 1.076293e-18, 1.075353e-18, 1.074913e-18, 1.0798e-18, 
    1.077057e-18, 1.081172e-18, 1.080944e-18, 1.079083e-18, 1.08097e-18, 
    1.062484e-18, 1.061948e-18, 1.060088e-18, 1.061544e-18, 1.058891e-18, 
    1.060376e-18, 1.061229e-18, 1.06452e-18, 1.065243e-18, 1.065913e-18, 
    1.067235e-18, 1.068931e-18, 1.071902e-18, 1.074484e-18, 1.07684e-18, 
    1.076667e-18, 1.076728e-18, 1.077254e-18, 1.075951e-18, 1.077467e-18, 
    1.077721e-18, 1.077057e-18, 1.080914e-18, 1.079813e-18, 1.08094e-18, 
    1.080223e-18, 1.062122e-18, 1.063023e-18, 1.062536e-18, 1.063451e-18, 
    1.062806e-18, 1.065671e-18, 1.06653e-18, 1.070542e-18, 1.068897e-18, 
    1.071516e-18, 1.069164e-18, 1.06958e-18, 1.0716e-18, 1.069291e-18, 
    1.074341e-18, 1.070917e-18, 1.077274e-18, 1.073858e-18, 1.077488e-18, 
    1.07683e-18, 1.07792e-18, 1.078895e-18, 1.080122e-18, 1.082384e-18, 
    1.08186e-18, 1.083751e-18, 1.064365e-18, 1.065532e-18, 1.06543e-18, 
    1.066651e-18, 1.067553e-18, 1.069509e-18, 1.072641e-18, 1.071464e-18, 
    1.073625e-18, 1.074058e-18, 1.070775e-18, 1.072791e-18, 1.066313e-18, 
    1.06736e-18, 1.066737e-18, 1.064457e-18, 1.071734e-18, 1.068002e-18, 
    1.074889e-18, 1.072871e-18, 1.078756e-18, 1.075831e-18, 1.081572e-18, 
    1.08402e-18, 1.086325e-18, 1.089011e-18, 1.066169e-18, 1.065377e-18, 
    1.066796e-18, 1.068758e-18, 1.070578e-18, 1.072994e-18, 1.073242e-18, 
    1.073694e-18, 1.074865e-18, 1.07585e-18, 1.073836e-18, 1.076097e-18, 
    1.067602e-18, 1.072058e-18, 1.065076e-18, 1.06718e-18, 1.068642e-18, 
    1.068002e-18, 1.071329e-18, 1.072113e-18, 1.075293e-18, 1.07365e-18, 
    1.083416e-18, 1.0791e-18, 1.091056e-18, 1.087721e-18, 1.0651e-18, 
    1.066167e-18, 1.069877e-18, 1.068112e-18, 1.073156e-18, 1.074395e-18, 
    1.075403e-18, 1.076689e-18, 1.076828e-18, 1.07759e-18, 1.076342e-18, 
    1.077541e-18, 1.072999e-18, 1.07503e-18, 1.069454e-18, 1.070812e-18, 
    1.070187e-18, 1.069502e-18, 1.071617e-18, 1.073868e-18, 1.073917e-18, 
    1.074638e-18, 1.076667e-18, 1.073176e-18, 1.08397e-18, 1.077309e-18, 
    1.06733e-18, 1.069382e-18, 1.069676e-18, 1.068881e-18, 1.074271e-18, 
    1.072319e-18, 1.077572e-18, 1.076154e-18, 1.078477e-18, 1.077323e-18, 
    1.077153e-18, 1.07567e-18, 1.074745e-18, 1.072409e-18, 1.070506e-18, 
    1.068997e-18, 1.069348e-18, 1.071006e-18, 1.074006e-18, 1.076841e-18, 
    1.07622e-18, 1.078301e-18, 1.07279e-18, 1.075102e-18, 1.074209e-18, 
    1.076538e-18, 1.071432e-18, 1.075778e-18, 1.07032e-18, 1.070799e-18, 
    1.072281e-18, 1.075258e-18, 1.075918e-18, 1.07662e-18, 1.076187e-18, 
    1.074082e-18, 1.073737e-18, 1.072245e-18, 1.071832e-18, 1.070695e-18, 
    1.069752e-18, 1.070613e-18, 1.071517e-18, 1.074083e-18, 1.076393e-18, 
    1.078909e-18, 1.079524e-18, 1.082457e-18, 1.080069e-18, 1.084007e-18, 
    1.080657e-18, 1.086454e-18, 1.076031e-18, 1.08056e-18, 1.072348e-18, 
    1.073235e-18, 1.074836e-18, 1.078507e-18, 1.076527e-18, 1.078842e-18, 
    1.073724e-18, 1.071062e-18, 1.070374e-18, 1.069088e-18, 1.070404e-18, 
    1.070297e-18, 1.071555e-18, 1.071151e-18, 1.074168e-18, 1.072548e-18, 
    1.077148e-18, 1.078824e-18, 1.083552e-18, 1.086445e-18, 1.089387e-18, 
    1.090684e-18, 1.091078e-18, 1.091243e-18 ;

 CWDN_TO_LITR3N =
  3.345153e-19, 3.353671e-19, 3.352017e-19, 3.35888e-19, 3.355075e-19, 
    3.359567e-19, 3.346882e-19, 3.354008e-19, 3.34946e-19, 3.345922e-19, 
    3.372179e-19, 3.359187e-19, 3.385662e-19, 3.377392e-19, 3.398152e-19, 
    3.384374e-19, 3.400928e-19, 3.397758e-19, 3.407301e-19, 3.404569e-19, 
    3.416753e-19, 3.408562e-19, 3.423066e-19, 3.4148e-19, 3.416092e-19, 
    3.408291e-19, 3.361806e-19, 3.370561e-19, 3.361286e-19, 3.362536e-19, 
    3.361976e-19, 3.355153e-19, 3.351709e-19, 3.344503e-19, 3.345813e-19, 
    3.351106e-19, 3.363097e-19, 3.359031e-19, 3.369281e-19, 3.36905e-19, 
    3.380442e-19, 3.375308e-19, 3.394432e-19, 3.389002e-19, 3.404683e-19, 
    3.400742e-19, 3.404497e-19, 3.403359e-19, 3.404512e-19, 3.398732e-19, 
    3.401209e-19, 3.396121e-19, 3.376269e-19, 3.382108e-19, 3.364678e-19, 
    3.354172e-19, 3.347194e-19, 3.342236e-19, 3.342937e-19, 3.344273e-19, 
    3.351137e-19, 3.357588e-19, 3.3625e-19, 3.365783e-19, 3.369016e-19, 
    3.378789e-19, 3.383962e-19, 3.395527e-19, 3.393444e-19, 3.396975e-19, 
    3.40035e-19, 3.406009e-19, 3.405079e-19, 3.40757e-19, 3.396884e-19, 
    3.403987e-19, 3.392257e-19, 3.395467e-19, 3.369885e-19, 3.360129e-19, 
    3.355969e-19, 3.352335e-19, 3.343476e-19, 3.349594e-19, 3.347182e-19, 
    3.352921e-19, 3.356563e-19, 3.354762e-19, 3.365872e-19, 3.361554e-19, 
    3.384269e-19, 3.374494e-19, 3.399957e-19, 3.393872e-19, 3.401415e-19, 
    3.397567e-19, 3.404157e-19, 3.398227e-19, 3.408498e-19, 3.410731e-19, 
    3.409205e-19, 3.41507e-19, 3.397897e-19, 3.404496e-19, 3.354711e-19, 
    3.355004e-19, 3.356374e-19, 3.350353e-19, 3.349985e-19, 3.344467e-19, 
    3.349378e-19, 3.351468e-19, 3.356774e-19, 3.359909e-19, 3.362889e-19, 
    3.369436e-19, 3.37674e-19, 3.386943e-19, 3.394267e-19, 3.399171e-19, 
    3.396164e-19, 3.398818e-19, 3.395851e-19, 3.39446e-19, 3.409894e-19, 
    3.401231e-19, 3.414227e-19, 3.413509e-19, 3.407629e-19, 3.41359e-19, 
    3.355211e-19, 3.353521e-19, 3.347646e-19, 3.352244e-19, 3.343866e-19, 
    3.348555e-19, 3.35125e-19, 3.361642e-19, 3.363926e-19, 3.36604e-19, 
    3.370216e-19, 3.375571e-19, 3.384953e-19, 3.393109e-19, 3.400547e-19, 
    3.400002e-19, 3.400194e-19, 3.401853e-19, 3.397741e-19, 3.402529e-19, 
    3.403331e-19, 3.401231e-19, 3.413412e-19, 3.409935e-19, 3.413493e-19, 
    3.41123e-19, 3.35407e-19, 3.356915e-19, 3.355378e-19, 3.358267e-19, 
    3.356231e-19, 3.365278e-19, 3.367988e-19, 3.38066e-19, 3.375465e-19, 
    3.383734e-19, 3.376306e-19, 3.377622e-19, 3.384e-19, 3.376708e-19, 
    3.392657e-19, 3.381844e-19, 3.401918e-19, 3.39113e-19, 3.402593e-19, 
    3.400515e-19, 3.403957e-19, 3.407037e-19, 3.410912e-19, 3.418053e-19, 
    3.416401e-19, 3.422371e-19, 3.361154e-19, 3.364838e-19, 3.364516e-19, 
    3.368371e-19, 3.371221e-19, 3.377396e-19, 3.387286e-19, 3.383569e-19, 
    3.390394e-19, 3.391762e-19, 3.381395e-19, 3.38776e-19, 3.367304e-19, 
    3.370611e-19, 3.368644e-19, 3.361443e-19, 3.384423e-19, 3.372638e-19, 
    3.394387e-19, 3.388014e-19, 3.406598e-19, 3.39736e-19, 3.415491e-19, 
    3.423222e-19, 3.430499e-19, 3.438982e-19, 3.36685e-19, 3.364348e-19, 
    3.36883e-19, 3.375024e-19, 3.380772e-19, 3.388403e-19, 3.389184e-19, 
    3.390612e-19, 3.394312e-19, 3.397421e-19, 3.391062e-19, 3.3982e-19, 
    3.371374e-19, 3.385446e-19, 3.363399e-19, 3.370042e-19, 3.37466e-19, 
    3.372637e-19, 3.383145e-19, 3.385618e-19, 3.395661e-19, 3.390472e-19, 
    3.421312e-19, 3.407685e-19, 3.445441e-19, 3.43491e-19, 3.363473e-19, 
    3.366843e-19, 3.378558e-19, 3.372986e-19, 3.388913e-19, 3.392827e-19, 
    3.396009e-19, 3.400071e-19, 3.400511e-19, 3.402917e-19, 3.398974e-19, 
    3.402762e-19, 3.388419e-19, 3.394832e-19, 3.377222e-19, 3.381511e-19, 
    3.379539e-19, 3.377374e-19, 3.384054e-19, 3.391161e-19, 3.391316e-19, 
    3.393593e-19, 3.4e-19, 3.388978e-19, 3.423063e-19, 3.402027e-19, 
    3.370516e-19, 3.376996e-19, 3.377925e-19, 3.375415e-19, 3.392434e-19, 
    3.386272e-19, 3.402858e-19, 3.39838e-19, 3.405717e-19, 3.402072e-19, 
    3.401535e-19, 3.396851e-19, 3.393933e-19, 3.386554e-19, 3.380546e-19, 
    3.375779e-19, 3.376888e-19, 3.382123e-19, 3.391597e-19, 3.400549e-19, 
    3.398589e-19, 3.40516e-19, 3.387759e-19, 3.395059e-19, 3.392238e-19, 
    3.399593e-19, 3.38347e-19, 3.397192e-19, 3.379957e-19, 3.38147e-19, 
    3.38615e-19, 3.395552e-19, 3.397635e-19, 3.399853e-19, 3.398485e-19, 
    3.391838e-19, 3.390749e-19, 3.386037e-19, 3.384733e-19, 3.381141e-19, 
    3.378164e-19, 3.380883e-19, 3.383737e-19, 3.391842e-19, 3.399136e-19, 
    3.40708e-19, 3.409025e-19, 3.418285e-19, 3.410743e-19, 3.42318e-19, 
    3.412601e-19, 3.430906e-19, 3.397992e-19, 3.412296e-19, 3.386363e-19, 
    3.389163e-19, 3.394219e-19, 3.40581e-19, 3.399559e-19, 3.406871e-19, 
    3.390707e-19, 3.382302e-19, 3.38013e-19, 3.376069e-19, 3.380223e-19, 
    3.379885e-19, 3.383858e-19, 3.382581e-19, 3.392111e-19, 3.386994e-19, 
    3.401521e-19, 3.406814e-19, 3.421744e-19, 3.430878e-19, 3.440169e-19, 
    3.444264e-19, 3.445511e-19, 3.446031e-19 ;

 CWDN_vr =
  1.022069e-07, 1.022068e-07, 1.022069e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022069e-07, 1.022068e-07, 1.022069e-07, 1.022069e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 1.022068e-07, 
    1.022068e-07, 1.022068e-07, 1.022068e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADSTEMC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 DEADSTEMN =
  6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05 ;

 DENIT =
  2.431536e-36, 2.080171e-35, 1.377042e-35, 7.51097e-35, 2.945023e-35, 
    8.881373e-35, 3.775778e-36, 2.262524e-35, 7.249973e-36, 2.95697e-36, 
    1.808846e-33, 8.093939e-35, 3.946951e-32, 6.045991e-33, 6.088165e-31, 
    2.958383e-32, 1.100823e-30, 5.589807e-31, 4.199307e-30, 2.372932e-30, 
    2.909635e-29, 5.454859e-30, 1.022441e-28, 1.959256e-29, 2.545516e-29, 
    5.157598e-30, 1.529097e-34, 1.237951e-33, 1.348288e-34, 1.824726e-34, 
    1.593225e-34, 3.003121e-35, 1.276494e-35, 2.058065e-36, 2.875827e-36, 
    1.096847e-35, 2.089805e-34, 7.787286e-35, 9.12848e-34, 8.643058e-34, 
    1.214609e-32, 3.736812e-33, 2.72498e-31, 8.287591e-32, 2.430399e-30, 
    1.057477e-30, 2.337914e-30, 1.840018e-30, 2.345202e-30, 6.887896e-31, 
    1.167867e-30, 3.928743e-31, 4.667509e-33, 1.773161e-32, 3.054395e-34, 
    2.358835e-35, 4.088082e-36, 1.149436e-36, 1.377033e-36, 1.940986e-36, 
    1.105402e-35, 5.469746e-35, 1.807634e-34, 3.977145e-34, 8.575428e-34, 
    8.34156e-33, 2.69561e-32, 3.457341e-31, 2.197837e-31, 4.725023e-31, 
    9.728318e-31, 3.209095e-30, 2.641e-30, 4.442478e-30, 4.630589e-31, 
    2.100941e-30, 1.695494e-31, 3.410151e-31, 1.055934e-33, 1.017697e-34, 
    3.678611e-35, 1.490986e-35, 1.581801e-36, 7.500951e-36, 4.076749e-36, 
    1.724691e-35, 4.25128e-35, 2.724771e-35, 4.063328e-34, 1.438516e-34, 
    2.887758e-32, 3.095547e-33, 8.94634e-31, 2.41262e-31, 1.219711e-30, 
    5.363627e-31, 2.177187e-30, 6.179375e-31, 5.384613e-30, 8.539326e-30, 
    6.233685e-30, 2.06851e-29, 5.758325e-31, 2.338045e-30, 2.691009e-35, 
    2.894075e-35, 4.057476e-35, 9.080108e-36, 8.27686e-36, 2.039305e-36, 
    7.101458e-36, 1.200639e-35, 4.477733e-35, 9.648016e-35, 1.986333e-34, 
    9.472638e-34, 5.205024e-33, 5.251311e-32, 2.62879e-31, 7.563291e-31, 
    3.964653e-31, 7.014704e-31, 3.705541e-31, 2.741184e-31, 7.187649e-30, 
    1.173657e-30, 1.743426e-29, 1.506449e-29, 4.497641e-30, 1.531475e-29, 
    3.04559e-35, 2.002432e-35, 4.583814e-36, 1.456866e-35, 1.747991e-36, 
    5.770927e-36, 1.137196e-35, 1.470528e-34, 2.549317e-34, 4.230895e-34, 
    1.138245e-33, 3.971221e-33, 3.365823e-32, 2.043549e-31, 1.014278e-30, 
    9.032062e-31, 9.408806e-31, 1.338794e-30, 5.567699e-31, 1.544329e-30, 
    1.829777e-30, 1.173308e-30, 1.477218e-29, 7.244453e-30, 1.501769e-29, 
    9.453937e-30, 2.295419e-35, 4.635668e-35, 3.173496e-35, 6.461318e-35, 
    3.918533e-35, 3.528461e-34, 6.730773e-34, 1.277267e-32, 3.875749e-33, 
    2.559798e-32, 4.706361e-33, 6.374028e-33, 2.720699e-32, 5.162966e-33, 
    1.852806e-31, 1.671785e-32, 1.357209e-30, 1.32692e-31, 1.565558e-30, 
    1.007367e-30, 2.086567e-30, 3.976023e-30, 8.858512e-30, 3.775103e-29, 
    2.707442e-29, 8.909693e-29, 1.30531e-34, 3.17464e-34, 2.936628e-34, 
    7.362291e-34, 1.441659e-33, 6.048335e-33, 5.665552e-32, 2.464709e-32, 
    1.126559e-31, 1.521901e-31, 1.507442e-32, 6.296677e-32, 5.718368e-34, 
    1.250379e-33, 7.855341e-34, 1.400796e-34, 2.989184e-32, 2.010164e-33, 
    2.698833e-31, 6.659578e-32, 3.628413e-30, 5.134083e-31, 2.252845e-29, 
    1.054976e-28, 4.337753e-28, 2.162218e-27, 5.131526e-34, 2.820386e-34, 
    8.205746e-34, 3.501788e-33, 1.309011e-32, 7.259584e-32, 8.627697e-32, 
    1.182309e-31, 2.654278e-31, 5.197211e-31, 1.305896e-31, 6.143558e-31, 
    1.497649e-33, 3.758781e-32, 2.246509e-34, 1.09386e-33, 3.217284e-33, 
    2.008247e-33, 2.239435e-32, 3.903964e-32, 3.558205e-31, 1.146259e-31, 
    7.23638e-29, 4.552815e-30, 7.106188e-27, 1.00624e-27, 2.285472e-34, 
    5.120692e-34, 7.901357e-33, 2.178861e-33, 8.125475e-32, 1.921216e-31, 
    3.833498e-31, 9.169636e-31, 1.006659e-30, 1.676492e-30, 7.251408e-31, 
    1.62218e-30, 7.285792e-32, 2.972194e-31, 5.810477e-33, 1.548275e-32, 
    9.881065e-33, 6.016816e-33, 2.748668e-32, 1.334958e-31, 1.379941e-31, 
    2.271224e-31, 9.0572e-31, 8.242193e-32, 1.024441e-28, 1.392712e-30, 
    1.22124e-33, 5.522901e-33, 6.830898e-33, 3.829655e-33, 1.76336e-31, 
    4.519103e-32, 1.655817e-30, 6.386244e-31, 3.018376e-30, 1.402101e-30, 
    1.25149e-30, 4.59802e-31, 2.444659e-31, 4.81349e-32, 1.243548e-32, 
    4.166146e-33, 5.380952e-33, 1.778853e-32, 1.468531e-31, 1.015282e-30, 
    6.682074e-31, 2.686088e-30, 6.2921e-32, 3.123257e-31, 1.689693e-31, 
    8.278788e-31, 2.41056e-32, 4.962282e-31, 1.086891e-32, 1.533495e-32, 
    4.397302e-32, 3.477105e-31, 5.442648e-31, 8.753326e-31, 6.531403e-31, 
    1.547918e-31, 1.218636e-31, 4.286784e-32, 3.203159e-32, 1.422964e-32, 
    7.213664e-33, 1.34234e-32, 2.560963e-32, 1.548728e-31, 7.510358e-31, 
    4.012579e-30, 6.003471e-30, 3.959985e-29, 8.568919e-30, 1.048367e-28, 
    1.256413e-29, 4.701216e-28, 5.885199e-31, 1.178497e-29, 4.611026e-32, 
    8.586307e-32, 2.603937e-31, 3.081409e-30, 8.217949e-31, 3.843672e-30, 
    1.207228e-31, 1.853259e-32, 1.130717e-32, 4.455016e-33, 1.154876e-32, 
    1.069319e-32, 2.629645e-32, 1.971957e-32, 1.642661e-31, 5.306551e-32, 
    1.247989e-30, 3.797551e-30, 7.874024e-29, 4.669595e-28, 2.693259e-27, 
    5.730218e-27, 7.194341e-27, 7.90995e-27 ;

 DISPVEGC =
  0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653 ;

 DISPVEGN =
  0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997 ;

 DSTDEP =
  2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12 ;

 DSTFLXT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_NFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_GRND_LAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 EFLX_LH_TOT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_LH_TOT_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_LH_TOT_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 ELAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 ER =
  7.624269e-08, 7.645139e-08, 7.641083e-08, 7.657911e-08, 7.648578e-08, 
    7.659595e-08, 7.628502e-08, 7.645966e-08, 7.634819e-08, 7.62615e-08, 
    7.690554e-08, 7.658662e-08, 7.723681e-08, 7.70335e-08, 7.754418e-08, 
    7.720516e-08, 7.761253e-08, 7.753444e-08, 7.776953e-08, 7.77022e-08, 
    7.800275e-08, 7.780061e-08, 7.815856e-08, 7.79545e-08, 7.798641e-08, 
    7.779394e-08, 7.665084e-08, 7.686582e-08, 7.663809e-08, 7.666875e-08, 
    7.6655e-08, 7.648769e-08, 7.640334e-08, 7.622676e-08, 7.625883e-08, 
    7.638853e-08, 7.668255e-08, 7.658277e-08, 7.683426e-08, 7.682858e-08, 
    7.710845e-08, 7.698227e-08, 7.745253e-08, 7.731892e-08, 7.7705e-08, 
    7.760792e-08, 7.770044e-08, 7.767239e-08, 7.77008e-08, 7.755842e-08, 
    7.761943e-08, 7.749413e-08, 7.700589e-08, 7.71494e-08, 7.67213e-08, 
    7.646373e-08, 7.629267e-08, 7.617125e-08, 7.618841e-08, 7.622113e-08, 
    7.638929e-08, 7.654739e-08, 7.666784e-08, 7.674839e-08, 7.682777e-08, 
    7.706788e-08, 7.719501e-08, 7.747953e-08, 7.742823e-08, 7.751517e-08, 
    7.759827e-08, 7.773771e-08, 7.771477e-08, 7.777619e-08, 7.75129e-08, 
    7.768788e-08, 7.739899e-08, 7.747801e-08, 7.684923e-08, 7.66097e-08, 
    7.650777e-08, 7.641862e-08, 7.620162e-08, 7.635147e-08, 7.629239e-08, 
    7.643295e-08, 7.652225e-08, 7.647809e-08, 7.67506e-08, 7.664466e-08, 
    7.720254e-08, 7.696229e-08, 7.758857e-08, 7.743876e-08, 7.762448e-08, 
    7.752973e-08, 7.769207e-08, 7.754596e-08, 7.779906e-08, 7.785415e-08, 
    7.78165e-08, 7.796114e-08, 7.753786e-08, 7.770043e-08, 7.647685e-08, 
    7.648405e-08, 7.651761e-08, 7.637008e-08, 7.636106e-08, 7.622587e-08, 
    7.634618e-08, 7.639739e-08, 7.652743e-08, 7.660432e-08, 7.667741e-08, 
    7.683809e-08, 7.701749e-08, 7.72683e-08, 7.744847e-08, 7.75692e-08, 
    7.749518e-08, 7.756054e-08, 7.748747e-08, 7.745323e-08, 7.78335e-08, 
    7.761999e-08, 7.794034e-08, 7.792262e-08, 7.777765e-08, 7.792462e-08, 
    7.648911e-08, 7.644767e-08, 7.630373e-08, 7.641638e-08, 7.621115e-08, 
    7.632602e-08, 7.639206e-08, 7.664685e-08, 7.670285e-08, 7.675474e-08, 
    7.685723e-08, 7.698873e-08, 7.721936e-08, 7.741998e-08, 7.76031e-08, 
    7.758969e-08, 7.759441e-08, 7.76353e-08, 7.7534e-08, 7.765193e-08, 
    7.767171e-08, 7.761997e-08, 7.792025e-08, 7.783448e-08, 7.792224e-08, 
    7.78664e-08, 7.646114e-08, 7.653087e-08, 7.649319e-08, 7.656404e-08, 
    7.651412e-08, 7.673605e-08, 7.680259e-08, 7.711383e-08, 7.698614e-08, 
    7.718939e-08, 7.70068e-08, 7.703915e-08, 7.719597e-08, 7.701667e-08, 
    7.74089e-08, 7.714296e-08, 7.763688e-08, 7.737135e-08, 7.765352e-08, 
    7.760231e-08, 7.768711e-08, 7.776304e-08, 7.785858e-08, 7.803479e-08, 
    7.7994e-08, 7.814135e-08, 7.663483e-08, 7.672524e-08, 7.671731e-08, 
    7.681193e-08, 7.68819e-08, 7.703356e-08, 7.727672e-08, 7.71853e-08, 
    7.735314e-08, 7.738683e-08, 7.713184e-08, 7.728839e-08, 7.678577e-08, 
    7.686698e-08, 7.681864e-08, 7.664195e-08, 7.720634e-08, 7.691673e-08, 
    7.745144e-08, 7.729462e-08, 7.775221e-08, 7.752466e-08, 7.797154e-08, 
    7.816244e-08, 7.834216e-08, 7.855203e-08, 7.677461e-08, 7.671318e-08, 
    7.682319e-08, 7.697533e-08, 7.711654e-08, 7.730418e-08, 7.732339e-08, 
    7.735854e-08, 7.744958e-08, 7.752611e-08, 7.736963e-08, 7.754529e-08, 
    7.688577e-08, 7.723148e-08, 7.668994e-08, 7.685301e-08, 7.696638e-08, 
    7.691667e-08, 7.717485e-08, 7.723568e-08, 7.748282e-08, 7.735509e-08, 
    7.811531e-08, 7.777906e-08, 7.871185e-08, 7.845127e-08, 7.669171e-08, 
    7.677441e-08, 7.706215e-08, 7.692525e-08, 7.731672e-08, 7.741303e-08, 
    7.749135e-08, 7.75914e-08, 7.760222e-08, 7.76615e-08, 7.756436e-08, 
    7.765767e-08, 7.730458e-08, 7.74624e-08, 7.702928e-08, 7.713471e-08, 
    7.708622e-08, 7.703301e-08, 7.719722e-08, 7.737208e-08, 7.737585e-08, 
    7.743191e-08, 7.758979e-08, 7.731831e-08, 7.815863e-08, 7.763973e-08, 
    7.686458e-08, 7.702379e-08, 7.704657e-08, 7.698489e-08, 7.740338e-08, 
    7.725177e-08, 7.766006e-08, 7.754974e-08, 7.77305e-08, 7.764068e-08, 
    7.762746e-08, 7.75121e-08, 7.744025e-08, 7.725872e-08, 7.711099e-08, 
    7.699384e-08, 7.702109e-08, 7.714976e-08, 7.738279e-08, 7.760318e-08, 
    7.755491e-08, 7.771676e-08, 7.728835e-08, 7.7468e-08, 7.739856e-08, 
    7.757962e-08, 7.718286e-08, 7.752063e-08, 7.709649e-08, 7.713369e-08, 
    7.724876e-08, 7.748016e-08, 7.75314e-08, 7.758604e-08, 7.755232e-08, 
    7.738871e-08, 7.736191e-08, 7.724597e-08, 7.721394e-08, 7.71256e-08, 
    7.705243e-08, 7.711927e-08, 7.718945e-08, 7.738879e-08, 7.756837e-08, 
    7.776411e-08, 7.781203e-08, 7.804059e-08, 7.785449e-08, 7.816151e-08, 
    7.790043e-08, 7.835236e-08, 7.754026e-08, 7.789281e-08, 7.725401e-08, 
    7.732286e-08, 7.744735e-08, 7.773286e-08, 7.757877e-08, 7.775899e-08, 
    7.736087e-08, 7.715419e-08, 7.710074e-08, 7.700096e-08, 7.710302e-08, 
    7.709473e-08, 7.719238e-08, 7.7161e-08, 7.739541e-08, 7.72695e-08, 
    7.762712e-08, 7.775758e-08, 7.812591e-08, 7.835159e-08, 7.858132e-08, 
    7.86827e-08, 7.871355e-08, 7.872645e-08 ;

 ERRH2O =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 ERRH2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ERRSEB =
  -2.007119e-14, -1.366582e-14, -3.241549e-15, -6.597626e-15, -4.265041e-15, 
    -1.884864e-14, -1.324156e-14, -8.251574e-15, -1.837742e-14, 
    -1.138665e-14, -1.210905e-14, -2.056087e-14, -1.180924e-14, 
    -1.664112e-14, -1.203695e-14, -1.671759e-14, -1.652374e-14, 
    -1.125482e-14, -1.30244e-14, -7.818122e-15, -2.180944e-14, -1.096261e-14, 
    -5.201353e-15, -6.019445e-15, -9.603353e-15, -1.483239e-14, 
    -1.025013e-14, -6.756047e-15, -1.661544e-14, -1.614295e-14, 
    -6.881167e-15, -1.112722e-14, -1.600763e-14, -1.13442e-14, -1.265143e-14, 
    -1.91349e-14, -1.479986e-14, -2.102611e-15, -1.61931e-14, -1.509392e-14, 
    -1.349152e-14, -9.467587e-15, -9.361921e-15, -1.319489e-14, 
    -9.602935e-15, -1.994978e-14, -9.692799e-16, -1.282387e-14, -1.60067e-14, 
    -1.964966e-14, -1.290968e-14, -1.226271e-14, -1.251061e-14, 
    -1.622766e-14, -6.261795e-15, -9.936405e-15, -1.259307e-14, 
    -1.766568e-14, -7.226534e-15, -7.191836e-15, -1.407728e-14, 
    -1.776976e-14, -1.866601e-14, -1.95773e-14, -1.6935e-14, -1.107892e-14, 
    -1.382747e-14, -4.030503e-15, -1.06531e-14, -1.643464e-14, -1.107834e-14, 
    -1.591279e-14, -1.568626e-14, -1.95338e-14, -1.181907e-14, -1.252906e-14, 
    -1.420834e-14, -1.793077e-14, -1.77925e-14, -1.145636e-14, -5.047017e-15, 
    -9.901436e-15, -6.38005e-15, -1.50444e-14, -4.322892e-15, -2.826569e-15, 
    -1.568549e-14, -1.305029e-14, -1.52943e-14, -1.554663e-14, -3.51218e-15, 
    -1.779581e-14, -1.002707e-14, -1.162984e-14, -7.506522e-15, 
    -9.874957e-15, -2.232139e-14, -1.907007e-14, -1.449535e-14, 
    -1.017113e-14, -9.20002e-15, -1.116339e-14, -7.6961e-15, -9.358887e-15, 
    -1.324198e-14, -8.399997e-15, -1.26799e-14, -1.478658e-14, -1.59689e-14, 
    -1.839882e-14, -9.68586e-15, -2.175982e-14, -9.506885e-15, -1.954163e-14, 
    -4.67566e-15, -1.263808e-14, -9.08237e-15, -1.357164e-14, -2.319897e-14, 
    -1.513274e-14, -7.721535e-15, -5.200644e-15, -1.03444e-14, -1.049187e-14, 
    -1.862618e-14, -1.298381e-14, -1.333174e-14, -1.311501e-14, 
    -1.738857e-14, -1.688002e-14, -1.265217e-14, -1.39654e-14, -1.205243e-14, 
    -1.524435e-14, -8.502917e-15, -1.496143e-14, -7.272767e-15, 
    -1.253273e-14, -1.338625e-14, -7.093512e-15, -1.267674e-14, 
    -1.262097e-14, -1.375574e-14, -3.941916e-15, -1.072792e-14, 
    -7.341345e-15, -1.145292e-14, -9.224558e-15, -1.394089e-14, -1.59955e-14, 
    -1.583335e-14, -7.115256e-15, -1.076913e-14, -1.230403e-14, -8.95914e-15, 
    -1.914874e-14, -9.636403e-15, -1.534415e-14, -8.035194e-15, 
    -1.887698e-14, -1.348808e-14, -4.568745e-15, -1.730229e-14, 
    -7.329457e-15, -1.078682e-14, -2.1635e-14, -1.330791e-14, -1.060414e-14, 
    -1.295378e-14, -1.206049e-14, -1.824246e-14, -9.663241e-15, 
    -7.016344e-15, -9.738152e-15, -1.496831e-14, -1.748319e-14, 
    -1.157735e-14, -2.102913e-14, -1.2381e-14, -1.602954e-14, -5.916491e-15, 
    -1.523324e-14, -8.025671e-15, -1.062633e-14, -1.612032e-14, 
    -1.492312e-14, -1.745233e-14, -1.810222e-14, -7.199849e-15, 
    -1.507294e-14, -1.737095e-14, -1.659519e-14, -1.272181e-14, 
    -1.113225e-14, -8.005447e-15, -1.156856e-14, -1.87056e-14, -1.955835e-14, 
    -1.314187e-14, -1.573696e-14, -8.066377e-15, -1.212809e-14, 
    -1.521929e-14, -1.345569e-14, -1.934479e-14, -1.179581e-14, 
    -1.175917e-14, -1.876593e-15, -9.687542e-15, -7.787882e-15, -9.85074e-15, 
    -5.33605e-15, -1.076245e-14, -1.728866e-14, -5.235323e-15, -1.874688e-14, 
    -1.014362e-14, -7.178552e-15, -8.675306e-15, -1.177484e-14, -7.06222e-16, 
    -1.312817e-14, -1.476245e-14, -1.506928e-14, -1.298148e-14, -1.39105e-14, 
    -1.249644e-14, -1.440014e-14, -1.551602e-14, -1.198664e-14, -1.21761e-14, 
    -1.366655e-14, -6.942706e-15, -1.295717e-14, -1.545866e-14, 
    -1.152939e-14, -9.027658e-15, -1.145598e-14, -1.181032e-14, 
    -1.603682e-14, -4.889895e-15, -1.75935e-14, -1.292395e-14, -8.923012e-15, 
    -1.673369e-14, -1.258512e-14, -1.108591e-14, -1.399409e-14, 
    -7.457182e-15, -1.64122e-14, -8.607935e-15, -8.878762e-15, -1.124589e-14, 
    -7.730245e-15, -5.600436e-15, -1.384944e-14, -3.981777e-15, 
    -1.505966e-14, -1.000202e-14, -1.050482e-14, -1.228205e-14, -1.05349e-14, 
    -5.721513e-15, -8.882818e-15, -1.09471e-14, -1.118786e-14, -1.237509e-14, 
    -1.048313e-14, -1.731227e-14, -1.368959e-14, -1.530431e-14, 
    -9.666309e-15, -1.323466e-14, -1.619833e-14, -1.313455e-14, 
    -1.514604e-14, -2.034377e-14, -1.057459e-14, -1.671918e-14, 
    -1.702701e-14, -1.732662e-14, -1.368996e-14, -1.672751e-14, 
    -1.321559e-14, -1.497206e-14, -2.460066e-14, -1.016085e-14, 
    -1.531155e-14, -5.891083e-16, -1.072591e-14, -1.537694e-14, -1.9883e-14, 
    -1.91562e-14, -9.263212e-15, -4.203211e-15, -1.027535e-14, -1.061499e-14, 
    -1.233196e-14, -6.525952e-15, -1.015936e-14, -1.472895e-14, -1.80287e-14, 
    -6.182305e-15, -1.315481e-14, -1.320038e-14, -1.150775e-14, 
    -1.673071e-14, -3.366315e-15, -9.274251e-15, -1.281183e-14, 
    -1.295025e-14, -1.444418e-14, -1.268325e-14, -6.590459e-15, 
    -1.366477e-14, -1.695281e-14, -1.255243e-14, -2.836847e-15, 
    -1.700572e-14, -1.336419e-14, -1.823606e-14, -6.164859e-15, 
    -1.129071e-14, -1.389389e-14, -1.526244e-14, -1.541568e-14, 
    -1.478356e-14, -1.911321e-14, -1.113325e-14, -9.102449e-15, 
    -6.848813e-15, -8.636871e-15, -7.142085e-15, -1.081356e-14, 
    -1.622819e-14, -3.96578e-15, -1.098838e-14, -1.551977e-14 ;

 ERRSOI =
  -8.048863e-11, -3.97242e-10, -3.187638e-10, -4.03303e-10, -2.853823e-10, 
    -2.161533e-10, -1.712507e-10, -3.063577e-10, -2.648181e-10, 
    -1.037775e-10, -3.834113e-10, -2.007011e-10, -3.231118e-10, 
    -2.849667e-10, -4.186552e-10, -3.046396e-10, -4.320107e-10, 
    -2.269567e-10, -4.096626e-10, -3.435573e-10, -1.865147e-10, 
    -3.289711e-10, -4.646109e-10, -2.680339e-10, -3.983319e-10, 
    -1.455538e-10, -4.804039e-10, -4.309356e-10, -4.679829e-10, 
    -2.216097e-10, -5.045026e-10, -1.305089e-10, -4.496219e-10, 
    -4.687175e-10, -4.733516e-10, -1.948928e-10, -3.317407e-10, 
    -2.224785e-10, -4.918345e-10, -4.364206e-10, -4.160843e-10, 
    -2.091114e-10, -2.13617e-10, -2.774738e-10, -3.621708e-10, -6.860227e-10, 
    -3.236457e-10, -2.523015e-10, -2.877982e-10, -5.536701e-10, 
    -4.475925e-10, -4.705755e-10, -6.016838e-10, -4.009116e-10, 
    -3.743745e-10, -4.205823e-10, -2.198752e-10, -3.735751e-10, 
    -1.973089e-10, -2.849583e-10, -1.611356e-10, -3.23965e-10, -2.394723e-10, 
    -2.953624e-10, -3.759499e-10, -3.649166e-10, -3.111579e-10, 
    -4.570612e-10, -2.305265e-10, -3.156915e-10, -4.312044e-10, -4.63283e-10, 
    -1.665717e-10, -3.479139e-10, -3.47553e-10, -4.434259e-10, -2.997262e-10, 
    -3.938031e-10, -3.116829e-10, -2.64079e-10, -1.651201e-10, -4.094064e-10, 
    -2.607516e-10, -2.287185e-10, -2.546865e-10, -3.986035e-10, 
    -3.444579e-10, -3.588518e-10, -2.407131e-10, -2.01996e-10, -3.524542e-10, 
    -4.479509e-10, -4.722838e-10, -3.360084e-10, -4.507024e-10, 
    -4.764674e-10, -5.201897e-10, -5.38838e-10, -2.46405e-10, -5.50967e-10, 
    -2.884743e-10, -6.740776e-11, -4.703515e-10, -1.061135e-10, 
    -3.788421e-10, -3.63254e-10, -3.219359e-10, -3.027329e-10, -3.522666e-10, 
    -3.7395e-10, -1.096604e-10, -2.518263e-10, -1.764514e-10, -3.120086e-10, 
    -2.247462e-10, -3.3298e-10, -5.478819e-10, -2.415503e-10, -4.069075e-10, 
    -7.926968e-11, -3.475163e-10, -5.839325e-11, -3.740478e-10, 
    -3.927928e-10, -3.34011e-10, -4.424542e-10, -3.914929e-10, -3.913092e-10, 
    -2.732514e-10, -2.425334e-10, -2.706682e-10, -2.278333e-10, 
    -3.148918e-10, -3.857851e-10, -2.249097e-10, -2.262659e-10, 
    -3.155241e-10, -4.957735e-10, -3.030754e-10, -4.452738e-10, -3.52092e-10, 
    -6.837193e-11, -3.477816e-10, -3.122415e-10, -4.420743e-10, -3.26337e-10, 
    -4.369317e-10, -3.818354e-10, -4.091886e-10, -1.742031e-10, 
    -4.364237e-10, -5.323872e-10, -3.391161e-10, -4.630843e-10, 
    -2.371777e-10, -3.002826e-10, -3.567231e-10, -2.793196e-10, 
    -4.014062e-10, -1.733798e-10, -3.736705e-10, -3.294552e-10, 
    -4.340439e-10, -4.643647e-10, -4.168675e-10, -4.287811e-10, 
    -4.252695e-10, -2.266924e-10, -3.232223e-10, -5.672741e-10, 
    -4.201224e-10, -3.846358e-10, -2.245262e-10, -3.260874e-10, 
    -4.160975e-10, -5.629146e-10, -1.891564e-10, -3.255737e-10, 
    -5.713998e-10, -4.851191e-10, -3.044425e-10, -3.278049e-10, 
    -4.016399e-10, -4.521125e-10, -3.019704e-10, -4.375414e-10, 
    -4.546751e-10, -4.355025e-10, -3.585881e-10, -3.156143e-10, 
    -1.657162e-10, -2.354308e-10, -4.262792e-10, -2.416524e-10, 
    -2.250975e-10, -5.115299e-10, -4.424844e-10, -3.978316e-10, -5.0998e-10, 
    -2.46782e-10, -3.665549e-10, -2.996438e-10, -4.571659e-10, -5.771656e-10, 
    -1.806364e-10, -2.726928e-10, -2.499393e-10, -3.683532e-11, 
    -3.669922e-10, -2.706201e-10, -2.35213e-10, -4.595605e-10, -4.636789e-10, 
    -1.790389e-10, -3.701636e-10, -3.185502e-10, -3.448923e-10, 
    -2.401118e-10, -3.378181e-10, -4.053013e-10, -1.458147e-10, 
    -2.935501e-10, -4.627987e-10, -1.769904e-10, -4.57855e-10, -5.78643e-10, 
    -4.194458e-10, -2.818347e-10, -3.804506e-10, -2.291996e-10, 
    -2.819111e-10, -3.719031e-10, -1.099823e-10, -1.264338e-10, -2.72408e-10, 
    -2.89765e-10, -3.922665e-10, -4.575852e-10, -3.336472e-10, -2.565268e-10, 
    -2.770858e-10, -6.718894e-10, -3.743198e-10, -3.250572e-10, -6.11653e-10, 
    -4.863034e-10, -3.368414e-10, -2.806706e-10, -3.228382e-10, 
    -4.888028e-10, -3.03749e-10, -3.508355e-10, -2.622868e-10, -3.514159e-10, 
    -3.452259e-10, -3.813019e-10, -6.654689e-11, -3.817796e-10, 
    -4.240483e-10, -4.710458e-10, -1.401679e-10, -3.265515e-10, 
    -3.720877e-10, -3.923254e-10, -2.335067e-10, -4.204855e-10, 
    -3.052902e-10, -3.423292e-10, -3.209962e-10, -3.190558e-10, 
    -3.604795e-10, -3.503365e-10, -4.084202e-10, -4.530886e-10, 
    -4.356056e-10, -1.306295e-10, -1.75136e-10, -2.533539e-10, -4.558277e-10, 
    -3.721091e-10, -2.816972e-10, -3.396096e-10, -1.271771e-10, 
    -3.058283e-10, -2.568376e-10, -3.854115e-10, -3.538196e-10, 
    -2.807986e-10, -1.766646e-10, -2.50865e-10, -3.415662e-10, -3.644123e-10, 
    -1.880697e-10, -3.168743e-10, -3.160603e-10, -3.785413e-10, -2.69903e-10, 
    -3.998442e-10, -1.516195e-10, -2.614735e-10, -4.630906e-10, 
    -3.135462e-10, -3.237159e-10, -4.514983e-10, -3.417157e-10, 
    -2.421217e-10, -3.499859e-10, -3.205066e-10, -2.859853e-10, 
    -1.422836e-11, -3.157095e-10, -3.601544e-10, -4.57829e-10, -2.487897e-10, 
    -2.087632e-10, -1.701543e-10, -1.682667e-10, -7.170208e-10, 
    -4.162676e-10, -3.101993e-10, -3.098456e-10, -3.228534e-10, 
    -2.680164e-10, -5.156883e-10, -3.402701e-10, -3.963124e-10, 
    -2.478806e-10, -4.728871e-10, -2.268202e-10, -4.638581e-10, 
    -2.709854e-10, -3.341628e-10, -3.322576e-10, -2.85404e-10, -2.075501e-10, 
    -8.186363e-11, -4.444162e-10, -4.48957e-10 ;

 ERRSOL =
  1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17 ;

 ESAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 FAREA_BURNED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCEV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4 =
  5.976281e-16, 5.914211e-16, 5.926296e-16, 5.876111e-16, 5.90397e-16, 
    5.871082e-16, 5.963718e-16, 5.911738e-16, 5.94494e-16, 5.970708e-16, 
    5.778332e-16, 5.87387e-16, 5.678625e-16, 5.739911e-16, 5.585617e-16, 
    5.688168e-16, 5.56488e-16, 5.588595e-16, 5.517164e-16, 5.537654e-16, 
    5.445999e-16, 5.507701e-16, 5.398351e-16, 5.460757e-16, 5.451002e-16, 
    5.509732e-16, 5.854692e-16, 5.790248e-16, 5.858501e-16, 5.849327e-16, 
    5.853447e-16, 5.903391e-16, 5.928503e-16, 5.981024e-16, 5.971502e-16, 
    5.932926e-16, 5.8452e-16, 5.875032e-16, 5.799783e-16, 5.801486e-16, 
    5.717351e-16, 5.755341e-16, 5.613418e-16, 5.653854e-16, 5.536799e-16, 
    5.566298e-16, 5.538184e-16, 5.546714e-16, 5.538072e-16, 5.581319e-16, 
    5.5628e-16, 5.600818e-16, 5.748233e-16, 5.705003e-16, 5.833611e-16, 
    5.910507e-16, 5.961439e-16, 5.99749e-16, 5.992398e-16, 5.982684e-16, 
    5.9327e-16, 5.885595e-16, 5.849616e-16, 5.82551e-16, 5.801731e-16, 
    5.729526e-16, 5.691239e-16, 5.605227e-16, 5.620786e-16, 5.594428e-16, 
    5.569231e-16, 5.526843e-16, 5.533828e-16, 5.515129e-16, 5.595131e-16, 
    5.541993e-16, 5.62964e-16, 5.605704e-16, 5.795223e-16, 5.86699e-16, 
    5.897381e-16, 5.923972e-16, 5.988481e-16, 5.943953e-16, 5.961518e-16, 
    5.919713e-16, 5.893096e-16, 5.906266e-16, 5.824851e-16, 5.856542e-16, 
    5.688967e-16, 5.761334e-16, 5.572171e-16, 5.617594e-16, 5.561271e-16, 
    5.590032e-16, 5.540723e-16, 5.585106e-16, 5.508169e-16, 5.491375e-16, 
    5.502852e-16, 5.458742e-16, 5.587563e-16, 5.53818e-16, 5.906633e-16, 
    5.904486e-16, 5.894482e-16, 5.938417e-16, 5.941103e-16, 5.981283e-16, 
    5.945539e-16, 5.930294e-16, 5.891555e-16, 5.868596e-16, 5.846749e-16, 
    5.798628e-16, 5.744738e-16, 5.669128e-16, 5.614652e-16, 5.578053e-16, 
    5.600505e-16, 5.580684e-16, 5.602839e-16, 5.613217e-16, 5.497667e-16, 
    5.562626e-16, 5.465092e-16, 5.470502e-16, 5.514683e-16, 5.469893e-16, 
    5.902978e-16, 5.915333e-16, 5.958154e-16, 5.924651e-16, 5.985654e-16, 
    5.951527e-16, 5.931873e-16, 5.855872e-16, 5.839143e-16, 5.823606e-16, 
    5.792892e-16, 5.753399e-16, 5.683907e-16, 5.623271e-16, 5.567765e-16, 
    5.571838e-16, 5.570404e-16, 5.557981e-16, 5.588733e-16, 5.552929e-16, 
    5.54691e-16, 5.562638e-16, 5.471227e-16, 5.497383e-16, 5.470617e-16, 
    5.487653e-16, 5.911319e-16, 5.890523e-16, 5.901762e-16, 5.880619e-16, 
    5.895514e-16, 5.829184e-16, 5.809253e-16, 5.71571e-16, 5.754175e-16, 
    5.692945e-16, 5.747969e-16, 5.738211e-16, 5.690928e-16, 5.744982e-16, 
    5.626611e-16, 5.706925e-16, 5.557499e-16, 5.637957e-16, 5.552445e-16, 
    5.568005e-16, 5.54224e-16, 5.519133e-16, 5.490035e-16, 5.436227e-16, 
    5.4487e-16, 5.40363e-16, 5.859482e-16, 5.832427e-16, 5.834818e-16, 
    5.806474e-16, 5.785484e-16, 5.7399e-16, 5.666596e-16, 5.694195e-16, 
    5.643506e-16, 5.633312e-16, 5.710314e-16, 5.663064e-16, 5.814306e-16, 
    5.789945e-16, 5.804458e-16, 5.857345e-16, 5.687828e-16, 5.775012e-16, 
    5.613749e-16, 5.661191e-16, 5.522429e-16, 5.591547e-16, 5.455562e-16, 
    5.397144e-16, 5.342054e-16, 5.277458e-16, 5.817654e-16, 5.836054e-16, 
    5.803103e-16, 5.757407e-16, 5.714915e-16, 5.658299e-16, 5.652501e-16, 
    5.641872e-16, 5.614322e-16, 5.591127e-16, 5.638503e-16, 5.585309e-16, 
    5.784276e-16, 5.680248e-16, 5.843e-16, 5.794129e-16, 5.760107e-16, 
    5.775046e-16, 5.697349e-16, 5.678995e-16, 5.604236e-16, 5.64292e-16, 
    5.41157e-16, 5.514239e-16, 5.228174e-16, 5.308488e-16, 5.842477e-16, 
    5.817721e-16, 5.731285e-16, 5.77247e-16, 5.654518e-16, 5.625379e-16, 
    5.601668e-16, 5.571305e-16, 5.56803e-16, 5.550017e-16, 5.579525e-16, 
    5.551187e-16, 5.658178e-16, 5.610435e-16, 5.741191e-16, 5.70944e-16, 
    5.724055e-16, 5.740069e-16, 5.690602e-16, 5.637756e-16, 5.636637e-16, 
    5.61966e-16, 5.571722e-16, 5.654039e-16, 5.398261e-16, 5.556571e-16, 
    5.790689e-16, 5.742814e-16, 5.735983e-16, 5.754559e-16, 5.628302e-16, 
    5.674132e-16, 5.550458e-16, 5.583959e-16, 5.529044e-16, 5.556349e-16, 
    5.560363e-16, 5.595376e-16, 5.617142e-16, 5.672031e-16, 5.716585e-16, 
    5.75187e-16, 5.743657e-16, 5.704899e-16, 5.634522e-16, 5.567728e-16, 
    5.582376e-16, 5.533222e-16, 5.663092e-16, 5.608728e-16, 5.629753e-16, 
    5.574889e-16, 5.694925e-16, 5.592717e-16, 5.720964e-16, 5.709755e-16, 
    5.675041e-16, 5.605028e-16, 5.589523e-16, 5.572935e-16, 5.583175e-16, 
    5.632734e-16, 5.640847e-16, 5.675888e-16, 5.685547e-16, 5.712196e-16, 
    5.734228e-16, 5.714097e-16, 5.692931e-16, 5.632718e-16, 5.578296e-16, 
    5.518802e-16, 5.504222e-16, 5.434418e-16, 5.491243e-16, 5.397374e-16, 
    5.477181e-16, 5.338856e-16, 5.586795e-16, 5.479548e-16, 5.673464e-16, 
    5.652663e-16, 5.614974e-16, 5.528296e-16, 5.575148e-16, 5.520349e-16, 
    5.641166e-16, 5.703555e-16, 5.719679e-16, 5.749726e-16, 5.718993e-16, 
    5.721493e-16, 5.692062e-16, 5.701525e-16, 5.630716e-16, 5.668783e-16, 
    5.560461e-16, 5.520786e-16, 5.408354e-16, 5.339131e-16, 5.268462e-16, 
    5.237186e-16, 5.227659e-16, 5.223674e-16 ;

 FCH4TOCO2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4_DFSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCOV =
  0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584 ;

 FCTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FGEV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FGR =
  -396.58, -397.6065, -397.4086, -398.23, -397.7746, -398.3122, -396.7943, 
    -397.6467, -397.1028, -396.6721, -399.8222, -398.2667, -401.4498, 
    -400.4582, -402.9492, -401.2952, -403.2826, -402.9022, -404.0486, 
    -403.7203, -405.1845, -404.2002, -405.9441, -404.9499, -405.1052, 
    -404.1676, -398.5805, -399.6284, -398.5182, -398.6677, -398.6008, 
    -397.7838, -397.3716, -396.5025, -396.6591, -397.2996, -398.735, 
    -398.2483, -399.476, -399.4483, -400.824, -400.1982, -402.5027, -401.851, 
    -403.734, -403.2606, -403.7117, -403.575, -403.7135, -403.0191, 
    -403.3166, -402.7056, -400.3134, -401.0237, -398.9243, -397.6661, 
    -396.8316, -396.2314, -396.3152, -396.4748, -397.3033, -398.0755, 
    -398.6636, -399.0568, -399.4443, -400.6251, -401.2459, -402.6341, 
    -402.3842, -402.808, -403.2135, -403.8933, -403.7816, -404.0809, 
    -402.7972, -403.6502, -402.2417, -402.627, -399.5473, -398.3797, 
    -397.8813, -397.4466, -396.3795, -397.1186, -396.8302, -397.5168, 
    -397.9527, -397.7372, -399.0676, -398.5504, -401.2827, -400.1004, 
    -403.1662, -402.4356, -403.3414, -402.8793, -403.6707, -402.9585, 
    -404.1925, -404.4608, -404.2774, -404.9825, -402.9189, -403.7115, 
    -397.7311, -397.7662, -397.9301, -397.2095, -397.1655, -396.4981, 
    -397.093, -397.3429, -397.9782, -398.3534, -398.7102, -399.4945, 
    -400.3697, -401.6038, -402.4829, -403.0719, -402.7109, -403.0296, 
    -402.6732, -402.5063, -404.3601, -403.3192, -404.8811, -404.7948, 
    -404.0879, -404.8046, -397.7909, -397.5887, -396.8857, -397.4359, 
    -396.4262, -396.9944, -397.3166, -398.5607, -398.8345, -399.0876, 
    -399.588, -400.2297, -401.365, -402.3438, -403.2372, -403.1718, 
    -403.1948, -403.3941, -402.9001, -403.4752, -403.5715, -403.3194, 
    -404.7833, -404.3652, -404.793, -404.5209, -397.6545, -397.9949, 
    -397.8109, -398.1567, -397.9129, -398.996, -399.3207, -400.8498, 
    -400.2169, -401.2187, -400.3178, -400.4857, -401.2501, -400.3763, 
    -402.2894, -400.9918, -403.4018, -402.1059, -403.4829, -403.2333, 
    -403.6468, -404.0168, -404.4827, -405.3412, -405.1425, -405.8606, 
    -398.5024, -398.9435, -398.9051, -399.3669, -399.7083, -400.4587, 
    -401.645, -401.1991, -402.0181, -402.1823, -400.9384, -401.7018, 
    -399.239, -399.635, -399.3995, -398.537, -401.3013, -399.8779, -402.4973, 
    -401.7324, -403.964, -402.8541, -405.033, -405.9625, -406.8388, -407.86, 
    -399.1847, -398.8849, -399.422, -400.1639, -400.8635, -401.779, 
    -401.8729, -402.0442, -402.4885, -402.8617, -402.098, -402.9553, 
    -399.726, -401.4241, -398.7712, -399.5668, -400.1204, -399.878, 
    -401.1483, -401.445, -402.6502, -402.0275, -405.7328, -404.0944, 
    -408.6385, -407.3696, -398.7801, -399.1838, -400.5979, -399.9199, 
    -401.8403, -402.3101, -402.6922, -403.1799, -403.2328, -403.5218, 
    -403.0482, -403.5032, -401.781, -402.5509, -400.438, -400.9522, 
    -400.7158, -400.4561, -401.2574, -402.1099, -402.1288, -402.4019, 
    -403.1703, -401.8481, -405.9428, -403.414, -399.6239, -400.4104, 
    -400.5221, -400.2111, -402.2629, -401.5233, -403.5148, -402.977, 
    -403.8583, -403.4203, -403.3559, -402.7933, -402.4428, -401.5571, 
    -400.8364, -400.2548, -400.3979, -401.0255, -402.1622, -403.2373, 
    -403.0018, -403.7914, -401.7019, -402.578, -402.2392, -403.1226, 
    -401.1871, -402.8333, -400.7659, -400.9474, -401.5087, -402.6369, 
    -402.8875, -403.1537, -402.9896, -402.1912, -402.0606, -401.4952, 
    -401.3387, -400.9079, -400.5509, -400.8769, -401.2191, -402.1918, 
    -403.0675, -404.022, -404.2558, -405.3685, -404.4618, -405.9568, 
    -404.6844, -406.887, -402.9297, -404.6484, -401.5345, -401.8703, 
    -402.477, -403.8691, -403.1184, -403.9966, -402.0556, -401.0468, 
    -400.7866, -400.2894, -400.7978, -400.7573, -401.2338, -401.0807, 
    -402.2241, -401.61, -403.3541, -403.9899, -405.7851, -406.8842, 
    -408.0034, -408.4968, -408.647, -408.7098 ;

 FGR12 =
  -52.00521, -52.07361, -52.06034, -52.11551, -52.08494, -52.12104, 
    -52.01912, -52.07629, -52.03981, -52.01142, -52.22263, -52.118, 
    -52.33203, -52.26507, -52.43359, -52.32158, -52.45625, -52.43048, 
    -52.50834, -52.48602, -52.58554, -52.51865, -52.63734, -52.56962, 
    -52.58015, -52.51643, -52.13913, -52.20956, -52.13493, -52.14497, 
    -52.14048, -52.08553, -52.05779, -52.00005, -52.01054, -52.05299, 
    -52.14949, -52.11678, -52.19946, -52.19759, -52.28978, -52.24817, 
    -52.40339, -52.35926, -52.48695, -52.4548, -52.48543, -52.47616, 
    -52.48555, -52.43841, -52.45859, -52.41716, -52.25592, -52.30325, 
    -52.16225, -52.07756, -52.0216, -51.98186, -51.98747, -51.99816, 
    -52.05325, -52.10515, -52.14473, -52.1712, -52.19733, -52.27624, 
    -52.31826, -52.41225, -52.39538, -52.42406, -52.45161, -52.49776, 
    -52.49018, -52.5105, -52.42337, -52.48123, -52.38573, -52.41182, 
    -52.20409, -52.12563, -52.09202, -52.06288, -51.99179, -52.04084, 
    -52.0215, -52.06761, -52.0969, -52.08244, -52.17193, -52.13711, 
    -52.32073, -52.24154, -52.44838, -52.39885, -52.46028, -52.42895, 
    -52.48263, -52.43431, -52.5181, -52.53633, -52.52387, -52.57185, 
    -52.43163, -52.48539, -52.08202, -52.08437, -52.09538, -52.04695, 
    -52.04399, -51.99974, -52.03915, -52.05592, -52.09863, -52.12385, 
    -52.14786, -52.20068, -52.25971, -52.34247, -52.40205, -52.44199, 
    -52.41753, -52.43913, -52.41497, -52.40366, -52.52947, -52.45877, 
    -52.56496, -52.55909, -52.51099, -52.55974, -52.08603, -52.07246, 
    -52.02524, -52.06218, -51.99493, -52.03252, -52.05414, -52.13775, 
    -52.15624, -52.17326, -52.207, -52.25028, -52.32635, -52.39259, 
    -52.45322, -52.44877, -52.45034, -52.46386, -52.43035, -52.46936, 
    -52.47589, -52.45879, -52.5583, -52.52986, -52.55896, -52.54046, 
    -52.07688, -52.09974, -52.08738, -52.11061, -52.09423, -52.16705, 
    -52.18893, -52.29147, -52.24942, -52.31643, -52.25624, -52.26693, 
    -52.31848, -52.25957, -52.38887, -52.30106, -52.46437, -52.37643, 
    -52.46989, -52.45296, -52.48104, -52.50616, -52.53785, -52.59625, 
    -52.58275, -52.63168, -52.13388, -52.16354, -52.16099, -52.19209, 
    -52.2151, -52.26512, -52.34529, -52.31516, -52.37056, -52.38168, 
    -52.29753, -52.34912, -52.18346, -52.21011, -52.19428, -52.1362, -52.322, 
    -52.22651, -52.40302, -52.35122, -52.50256, -52.4272, -52.57529, 
    -52.63857, -52.69848, -52.76824, -52.1798, -52.15964, -52.19582, 
    -52.2458, -52.29246, -52.35435, -52.36074, -52.37233, -52.40244, 
    -52.42774, -52.37594, -52.43408, -52.21619, -52.33032, -52.15197, 
    -52.2055, -52.24288, -52.22654, -52.31172, -52.33178, -52.41337, 
    -52.37122, -52.62288, -52.51139, -52.82161, -52.73471, -52.15258, 
    -52.17977, -52.27448, -52.22938, -52.35853, -52.39033, -52.41625, 
    -52.4493, -52.45292, -52.47252, -52.4404, -52.47127, -52.3545, -52.40665, 
    -52.26373, -52.29844, -52.28249, -52.26496, -52.3191, -52.37673, 
    -52.37807, -52.39655, -52.44848, -52.35908, -52.6371, -52.46508, 
    -52.20944, -52.26179, -52.26939, -52.24905, -52.38714, -52.33707, 
    -52.47205, -52.43557, -52.49539, -52.46565, -52.46126, -52.42311, 
    -52.39933, -52.33935, -52.29061, -52.25201, -52.26103, -52.30339, 
    -52.38029, -52.45319, -52.43721, -52.49084, -52.34917, -52.40848, 
    -52.38552, -52.44543, -52.31435, -52.42564, -52.28588, -52.29814, 
    -52.33609, -52.41243, -52.42949, -52.44752, -52.43641, -52.38227, 
    -52.37343, -52.33518, -52.32457, -52.29548, -52.27136, -52.29337, 
    -52.31649, -52.38231, -52.44169, -52.50649, -52.52243, -52.59803, 
    -52.53635, -52.63805, -52.5514, -52.70162, -52.43227, -52.54899, 
    -52.33784, -52.36057, -52.40162, -52.49605, -52.44516, -52.50473, 
    -52.37309, -52.30482, -52.28727, -52.25433, -52.28802, -52.2853, 
    -52.3175, -52.30716, -52.38451, -52.34296, -52.46114, -52.5043, 
    -52.62652, -52.70152, -52.77813, -52.81194, -52.82223, -52.82654 ;

 FGR_R =
  -396.58, -397.6065, -397.4086, -398.23, -397.7746, -398.3122, -396.7943, 
    -397.6467, -397.1028, -396.6721, -399.8222, -398.2667, -401.4498, 
    -400.4582, -402.9492, -401.2952, -403.2826, -402.9022, -404.0486, 
    -403.7203, -405.1845, -404.2002, -405.9441, -404.9499, -405.1052, 
    -404.1676, -398.5805, -399.6284, -398.5182, -398.6677, -398.6008, 
    -397.7838, -397.3716, -396.5025, -396.6591, -397.2996, -398.735, 
    -398.2483, -399.476, -399.4483, -400.824, -400.1982, -402.5027, -401.851, 
    -403.734, -403.2606, -403.7117, -403.575, -403.7135, -403.0191, 
    -403.3166, -402.7056, -400.3134, -401.0237, -398.9243, -397.6661, 
    -396.8316, -396.2314, -396.3152, -396.4748, -397.3033, -398.0755, 
    -398.6636, -399.0568, -399.4443, -400.6251, -401.2459, -402.6341, 
    -402.3842, -402.808, -403.2135, -403.8933, -403.7816, -404.0809, 
    -402.7972, -403.6502, -402.2417, -402.627, -399.5473, -398.3797, 
    -397.8813, -397.4466, -396.3795, -397.1186, -396.8302, -397.5168, 
    -397.9527, -397.7372, -399.0676, -398.5504, -401.2827, -400.1004, 
    -403.1662, -402.4356, -403.3414, -402.8793, -403.6707, -402.9585, 
    -404.1925, -404.4608, -404.2774, -404.9825, -402.9189, -403.7115, 
    -397.7311, -397.7662, -397.9301, -397.2095, -397.1655, -396.4981, 
    -397.093, -397.3429, -397.9782, -398.3534, -398.7102, -399.4945, 
    -400.3697, -401.6038, -402.4829, -403.0719, -402.7109, -403.0296, 
    -402.6732, -402.5063, -404.3601, -403.3192, -404.8811, -404.7948, 
    -404.0879, -404.8046, -397.7909, -397.5887, -396.8857, -397.4359, 
    -396.4262, -396.9944, -397.3166, -398.5607, -398.8345, -399.0876, 
    -399.588, -400.2297, -401.365, -402.3438, -403.2372, -403.1718, 
    -403.1948, -403.3941, -402.9001, -403.4752, -403.5715, -403.3194, 
    -404.7833, -404.3652, -404.793, -404.5209, -397.6545, -397.9949, 
    -397.8109, -398.1567, -397.9129, -398.996, -399.3207, -400.8498, 
    -400.2169, -401.2187, -400.3178, -400.4857, -401.2501, -400.3763, 
    -402.2894, -400.9918, -403.4018, -402.1059, -403.4829, -403.2333, 
    -403.6468, -404.0168, -404.4827, -405.3412, -405.1425, -405.8606, 
    -398.5024, -398.9435, -398.9051, -399.3669, -399.7083, -400.4587, 
    -401.645, -401.1991, -402.0181, -402.1823, -400.9384, -401.7018, 
    -399.239, -399.635, -399.3995, -398.537, -401.3013, -399.8779, -402.4973, 
    -401.7324, -403.964, -402.8541, -405.033, -405.9625, -406.8388, -407.86, 
    -399.1847, -398.8849, -399.422, -400.1639, -400.8635, -401.779, 
    -401.8729, -402.0442, -402.4885, -402.8617, -402.098, -402.9553, 
    -399.726, -401.4241, -398.7712, -399.5668, -400.1204, -399.878, 
    -401.1483, -401.445, -402.6502, -402.0275, -405.7328, -404.0944, 
    -408.6385, -407.3696, -398.7801, -399.1838, -400.5979, -399.9199, 
    -401.8403, -402.3101, -402.6922, -403.1799, -403.2328, -403.5218, 
    -403.0482, -403.5032, -401.781, -402.5509, -400.438, -400.9522, 
    -400.7158, -400.4561, -401.2574, -402.1099, -402.1288, -402.4019, 
    -403.1703, -401.8481, -405.9428, -403.414, -399.6239, -400.4104, 
    -400.5221, -400.2111, -402.2629, -401.5233, -403.5148, -402.977, 
    -403.8583, -403.4203, -403.3559, -402.7933, -402.4428, -401.5571, 
    -400.8364, -400.2548, -400.3979, -401.0255, -402.1622, -403.2373, 
    -403.0018, -403.7914, -401.7019, -402.578, -402.2392, -403.1226, 
    -401.1871, -402.8333, -400.7659, -400.9474, -401.5087, -402.6369, 
    -402.8875, -403.1537, -402.9896, -402.1912, -402.0606, -401.4952, 
    -401.3387, -400.9079, -400.5509, -400.8769, -401.2191, -402.1918, 
    -403.0675, -404.022, -404.2558, -405.3685, -404.4618, -405.9568, 
    -404.6844, -406.887, -402.9297, -404.6484, -401.5345, -401.8703, 
    -402.477, -403.8691, -403.1184, -403.9966, -402.0556, -401.0468, 
    -400.7866, -400.2894, -400.7978, -400.7573, -401.2338, -401.0807, 
    -402.2241, -401.61, -403.3541, -403.9899, -405.7851, -406.8842, 
    -408.0034, -408.4968, -408.647, -408.7098 ;

 FGR_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FIRA =
  48.64412, 48.71832, 48.70387, 48.76385, 48.7306, 48.76985, 48.65901, 
    48.72125, 48.68153, 48.65086, 48.88011, 48.76653, 48.99666, 48.92426, 
    49.10614, 48.98536, 49.1305, 49.10272, 49.18645, 49.16247, 49.26938, 
    49.19751, 49.32486, 49.25225, 49.26359, 49.19513, 48.78945, 48.86595, 
    48.7849, 48.79582, 48.79093, 48.73127, 48.70115, 48.63847, 48.6499, 
    48.6959, 48.80073, 48.76519, 48.85485, 48.85283, 48.95097, 48.9076, 
    49.07355, 49.02597, 49.16347, 49.1289, 49.16184, 49.15186, 49.16197, 
    49.11126, 49.13298, 49.08837, 48.916, 48.96555, 48.81456, 48.72265, 
    48.66173, 48.61866, 48.62479, 48.63644, 48.69617, 48.75257, 48.79552, 
    48.82424, 48.85254, 48.93643, 48.98177, 49.08314, 49.0649, 49.09584, 
    49.12546, 49.17511, 49.16694, 49.1888, 49.09506, 49.15735, 49.0545, 
    49.08263, 48.86003, 48.77479, 48.73837, 48.70664, 48.62949, 48.68269, 
    48.66162, 48.71177, 48.7436, 48.72787, 48.82502, 48.78725, 48.98446, 
    48.90045, 49.12201, 49.06865, 49.1348, 49.10106, 49.15885, 49.10684, 
    49.19695, 49.21654, 49.20315, 49.25465, 49.10395, 49.16182, 48.72742, 
    48.72998, 48.74196, 48.68932, 48.68611, 48.63815, 48.68082, 48.69907, 
    48.74546, 48.77287, 48.79892, 48.8562, 48.92011, 49.0079, 49.07211, 
    49.11512, 49.08876, 49.11203, 49.08601, 49.07382, 49.20919, 49.13317, 
    49.24724, 49.24094, 49.18931, 49.24165, 48.73179, 48.71702, 48.66568, 
    48.70586, 48.6329, 48.67362, 48.69714, 48.788, 48.808, 48.82648, 
    48.86303, 48.90989, 48.99047, 49.06195, 49.12719, 49.12241, 49.1241, 
    49.13865, 49.10257, 49.14457, 49.1516, 49.13319, 49.24009, 49.20956, 
    49.24081, 49.22093, 48.72183, 48.74669, 48.73325, 48.7585, 48.7407, 
    48.81979, 48.84349, 48.95285, 48.90896, 48.97979, 48.91634, 48.92627, 
    48.98207, 48.91829, 49.05797, 48.96321, 49.13921, 49.04456, 49.14513, 
    49.12691, 49.1571, 49.18412, 49.21814, 49.28083, 49.26632, 49.31876, 
    48.78375, 48.81596, 48.81316, 48.84689, 48.87181, 48.9243, 49.01092, 
    48.97837, 49.03817, 49.05016, 48.95933, 49.01506, 48.83754, 48.86645, 
    48.84927, 48.78627, 48.98582, 48.88419, 49.07316, 49.01731, 49.18026, 
    49.09921, 49.25833, 49.32619, 49.39021, 49.46478, 48.83357, 48.81169, 
    48.85091, 48.90508, 48.95386, 49.02071, 49.02757, 49.04007, 49.07252, 
    49.09977, 49.04399, 49.1066, 48.87308, 48.99479, 48.80338, 48.86147, 
    48.90191, 48.8842, 48.97466, 48.99632, 49.08432, 49.03886, 49.30941, 
    49.18978, 49.52164, 49.42897, 48.80403, 48.83352, 48.93446, 48.88727, 
    49.02519, 49.05949, 49.08739, 49.123, 49.12687, 49.14797, 49.11339, 
    49.14662, 49.02085, 49.07707, 48.92279, 48.96033, 48.94308, 48.92412, 
    48.98262, 49.04486, 49.04625, 49.06619, 49.12226, 49.02576, 49.32474, 
    49.14006, 48.86566, 48.92076, 48.92893, 48.90854, 49.05605, 49.00204, 
    49.14746, 49.10819, 49.17255, 49.14056, 49.13586, 49.09478, 49.06918, 
    49.00451, 48.95188, 48.91174, 48.91987, 48.96569, 49.04868, 49.12719, 
    49.10999, 49.16766, 49.01508, 49.07904, 49.05431, 49.11882, 48.97749, 
    49.09766, 48.94674, 48.95999, 49.00097, 49.08334, 49.10165, 49.12109, 
    49.10911, 49.0508, 49.04127, 48.99999, 48.98856, 48.95711, 48.93103, 
    48.95484, 48.97982, 49.05085, 49.11479, 49.1845, 49.20158, 49.28281, 
    49.2166, 49.32575, 49.23283, 49.3937, 49.10471, 49.23022, 49.00285, 
    49.02738, 49.07167, 49.17332, 49.11852, 49.18264, 49.0409, 48.96724, 
    48.94825, 48.91426, 48.94906, 48.94611, 48.9809, 48.96972, 49.05321, 
    49.00837, 49.13572, 49.18215, 49.31325, 49.39351, 49.47526, 49.5113, 
    49.52227, 49.52686 ;

 FIRA_R =
  48.64412, 48.71832, 48.70387, 48.76385, 48.7306, 48.76985, 48.65901, 
    48.72125, 48.68153, 48.65086, 48.88011, 48.76653, 48.99666, 48.92426, 
    49.10614, 48.98536, 49.1305, 49.10272, 49.18645, 49.16247, 49.26938, 
    49.19751, 49.32486, 49.25225, 49.26359, 49.19513, 48.78945, 48.86595, 
    48.7849, 48.79582, 48.79093, 48.73127, 48.70115, 48.63847, 48.6499, 
    48.6959, 48.80073, 48.76519, 48.85485, 48.85283, 48.95097, 48.9076, 
    49.07355, 49.02597, 49.16347, 49.1289, 49.16184, 49.15186, 49.16197, 
    49.11126, 49.13298, 49.08837, 48.916, 48.96555, 48.81456, 48.72265, 
    48.66173, 48.61866, 48.62479, 48.63644, 48.69617, 48.75257, 48.79552, 
    48.82424, 48.85254, 48.93643, 48.98177, 49.08314, 49.0649, 49.09584, 
    49.12546, 49.17511, 49.16694, 49.1888, 49.09506, 49.15735, 49.0545, 
    49.08263, 48.86003, 48.77479, 48.73837, 48.70664, 48.62949, 48.68269, 
    48.66162, 48.71177, 48.7436, 48.72787, 48.82502, 48.78725, 48.98446, 
    48.90045, 49.12201, 49.06865, 49.1348, 49.10106, 49.15885, 49.10684, 
    49.19695, 49.21654, 49.20315, 49.25465, 49.10395, 49.16182, 48.72742, 
    48.72998, 48.74196, 48.68932, 48.68611, 48.63815, 48.68082, 48.69907, 
    48.74546, 48.77287, 48.79892, 48.8562, 48.92011, 49.0079, 49.07211, 
    49.11512, 49.08876, 49.11203, 49.08601, 49.07382, 49.20919, 49.13317, 
    49.24724, 49.24094, 49.18931, 49.24165, 48.73179, 48.71702, 48.66568, 
    48.70586, 48.6329, 48.67362, 48.69714, 48.788, 48.808, 48.82648, 
    48.86303, 48.90989, 48.99047, 49.06195, 49.12719, 49.12241, 49.1241, 
    49.13865, 49.10257, 49.14457, 49.1516, 49.13319, 49.24009, 49.20956, 
    49.24081, 49.22093, 48.72183, 48.74669, 48.73325, 48.7585, 48.7407, 
    48.81979, 48.84349, 48.95285, 48.90896, 48.97979, 48.91634, 48.92627, 
    48.98207, 48.91829, 49.05797, 48.96321, 49.13921, 49.04456, 49.14513, 
    49.12691, 49.1571, 49.18412, 49.21814, 49.28083, 49.26632, 49.31876, 
    48.78375, 48.81596, 48.81316, 48.84689, 48.87181, 48.9243, 49.01092, 
    48.97837, 49.03817, 49.05016, 48.95933, 49.01506, 48.83754, 48.86645, 
    48.84927, 48.78627, 48.98582, 48.88419, 49.07316, 49.01731, 49.18026, 
    49.09921, 49.25833, 49.32619, 49.39021, 49.46478, 48.83357, 48.81169, 
    48.85091, 48.90508, 48.95386, 49.02071, 49.02757, 49.04007, 49.07252, 
    49.09977, 49.04399, 49.1066, 48.87308, 48.99479, 48.80338, 48.86147, 
    48.90191, 48.8842, 48.97466, 48.99632, 49.08432, 49.03886, 49.30941, 
    49.18978, 49.52164, 49.42897, 48.80403, 48.83352, 48.93446, 48.88727, 
    49.02519, 49.05949, 49.08739, 49.123, 49.12687, 49.14797, 49.11339, 
    49.14662, 49.02085, 49.07707, 48.92279, 48.96033, 48.94308, 48.92412, 
    48.98262, 49.04486, 49.04625, 49.06619, 49.12226, 49.02576, 49.32474, 
    49.14006, 48.86566, 48.92076, 48.92893, 48.90854, 49.05605, 49.00204, 
    49.14746, 49.10819, 49.17255, 49.14056, 49.13586, 49.09478, 49.06918, 
    49.00451, 48.95188, 48.91174, 48.91987, 48.96569, 49.04868, 49.12719, 
    49.10999, 49.16766, 49.01508, 49.07904, 49.05431, 49.11882, 48.97749, 
    49.09766, 48.94674, 48.95999, 49.00097, 49.08334, 49.10165, 49.12109, 
    49.10911, 49.0508, 49.04127, 48.99999, 48.98856, 48.95711, 48.93103, 
    48.95484, 48.97982, 49.05085, 49.11479, 49.1845, 49.20158, 49.28281, 
    49.2166, 49.32575, 49.23283, 49.3937, 49.10471, 49.23022, 49.00285, 
    49.02738, 49.07167, 49.17332, 49.11852, 49.18264, 49.0409, 48.96724, 
    48.94825, 48.91426, 48.94906, 48.94611, 48.9809, 48.96972, 49.05321, 
    49.00837, 49.13572, 49.18215, 49.31325, 49.39351, 49.47526, 49.5113, 
    49.52227, 49.52686 ;

 FIRA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FIRE =
  262.9903, 263.0645, 263.05, 263.11, 263.0768, 263.116, 263.0052, 263.0674, 
    263.0277, 262.997, 263.2263, 263.1127, 263.3428, 263.2704, 263.4523, 
    263.3315, 263.4767, 263.4489, 263.5326, 263.5086, 263.6155, 263.5437, 
    263.671, 263.5984, 263.6097, 263.5413, 263.1356, 263.2121, 263.131, 
    263.142, 263.1371, 263.0774, 263.0473, 262.9846, 262.996, 263.0421, 
    263.1469, 263.1113, 263.201, 263.199, 263.2971, 263.2538, 263.4197, 
    263.3721, 263.5096, 263.475, 263.508, 263.498, 263.5081, 263.4574, 
    263.4791, 263.4345, 263.2621, 263.3117, 263.1607, 263.0688, 263.0079, 
    262.9648, 262.9709, 262.9826, 263.0423, 263.0987, 263.1417, 263.1704, 
    263.1987, 263.2826, 263.3279, 263.4293, 263.411, 263.442, 263.4716, 
    263.5212, 263.5131, 263.5349, 263.4412, 263.5035, 263.4006, 263.4288, 
    263.2062, 263.1209, 263.0845, 263.0528, 262.9756, 263.0288, 263.0078, 
    263.0579, 263.0898, 263.074, 263.1712, 263.1334, 263.3306, 263.2466, 
    263.4681, 263.4148, 263.4809, 263.4472, 263.505, 263.453, 263.5431, 
    263.5627, 263.5493, 263.6008, 263.4501, 263.508, 263.0736, 263.0761, 
    263.0881, 263.0355, 263.0323, 262.9843, 263.0269, 263.0452, 263.0916, 
    263.119, 263.1451, 263.2023, 263.2663, 263.354, 263.4182, 263.4613, 
    263.4349, 263.4582, 263.4322, 263.42, 263.5553, 263.4793, 263.5934, 
    263.5871, 263.5355, 263.5878, 263.0779, 263.0632, 263.0118, 263.052, 
    262.979, 263.0198, 263.0433, 263.1342, 263.1541, 263.1726, 263.2092, 
    263.256, 263.3366, 263.4081, 263.4733, 263.4686, 263.4702, 263.4848, 
    263.4487, 263.4907, 263.4977, 263.4793, 263.5862, 263.5557, 263.5869, 
    263.5671, 263.068, 263.0928, 263.0794, 263.1046, 263.0869, 263.1659, 
    263.1896, 263.299, 263.2551, 263.3259, 263.2625, 263.2724, 263.3282, 
    263.2644, 263.4041, 263.3094, 263.4854, 263.3907, 263.4913, 263.4731, 
    263.5032, 263.5303, 263.5643, 263.627, 263.6125, 263.6649, 263.1299, 
    263.1621, 263.1593, 263.193, 263.218, 263.2704, 263.3571, 263.3245, 
    263.3843, 263.3963, 263.3055, 263.3612, 263.1837, 263.2126, 263.1954, 
    263.1324, 263.332, 263.2303, 263.4193, 263.3635, 263.5264, 263.4453, 
    263.6045, 263.6723, 263.7364, 263.8109, 263.1797, 263.1578, 263.1971, 
    263.2512, 263.3, 263.3669, 263.3737, 263.3862, 263.4187, 263.4459, 
    263.3901, 263.4528, 263.2192, 263.3409, 263.1495, 263.2076, 263.248, 
    263.2303, 263.3208, 263.3425, 263.4305, 263.385, 263.6555, 263.5359, 
    263.8678, 263.7751, 263.1502, 263.1797, 263.2806, 263.2334, 263.3713, 
    263.4056, 263.4335, 263.4691, 263.473, 263.4941, 263.4595, 263.4928, 
    263.367, 263.4232, 263.2689, 263.3065, 263.2892, 263.2703, 263.3288, 
    263.391, 263.3924, 263.4123, 263.4684, 263.3719, 263.6709, 263.4862, 
    263.2118, 263.2669, 263.2751, 263.2547, 263.4022, 263.3482, 263.4936, 
    263.4543, 263.5187, 263.4867, 263.482, 263.4409, 263.4153, 263.3506, 
    263.298, 263.2579, 263.266, 263.3118, 263.3948, 263.4733, 263.4561, 
    263.5138, 263.3612, 263.4252, 263.4005, 263.465, 263.3236, 263.4438, 
    263.2929, 263.3061, 263.3471, 263.4295, 263.4478, 263.4672, 263.4553, 
    263.3969, 263.3874, 263.3461, 263.3347, 263.3033, 263.2772, 263.301, 
    263.326, 263.397, 263.4609, 263.5306, 263.5477, 263.6289, 263.5627, 
    263.6719, 263.579, 263.7398, 263.4509, 263.5764, 263.349, 263.3735, 
    263.4178, 263.5195, 263.4647, 263.5288, 263.3871, 263.3134, 263.2944, 
    263.2604, 263.2952, 263.2922, 263.3271, 263.3159, 263.3994, 263.3545, 
    263.4819, 263.5283, 263.6594, 263.7397, 263.8214, 263.8575, 263.8684, 
    263.873 ;

 FIRE_R =
  262.9903, 263.0645, 263.05, 263.11, 263.0768, 263.116, 263.0052, 263.0674, 
    263.0277, 262.997, 263.2263, 263.1127, 263.3428, 263.2704, 263.4523, 
    263.3315, 263.4767, 263.4489, 263.5326, 263.5086, 263.6155, 263.5437, 
    263.671, 263.5984, 263.6097, 263.5413, 263.1356, 263.2121, 263.131, 
    263.142, 263.1371, 263.0774, 263.0473, 262.9846, 262.996, 263.0421, 
    263.1469, 263.1113, 263.201, 263.199, 263.2971, 263.2538, 263.4197, 
    263.3721, 263.5096, 263.475, 263.508, 263.498, 263.5081, 263.4574, 
    263.4791, 263.4345, 263.2621, 263.3117, 263.1607, 263.0688, 263.0079, 
    262.9648, 262.9709, 262.9826, 263.0423, 263.0987, 263.1417, 263.1704, 
    263.1987, 263.2826, 263.3279, 263.4293, 263.411, 263.442, 263.4716, 
    263.5212, 263.5131, 263.5349, 263.4412, 263.5035, 263.4006, 263.4288, 
    263.2062, 263.1209, 263.0845, 263.0528, 262.9756, 263.0288, 263.0078, 
    263.0579, 263.0898, 263.074, 263.1712, 263.1334, 263.3306, 263.2466, 
    263.4681, 263.4148, 263.4809, 263.4472, 263.505, 263.453, 263.5431, 
    263.5627, 263.5493, 263.6008, 263.4501, 263.508, 263.0736, 263.0761, 
    263.0881, 263.0355, 263.0323, 262.9843, 263.0269, 263.0452, 263.0916, 
    263.119, 263.1451, 263.2023, 263.2663, 263.354, 263.4182, 263.4613, 
    263.4349, 263.4582, 263.4322, 263.42, 263.5553, 263.4793, 263.5934, 
    263.5871, 263.5355, 263.5878, 263.0779, 263.0632, 263.0118, 263.052, 
    262.979, 263.0198, 263.0433, 263.1342, 263.1541, 263.1726, 263.2092, 
    263.256, 263.3366, 263.4081, 263.4733, 263.4686, 263.4702, 263.4848, 
    263.4487, 263.4907, 263.4977, 263.4793, 263.5862, 263.5557, 263.5869, 
    263.5671, 263.068, 263.0928, 263.0794, 263.1046, 263.0869, 263.1659, 
    263.1896, 263.299, 263.2551, 263.3259, 263.2625, 263.2724, 263.3282, 
    263.2644, 263.4041, 263.3094, 263.4854, 263.3907, 263.4913, 263.4731, 
    263.5032, 263.5303, 263.5643, 263.627, 263.6125, 263.6649, 263.1299, 
    263.1621, 263.1593, 263.193, 263.218, 263.2704, 263.3571, 263.3245, 
    263.3843, 263.3963, 263.3055, 263.3612, 263.1837, 263.2126, 263.1954, 
    263.1324, 263.332, 263.2303, 263.4193, 263.3635, 263.5264, 263.4453, 
    263.6045, 263.6723, 263.7364, 263.8109, 263.1797, 263.1578, 263.1971, 
    263.2512, 263.3, 263.3669, 263.3737, 263.3862, 263.4187, 263.4459, 
    263.3901, 263.4528, 263.2192, 263.3409, 263.1495, 263.2076, 263.248, 
    263.2303, 263.3208, 263.3425, 263.4305, 263.385, 263.6555, 263.5359, 
    263.8678, 263.7751, 263.1502, 263.1797, 263.2806, 263.2334, 263.3713, 
    263.4056, 263.4335, 263.4691, 263.473, 263.4941, 263.4595, 263.4928, 
    263.367, 263.4232, 263.2689, 263.3065, 263.2892, 263.2703, 263.3288, 
    263.391, 263.3924, 263.4123, 263.4684, 263.3719, 263.6709, 263.4862, 
    263.2118, 263.2669, 263.2751, 263.2547, 263.4022, 263.3482, 263.4936, 
    263.4543, 263.5187, 263.4867, 263.482, 263.4409, 263.4153, 263.3506, 
    263.298, 263.2579, 263.266, 263.3118, 263.3948, 263.4733, 263.4561, 
    263.5138, 263.3612, 263.4252, 263.4005, 263.465, 263.3236, 263.4438, 
    263.2929, 263.3061, 263.3471, 263.4295, 263.4478, 263.4672, 263.4553, 
    263.3969, 263.3874, 263.3461, 263.3347, 263.3033, 263.2772, 263.301, 
    263.326, 263.397, 263.4609, 263.5306, 263.5477, 263.6289, 263.5627, 
    263.6719, 263.579, 263.7398, 263.4509, 263.5764, 263.349, 263.3735, 
    263.4178, 263.5195, 263.4647, 263.5288, 263.3871, 263.3134, 263.2944, 
    263.2604, 263.2952, 263.2922, 263.3271, 263.3159, 263.3994, 263.3545, 
    263.4819, 263.5283, 263.6594, 263.7397, 263.8214, 263.8575, 263.8684, 
    263.873 ;

 FIRE_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FLDS =
  214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461 ;

 FPG =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI_vr =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WJ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROST_TABLE =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 FSA =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 FSAT =
  0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584 ;

 FSA_R =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 FSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSDS =
  1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347 ;

 FSDSND =
  0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532 ;

 FSDSNDLN =
  0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495 ;

 FSDSNI =
  0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819 ;

 FSDSVD =
  0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128 ;

 FSDSVDLN =
  0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609 ;

 FSDSVI =
  0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223 ;

 FSDSVILN =
  0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376 ;

 FSH =
  347.9881, 348.9405, 348.757, 349.5184, 349.0963, 349.5947, 348.1876, 
    348.9778, 348.4735, 348.0735, 350.9944, 349.5525, 352.5055, 351.5862, 
    353.8953, 352.3621, 354.2044, 353.8517, 354.9145, 354.6101, 355.9674, 
    355.055, 356.6715, 355.7499, 355.8939, 355.0247, 349.8433, 350.8148, 
    349.7856, 349.9242, 349.8622, 349.1048, 348.7227, 347.9163, 348.0615, 
    348.6559, 349.9865, 349.5354, 350.6734, 350.6477, 351.9253, 351.3429, 
    353.4814, 352.8774, 354.6229, 354.184, 354.6021, 354.4754, 354.6038, 
    353.9601, 354.2359, 353.6696, 351.4496, 352.1104, 350.162, 348.9957, 
    348.2221, 347.665, 347.7427, 347.8907, 348.6594, 349.3752, 349.9204, 
    350.2849, 350.644, 351.7409, 352.3164, 353.6032, 353.3716, 353.7644, 
    354.1403, 354.7705, 354.6669, 354.9444, 353.7544, 354.5452, 353.2395, 
    353.5967, 350.7396, 349.6572, 349.1952, 348.7922, 347.8024, 348.4882, 
    348.2208, 348.8574, 349.2614, 349.0617, 350.2949, 349.8154, 352.3505, 
    351.2523, 354.0965, 353.4192, 354.2589, 353.8306, 354.5642, 353.904, 
    355.0478, 355.2965, 355.1265, 355.7802, 353.8673, 354.6019, 349.056, 
    349.0885, 349.2405, 348.5724, 348.5317, 347.9122, 348.4644, 348.6961, 
    349.285, 349.6328, 349.9636, 350.6906, 351.5018, 352.6481, 353.4631, 
    354.009, 353.6744, 353.9698, 353.6395, 353.4848, 355.2032, 354.2383, 
    355.6862, 355.6062, 354.9509, 355.6152, 349.1115, 348.924, 348.2723, 
    348.7823, 347.8456, 348.3731, 348.6718, 349.825, 350.0788, 350.3134, 
    350.7773, 351.3721, 352.4268, 353.3341, 354.1623, 354.1017, 354.123, 
    354.3077, 353.8498, 354.3829, 354.4722, 354.2385, 355.5955, 355.2079, 
    355.6045, 355.3522, 348.985, 349.3005, 349.13, 349.4505, 349.2245, 
    350.2285, 350.5295, 351.9493, 351.3603, 352.2912, 351.4538, 351.6118, 
    352.3203, 351.5103, 353.2837, 352.0808, 354.3149, 353.1136, 354.3901, 
    354.1587, 354.542, 354.885, 355.3168, 356.1126, 355.9285, 356.5941, 
    349.771, 350.1798, 350.1442, 350.5723, 350.8888, 351.5867, 352.6864, 
    352.2731, 353.0322, 353.1844, 352.0313, 352.739, 350.4537, 350.8208, 
    350.6026, 349.803, 352.3678, 351.046, 353.4765, 352.7674, 354.8361, 
    353.8072, 355.827, 356.6886, 357.5009, 358.4475, 350.4034, 350.1255, 
    350.6234, 351.3111, 351.9619, 352.8106, 352.8976, 353.0564, 353.4682, 
    353.8142, 353.1063, 353.9009, 350.9052, 352.4816, 350.0201, 350.7576, 
    351.2708, 351.0461, 352.2259, 352.501, 353.6182, 353.041, 356.4756, 
    354.9569, 359.1691, 357.993, 350.0284, 350.4026, 351.7157, 351.0849, 
    352.8674, 353.3029, 353.6571, 354.1092, 354.1583, 354.4261, 353.9871, 
    354.4089, 352.8124, 353.5261, 351.5674, 352.0441, 351.825, 351.5843, 
    352.327, 353.1173, 353.1348, 353.3881, 354.1003, 352.8746, 356.6704, 
    354.3262, 350.8106, 351.5419, 351.6455, 351.3549, 353.2592, 352.5736, 
    354.4196, 353.9211, 354.7381, 354.3321, 354.2723, 353.7509, 353.4259, 
    352.6049, 351.9368, 351.3954, 351.5303, 352.1122, 353.1658, 354.1624, 
    353.9441, 354.676, 352.7391, 353.5512, 353.2372, 354.056, 352.2619, 
    353.7879, 351.8714, 352.0397, 352.56, 353.6059, 353.8381, 354.0849, 
    353.9327, 353.1927, 353.0717, 352.5475, 352.4024, 352.0031, 351.6721, 
    351.9744, 352.2916, 353.1932, 354.005, 354.8898, 355.1065, 356.138, 
    355.2975, 356.6833, 355.5039, 357.5456, 353.8773, 355.4705, 352.5839, 
    352.8953, 353.4576, 354.7481, 354.0522, 354.8663, 353.067, 352.1319, 
    351.8907, 351.4275, 351.901, 351.8635, 352.3052, 352.1633, 353.2232, 
    352.654, 354.2706, 354.86, 356.5241, 357.543, 358.5804, 359.0378, 
    359.1771, 359.2352 ;

 FSH_G =
  354.7173, 355.6701, 355.4866, 356.2484, 355.826, 356.3247, 354.9168, 
    355.7074, 355.2029, 354.8027, 357.7251, 356.2824, 359.237, 358.3173, 
    360.6276, 359.0936, 360.9369, 360.584, 361.6474, 361.3429, 362.7009, 
    361.7879, 363.4054, 362.4832, 362.6273, 361.7577, 356.5735, 357.5454, 
    356.5157, 356.6544, 356.5923, 355.8346, 355.4522, 354.6454, 354.7906, 
    355.3854, 356.7167, 356.2654, 357.404, 357.3783, 358.6566, 358.0739, 
    360.2135, 359.6092, 361.3556, 360.9165, 361.3349, 361.2081, 361.3365, 
    360.6925, 360.9684, 360.4018, 358.1807, 358.8418, 356.8923, 355.7254, 
    354.9514, 354.3939, 354.4716, 354.6197, 355.3889, 356.1051, 356.6506, 
    357.0153, 357.3746, 358.4721, 359.0479, 360.3354, 360.1037, 360.4967, 
    360.8728, 361.5034, 361.3997, 361.6773, 360.4867, 361.2779, 359.9715, 
    360.3289, 357.4702, 356.3872, 355.9249, 355.5218, 354.5314, 355.2176, 
    354.9501, 355.5869, 355.9912, 355.7914, 357.0252, 356.5456, 359.082, 
    357.9832, 360.8289, 360.1513, 360.9914, 360.5629, 361.2969, 360.6363, 
    361.7808, 362.0296, 361.8595, 362.5136, 360.5996, 361.3347, 355.7857, 
    355.8183, 355.9703, 355.3019, 355.2611, 354.6413, 355.1938, 355.4256, 
    356.0148, 356.3629, 356.6938, 357.4212, 358.2329, 359.3798, 360.1952, 
    360.7415, 360.4066, 360.7022, 360.3717, 360.2169, 361.9362, 360.9709, 
    362.4195, 362.3395, 361.6838, 362.3485, 355.8412, 355.6536, 355.0016, 
    355.5119, 354.5747, 355.1024, 355.4013, 356.5551, 356.8091, 357.0438, 
    357.5079, 358.1031, 359.1584, 360.0662, 360.8948, 360.8341, 360.8554, 
    361.0403, 360.5821, 361.1155, 361.2048, 360.971, 362.3287, 361.941, 
    362.3378, 362.0854, 355.7146, 356.0303, 355.8597, 356.1804, 355.9543, 
    356.9589, 357.2599, 358.6805, 358.0912, 359.0227, 358.1848, 358.3429, 
    359.0518, 358.2414, 360.0157, 358.8122, 361.0475, 359.8455, 361.1227, 
    360.8912, 361.2747, 361.6179, 362.0499, 362.8462, 362.6619, 363.3279, 
    356.5011, 356.9102, 356.8745, 357.3029, 357.6195, 358.3178, 359.418, 
    359.0045, 359.7641, 359.9164, 358.7626, 359.4707, 357.1842, 357.5515, 
    357.3331, 356.5331, 359.0993, 357.7767, 360.2086, 359.4991, 361.5689, 
    360.5395, 362.5604, 363.4225, 364.2353, 365.1823, 357.1338, 356.8558, 
    357.3539, 358.042, 358.6932, 359.5423, 359.6294, 359.7883, 360.2003, 
    360.5465, 359.8382, 360.6333, 357.6359, 359.2132, 356.7504, 357.4882, 
    358.0016, 357.7768, 358.9573, 359.2326, 360.3503, 359.7729, 363.2094, 
    361.6898, 365.9044, 364.7275, 356.7586, 357.1331, 358.4468, 357.8157, 
    359.5992, 360.0349, 360.3893, 360.8416, 360.8907, 361.1587, 360.7195, 
    361.1415, 359.5442, 360.2582, 358.2985, 358.7755, 358.5562, 358.3154, 
    359.0585, 359.8492, 359.8668, 360.1201, 360.8327, 359.6064, 363.4042, 
    361.0587, 357.5412, 358.273, 358.3766, 358.0858, 359.9912, 359.3052, 
    361.1523, 360.6534, 361.4709, 361.0647, 361.0049, 360.4831, 360.158, 
    359.3365, 358.6681, 358.1263, 358.2614, 358.8435, 359.8977, 360.8949, 
    360.6764, 361.4088, 359.4708, 360.2834, 359.9691, 360.7885, 358.9934, 
    360.5202, 358.6027, 358.771, 359.2916, 360.338, 360.5704, 360.8173, 
    360.6651, 359.9246, 359.8035, 359.2791, 359.134, 358.7344, 358.4033, 
    358.7057, 359.0231, 359.9252, 360.7374, 361.6227, 361.8395, 362.8715, 
    362.0306, 363.4171, 362.2371, 364.2799, 360.6096, 362.2036, 359.3155, 
    359.627, 360.1897, 361.4809, 360.7846, 361.5992, 359.7989, 358.8633, 
    358.6219, 358.1584, 358.6322, 358.5947, 359.0367, 358.8947, 359.9551, 
    359.3856, 361.0032, 361.5929, 363.2579, 364.2773, 365.3153, 365.773, 
    365.9123, 365.9705 ;

 FSH_NODYNLNDUSE =
  347.9881, 348.9405, 348.757, 349.5184, 349.0963, 349.5947, 348.1876, 
    348.9778, 348.4735, 348.0735, 350.9944, 349.5525, 352.5055, 351.5862, 
    353.8953, 352.3621, 354.2044, 353.8517, 354.9145, 354.6101, 355.9674, 
    355.055, 356.6715, 355.7499, 355.8939, 355.0247, 349.8433, 350.8148, 
    349.7856, 349.9242, 349.8622, 349.1048, 348.7227, 347.9163, 348.0615, 
    348.6559, 349.9865, 349.5354, 350.6734, 350.6477, 351.9253, 351.3429, 
    353.4814, 352.8774, 354.6229, 354.184, 354.6021, 354.4754, 354.6038, 
    353.9601, 354.2359, 353.6696, 351.4496, 352.1104, 350.162, 348.9957, 
    348.2221, 347.665, 347.7427, 347.8907, 348.6594, 349.3752, 349.9204, 
    350.2849, 350.644, 351.7409, 352.3164, 353.6032, 353.3716, 353.7644, 
    354.1403, 354.7705, 354.6669, 354.9444, 353.7544, 354.5452, 353.2395, 
    353.5967, 350.7396, 349.6572, 349.1952, 348.7922, 347.8024, 348.4882, 
    348.2208, 348.8574, 349.2614, 349.0617, 350.2949, 349.8154, 352.3505, 
    351.2523, 354.0965, 353.4192, 354.2589, 353.8306, 354.5642, 353.904, 
    355.0478, 355.2965, 355.1265, 355.7802, 353.8673, 354.6019, 349.056, 
    349.0885, 349.2405, 348.5724, 348.5317, 347.9122, 348.4644, 348.6961, 
    349.285, 349.6328, 349.9636, 350.6906, 351.5018, 352.6481, 353.4631, 
    354.009, 353.6744, 353.9698, 353.6395, 353.4848, 355.2032, 354.2383, 
    355.6862, 355.6062, 354.9509, 355.6152, 349.1115, 348.924, 348.2723, 
    348.7823, 347.8456, 348.3731, 348.6718, 349.825, 350.0788, 350.3134, 
    350.7773, 351.3721, 352.4268, 353.3341, 354.1623, 354.1017, 354.123, 
    354.3077, 353.8498, 354.3829, 354.4722, 354.2385, 355.5955, 355.2079, 
    355.6045, 355.3522, 348.985, 349.3005, 349.13, 349.4505, 349.2245, 
    350.2285, 350.5295, 351.9493, 351.3603, 352.2912, 351.4538, 351.6118, 
    352.3203, 351.5103, 353.2837, 352.0808, 354.3149, 353.1136, 354.3901, 
    354.1587, 354.542, 354.885, 355.3168, 356.1126, 355.9285, 356.5941, 
    349.771, 350.1798, 350.1442, 350.5723, 350.8888, 351.5867, 352.6864, 
    352.2731, 353.0322, 353.1844, 352.0313, 352.739, 350.4537, 350.8208, 
    350.6026, 349.803, 352.3678, 351.046, 353.4765, 352.7674, 354.8361, 
    353.8072, 355.827, 356.6886, 357.5009, 358.4475, 350.4034, 350.1255, 
    350.6234, 351.3111, 351.9619, 352.8106, 352.8976, 353.0564, 353.4682, 
    353.8142, 353.1063, 353.9009, 350.9052, 352.4816, 350.0201, 350.7576, 
    351.2708, 351.0461, 352.2259, 352.501, 353.6182, 353.041, 356.4756, 
    354.9569, 359.1691, 357.993, 350.0284, 350.4026, 351.7157, 351.0849, 
    352.8674, 353.3029, 353.6571, 354.1092, 354.1583, 354.4261, 353.9871, 
    354.4089, 352.8124, 353.5261, 351.5674, 352.0441, 351.825, 351.5843, 
    352.327, 353.1173, 353.1348, 353.3881, 354.1003, 352.8746, 356.6704, 
    354.3262, 350.8106, 351.5419, 351.6455, 351.3549, 353.2592, 352.5736, 
    354.4196, 353.9211, 354.7381, 354.3321, 354.2723, 353.7509, 353.4259, 
    352.6049, 351.9368, 351.3954, 351.5303, 352.1122, 353.1658, 354.1624, 
    353.9441, 354.676, 352.7391, 353.5512, 353.2372, 354.056, 352.2619, 
    353.7879, 351.8714, 352.0397, 352.56, 353.6059, 353.8381, 354.0849, 
    353.9327, 353.1927, 353.0717, 352.5475, 352.4024, 352.0031, 351.6721, 
    351.9744, 352.2916, 353.1932, 354.005, 354.8898, 355.1065, 356.138, 
    355.2975, 356.6833, 355.5039, 357.5456, 353.8773, 355.4705, 352.5839, 
    352.8953, 353.4576, 354.7481, 354.0522, 354.8663, 353.067, 352.1319, 
    351.8907, 351.4275, 351.901, 351.8635, 352.3052, 352.1633, 353.2232, 
    352.654, 354.2706, 354.86, 356.5241, 357.543, 358.5804, 359.0378, 
    359.1771, 359.2352 ;

 FSH_R =
  347.9881, 348.9405, 348.757, 349.5184, 349.0963, 349.5947, 348.1876, 
    348.9778, 348.4735, 348.0735, 350.9944, 349.5525, 352.5055, 351.5862, 
    353.8953, 352.3621, 354.2044, 353.8517, 354.9145, 354.6101, 355.9674, 
    355.055, 356.6715, 355.7499, 355.8939, 355.0247, 349.8433, 350.8148, 
    349.7856, 349.9242, 349.8622, 349.1048, 348.7227, 347.9163, 348.0615, 
    348.6559, 349.9865, 349.5354, 350.6734, 350.6477, 351.9253, 351.3429, 
    353.4814, 352.8774, 354.6229, 354.184, 354.6021, 354.4754, 354.6038, 
    353.9601, 354.2359, 353.6696, 351.4496, 352.1104, 350.162, 348.9957, 
    348.2221, 347.665, 347.7427, 347.8907, 348.6594, 349.3752, 349.9204, 
    350.2849, 350.644, 351.7409, 352.3164, 353.6032, 353.3716, 353.7644, 
    354.1403, 354.7705, 354.6669, 354.9444, 353.7544, 354.5452, 353.2395, 
    353.5967, 350.7396, 349.6572, 349.1952, 348.7922, 347.8024, 348.4882, 
    348.2208, 348.8574, 349.2614, 349.0617, 350.2949, 349.8154, 352.3505, 
    351.2523, 354.0965, 353.4192, 354.2589, 353.8306, 354.5642, 353.904, 
    355.0478, 355.2965, 355.1265, 355.7802, 353.8673, 354.6019, 349.056, 
    349.0885, 349.2405, 348.5724, 348.5317, 347.9122, 348.4644, 348.6961, 
    349.285, 349.6328, 349.9636, 350.6906, 351.5018, 352.6481, 353.4631, 
    354.009, 353.6744, 353.9698, 353.6395, 353.4848, 355.2032, 354.2383, 
    355.6862, 355.6062, 354.9509, 355.6152, 349.1115, 348.924, 348.2723, 
    348.7823, 347.8456, 348.3731, 348.6718, 349.825, 350.0788, 350.3134, 
    350.7773, 351.3721, 352.4268, 353.3341, 354.1623, 354.1017, 354.123, 
    354.3077, 353.8498, 354.3829, 354.4722, 354.2385, 355.5955, 355.2079, 
    355.6045, 355.3522, 348.985, 349.3005, 349.13, 349.4505, 349.2245, 
    350.2285, 350.5295, 351.9493, 351.3603, 352.2912, 351.4538, 351.6118, 
    352.3203, 351.5103, 353.2837, 352.0808, 354.3149, 353.1136, 354.3901, 
    354.1587, 354.542, 354.885, 355.3168, 356.1126, 355.9285, 356.5941, 
    349.771, 350.1798, 350.1442, 350.5723, 350.8888, 351.5867, 352.6864, 
    352.2731, 353.0322, 353.1844, 352.0313, 352.739, 350.4537, 350.8208, 
    350.6026, 349.803, 352.3678, 351.046, 353.4765, 352.7674, 354.8361, 
    353.8072, 355.827, 356.6886, 357.5009, 358.4475, 350.4034, 350.1255, 
    350.6234, 351.3111, 351.9619, 352.8106, 352.8976, 353.0564, 353.4682, 
    353.8142, 353.1063, 353.9009, 350.9052, 352.4816, 350.0201, 350.7576, 
    351.2708, 351.0461, 352.2259, 352.501, 353.6182, 353.041, 356.4756, 
    354.9569, 359.1691, 357.993, 350.0284, 350.4026, 351.7157, 351.0849, 
    352.8674, 353.3029, 353.6571, 354.1092, 354.1583, 354.4261, 353.9871, 
    354.4089, 352.8124, 353.5261, 351.5674, 352.0441, 351.825, 351.5843, 
    352.327, 353.1173, 353.1348, 353.3881, 354.1003, 352.8746, 356.6704, 
    354.3262, 350.8106, 351.5419, 351.6455, 351.3549, 353.2592, 352.5736, 
    354.4196, 353.9211, 354.7381, 354.3321, 354.2723, 353.7509, 353.4259, 
    352.6049, 351.9368, 351.3954, 351.5303, 352.1122, 353.1658, 354.1624, 
    353.9441, 354.676, 352.7391, 353.5512, 353.2372, 354.056, 352.2619, 
    353.7879, 351.8714, 352.0397, 352.56, 353.6059, 353.8381, 354.0849, 
    353.9327, 353.1927, 353.0717, 352.5475, 352.4024, 352.0031, 351.6721, 
    351.9744, 352.2916, 353.1932, 354.005, 354.8898, 355.1065, 356.138, 
    355.2975, 356.6833, 355.5039, 357.5456, 353.8773, 355.4705, 352.5839, 
    352.8953, 353.4576, 354.7481, 354.0522, 354.8663, 353.067, 352.1319, 
    351.8907, 351.4275, 351.901, 351.8635, 352.3052, 352.1633, 353.2232, 
    352.654, 354.2706, 354.86, 356.5241, 357.543, 358.5804, 359.0378, 
    359.1771, 359.2352 ;

 FSH_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSH_V =
  -6.729109, -6.729638, -6.72954, -6.729949, -6.729727, -6.729991, -6.729233, 
    -6.729654, -6.729388, -6.729162, -6.730729, -6.729969, -6.731568, 
    -6.731074, -6.73233, -6.731484, -6.732502, -6.732317, -6.732904, 
    -6.732737, -6.733465, -6.732982, -6.733862, -6.733356, -6.73343, 
    -6.732964, -6.730132, -6.73063, -6.7301, -6.730172, -6.730142, -6.729727, 
    -6.729511, -6.729077, -6.729156, -6.729482, -6.730204, -6.729966, 
    -6.730588, -6.730575, -6.731261, -6.73095, -6.732113, -6.731785, 
    -6.732744, -6.732501, -6.73273, -6.732662, -6.732731, -6.732376, 
    -6.732527, -6.732218, -6.731006, -6.731359, -6.730303, -6.729653, 
    -6.729249, -6.72894, -6.728981, -6.729059, -6.729484, -6.729879, 
    -6.730177, -6.730375, -6.730572, -6.73114, -6.731464, -6.732174, 
    -6.732056, -6.732264, -6.732477, -6.732822, -6.732767, -6.732916, 
    -6.732265, -6.732695, -6.731986, -6.732178, -6.730587, -6.730032, 
    -6.729764, -6.729558, -6.729013, -6.729392, -6.729247, -6.729599, 
    -6.729817, -6.729711, -6.730381, -6.730119, -6.731484, -6.730896, 
    -6.732452, -6.732081, -6.732543, -6.732309, -6.732707, -6.732349, 
    -6.732975, -6.733107, -6.733016, -6.733379, -6.732328, -6.732727, 
    -6.729706, -6.729723, -6.729807, -6.729436, -6.729416, -6.729074, 
    -6.729383, -6.729506, -6.729833, -6.730019, -6.730198, -6.730594, 
    -6.73103, -6.731651, -6.732104, -6.732407, -6.732224, -6.732385, 
    -6.732203, -6.73212, -6.733055, -6.732526, -6.733327, -6.733284, 
    -6.732918, -6.733289, -6.729735, -6.729636, -6.729278, -6.729558, 
    -6.729038, -6.729331, -6.729488, -6.730116, -6.730263, -6.730388, 
    -6.730643, -6.730966, -6.731532, -6.73203, -6.732491, -6.732458, 
    -6.73247, -6.732568, -6.732318, -6.73261, -6.732656, -6.732531, 
    -6.733278, -6.733065, -6.733283, -6.733145, -6.729669, -6.729839, 
    -6.729746, -6.729918, -6.729794, -6.730333, -6.730495, -6.731264, 
    -6.730958, -6.731456, -6.731011, -6.731088, -6.731456, -6.731039, 
    -6.731995, -6.731332, -6.732572, -6.731894, -6.732614, -6.732489, 
    -6.7327, -6.732884, -6.733124, -6.733556, -6.733458, -6.733825, 
    -6.730095, -6.730311, -6.730299, -6.730531, -6.730701, -6.731079, 
    -6.731677, -6.731454, -6.731871, -6.731952, -6.731324, -6.731702, 
    -6.730462, -6.730655, -6.730545, -6.730108, -6.731496, -6.730778, 
    -6.732111, -6.731723, -6.732857, -6.732285, -6.733401, -6.733861, 
    -6.734328, -6.734835, -6.730437, -6.730289, -6.730561, -6.730924, 
    -6.731281, -6.731745, -6.731797, -6.731882, -6.732111, -6.732299, 
    -6.731902, -6.732347, -6.730685, -6.731561, -6.730227, -6.730618, 
    -6.730906, -6.730787, -6.731431, -6.73158, -6.732184, -6.731876, 
    -6.733741, -6.732913, -6.735246, -6.734588, -6.730236, -6.730441, 
    -6.731143, -6.730809, -6.73178, -6.732016, -6.732214, -6.732456, 
    -6.732488, -6.732632, -6.732395, -6.732625, -6.731746, -6.73214, 
    -6.731071, -6.731327, -6.731211, -6.73108, -6.731485, -6.731906, 
    -6.731926, -6.732059, -6.732414, -6.731784, -6.733827, -6.732543, 
    -6.730663, -6.731041, -6.73111, -6.73096, -6.731992, -6.731616, -6.73263, 
    -6.732358, -6.732807, -6.732583, -6.732549, -6.732265, -6.732084, 
    -6.731631, -6.731266, -6.730983, -6.73105, -6.731362, -6.731935, 
    -6.732485, -6.732363, -6.732773, -6.731709, -6.732149, -6.731975, 
    -6.73243, -6.731446, -6.732249, -6.731237, -6.731328, -6.731609, 
    -6.732171, -6.732313, -6.732443, -6.732365, -6.731951, -6.731888, 
    -6.731605, -6.731521, -6.731309, -6.731128, -6.73129, -6.731459, 
    -6.731956, -6.732399, -6.732885, -6.733009, -6.733551, -6.733094, 
    -6.733832, -6.733181, -6.734321, -6.732313, -6.733184, -6.731626, 
    -6.731796, -6.732092, -6.732797, -6.732429, -6.732865, -6.731887, 
    -6.731367, -6.731246, -6.730998, -6.731252, -6.731232, -6.731474, 
    -6.731397, -6.731973, -6.731664, -6.732545, -6.732864, -6.733782, 
    -6.734339, -6.734925, -6.735178, -6.735256, -6.735288 ;

 FSM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSNO_EFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSR =
  1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179 ;

 FSRND =
  0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234 ;

 FSRNDLN =
  0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495 ;

 FSRNI =
  0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666 ;

 FSRVD =
  0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223 ;

 FSRVDLN =
  0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609 ;

 FSRVI =
  0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671 ;

 FUELC =
  0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806 ;

 F_DENIT =
  2.431536e-36, 2.080171e-35, 1.377042e-35, 7.51097e-35, 2.945023e-35, 
    8.881373e-35, 3.775778e-36, 2.262524e-35, 7.249973e-36, 2.95697e-36, 
    1.808846e-33, 8.093939e-35, 3.946951e-32, 6.045991e-33, 6.088165e-31, 
    2.958383e-32, 1.100823e-30, 5.589807e-31, 4.199307e-30, 2.372932e-30, 
    2.909635e-29, 5.454859e-30, 1.022441e-28, 1.959256e-29, 2.545516e-29, 
    5.157598e-30, 1.529097e-34, 1.237951e-33, 1.348288e-34, 1.824726e-34, 
    1.593225e-34, 3.003121e-35, 1.276494e-35, 2.058065e-36, 2.875827e-36, 
    1.096847e-35, 2.089805e-34, 7.787286e-35, 9.12848e-34, 8.643058e-34, 
    1.214609e-32, 3.736812e-33, 2.72498e-31, 8.287591e-32, 2.430399e-30, 
    1.057477e-30, 2.337914e-30, 1.840018e-30, 2.345202e-30, 6.887896e-31, 
    1.167867e-30, 3.928743e-31, 4.667509e-33, 1.773161e-32, 3.054395e-34, 
    2.358835e-35, 4.088082e-36, 1.149436e-36, 1.377033e-36, 1.940986e-36, 
    1.105402e-35, 5.469746e-35, 1.807634e-34, 3.977145e-34, 8.575428e-34, 
    8.34156e-33, 2.69561e-32, 3.457341e-31, 2.197837e-31, 4.725023e-31, 
    9.728318e-31, 3.209095e-30, 2.641e-30, 4.442478e-30, 4.630589e-31, 
    2.100941e-30, 1.695494e-31, 3.410151e-31, 1.055934e-33, 1.017697e-34, 
    3.678611e-35, 1.490986e-35, 1.581801e-36, 7.500951e-36, 4.076749e-36, 
    1.724691e-35, 4.25128e-35, 2.724771e-35, 4.063328e-34, 1.438516e-34, 
    2.887758e-32, 3.095547e-33, 8.94634e-31, 2.41262e-31, 1.219711e-30, 
    5.363627e-31, 2.177187e-30, 6.179375e-31, 5.384613e-30, 8.539326e-30, 
    6.233685e-30, 2.06851e-29, 5.758325e-31, 2.338045e-30, 2.691009e-35, 
    2.894075e-35, 4.057476e-35, 9.080108e-36, 8.27686e-36, 2.039305e-36, 
    7.101458e-36, 1.200639e-35, 4.477733e-35, 9.648016e-35, 1.986333e-34, 
    9.472638e-34, 5.205024e-33, 5.251311e-32, 2.62879e-31, 7.563291e-31, 
    3.964653e-31, 7.014704e-31, 3.705541e-31, 2.741184e-31, 7.187649e-30, 
    1.173657e-30, 1.743426e-29, 1.506449e-29, 4.497641e-30, 1.531475e-29, 
    3.04559e-35, 2.002432e-35, 4.583814e-36, 1.456866e-35, 1.747991e-36, 
    5.770927e-36, 1.137196e-35, 1.470528e-34, 2.549317e-34, 4.230895e-34, 
    1.138245e-33, 3.971221e-33, 3.365823e-32, 2.043549e-31, 1.014278e-30, 
    9.032062e-31, 9.408806e-31, 1.338794e-30, 5.567699e-31, 1.544329e-30, 
    1.829777e-30, 1.173308e-30, 1.477218e-29, 7.244453e-30, 1.501769e-29, 
    9.453937e-30, 2.295419e-35, 4.635668e-35, 3.173496e-35, 6.461318e-35, 
    3.918533e-35, 3.528461e-34, 6.730773e-34, 1.277267e-32, 3.875749e-33, 
    2.559798e-32, 4.706361e-33, 6.374028e-33, 2.720699e-32, 5.162966e-33, 
    1.852806e-31, 1.671785e-32, 1.357209e-30, 1.32692e-31, 1.565558e-30, 
    1.007367e-30, 2.086567e-30, 3.976023e-30, 8.858512e-30, 3.775103e-29, 
    2.707442e-29, 8.909693e-29, 1.30531e-34, 3.17464e-34, 2.936628e-34, 
    7.362291e-34, 1.441659e-33, 6.048335e-33, 5.665552e-32, 2.464709e-32, 
    1.126559e-31, 1.521901e-31, 1.507442e-32, 6.296677e-32, 5.718368e-34, 
    1.250379e-33, 7.855341e-34, 1.400796e-34, 2.989184e-32, 2.010164e-33, 
    2.698833e-31, 6.659578e-32, 3.628413e-30, 5.134083e-31, 2.252845e-29, 
    1.054976e-28, 4.337753e-28, 2.162218e-27, 5.131526e-34, 2.820386e-34, 
    8.205746e-34, 3.501788e-33, 1.309011e-32, 7.259584e-32, 8.627697e-32, 
    1.182309e-31, 2.654278e-31, 5.197211e-31, 1.305896e-31, 6.143558e-31, 
    1.497649e-33, 3.758781e-32, 2.246509e-34, 1.09386e-33, 3.217284e-33, 
    2.008247e-33, 2.239435e-32, 3.903964e-32, 3.558205e-31, 1.146259e-31, 
    7.23638e-29, 4.552815e-30, 7.106188e-27, 1.00624e-27, 2.285472e-34, 
    5.120692e-34, 7.901357e-33, 2.178861e-33, 8.125475e-32, 1.921216e-31, 
    3.833498e-31, 9.169636e-31, 1.006659e-30, 1.676492e-30, 7.251408e-31, 
    1.62218e-30, 7.285792e-32, 2.972194e-31, 5.810477e-33, 1.548275e-32, 
    9.881065e-33, 6.016816e-33, 2.748668e-32, 1.334958e-31, 1.379941e-31, 
    2.271224e-31, 9.0572e-31, 8.242193e-32, 1.024441e-28, 1.392712e-30, 
    1.22124e-33, 5.522901e-33, 6.830898e-33, 3.829655e-33, 1.76336e-31, 
    4.519103e-32, 1.655817e-30, 6.386244e-31, 3.018376e-30, 1.402101e-30, 
    1.25149e-30, 4.59802e-31, 2.444659e-31, 4.81349e-32, 1.243548e-32, 
    4.166146e-33, 5.380952e-33, 1.778853e-32, 1.468531e-31, 1.015282e-30, 
    6.682074e-31, 2.686088e-30, 6.2921e-32, 3.123257e-31, 1.689693e-31, 
    8.278788e-31, 2.41056e-32, 4.962282e-31, 1.086891e-32, 1.533495e-32, 
    4.397302e-32, 3.477105e-31, 5.442648e-31, 8.753326e-31, 6.531403e-31, 
    1.547918e-31, 1.218636e-31, 4.286784e-32, 3.203159e-32, 1.422964e-32, 
    7.213664e-33, 1.34234e-32, 2.560963e-32, 1.548728e-31, 7.510358e-31, 
    4.012579e-30, 6.003471e-30, 3.959985e-29, 8.568919e-30, 1.048367e-28, 
    1.256413e-29, 4.701216e-28, 5.885199e-31, 1.178497e-29, 4.611026e-32, 
    8.586307e-32, 2.603937e-31, 3.081409e-30, 8.217949e-31, 3.843672e-30, 
    1.207228e-31, 1.853259e-32, 1.130717e-32, 4.455016e-33, 1.154876e-32, 
    1.069319e-32, 2.629645e-32, 1.971957e-32, 1.642661e-31, 5.306551e-32, 
    1.247989e-30, 3.797551e-30, 7.874024e-29, 4.669595e-28, 2.693259e-27, 
    5.730218e-27, 7.194341e-27, 7.90995e-27 ;

 F_DENIT_vr =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1.967257e-35, 1.682981e-34, 1.114108e-34, 6.076818e-34, 2.382698e-34, 
    7.185555e-34, 3.054827e-35, 1.830516e-34, 5.865657e-35, 2.392363e-35, 
    1.463464e-32, 6.548475e-34, 3.193316e-31, 4.891564e-32, 4.925685e-30, 
    2.393507e-31, 8.906308e-30, 4.522484e-30, 3.397488e-29, 1.919842e-29, 
    2.354066e-28, 4.413303e-29, 8.272155e-28, 1.585154e-28, 2.059473e-28, 
    4.172802e-29, 1.23713e-33, 1.001576e-32, 1.090845e-33, 1.476311e-33, 
    1.289013e-33, 2.429702e-34, 1.032759e-34, 1.665096e-35, 2.326714e-35, 
    8.874144e-35, 1.690776e-33, 6.300374e-34, 7.38548e-33, 6.992745e-33, 
    9.826902e-32, 3.023302e-32, 2.20467e-30, 6.705151e-31, 1.966336e-29, 
    8.555611e-30, 1.891511e-29, 1.488683e-29, 1.897407e-29, 5.572714e-30, 
    9.448731e-30, 3.178585e-30, 3.776291e-32, 1.434592e-31, 2.471186e-33, 
    1.908437e-34, 3.3075e-35, 9.29962e-36, 1.114101e-35, 1.570372e-35, 
    8.943358e-35, 4.425348e-34, 1.462483e-33, 3.217745e-33, 6.938028e-33, 
    6.748815e-32, 2.180907e-31, 2.797193e-30, 1.77818e-30, 3.822822e-30, 
    7.870784e-30, 2.596347e-29, 2.136725e-29, 3.594227e-29, 3.74642e-30, 
    1.699785e-29, 1.371755e-30, 2.759014e-30, 8.543131e-33, 8.233769e-34, 
    2.976213e-34, 1.206296e-34, 1.279771e-35, 6.068712e-35, 3.298331e-35, 
    1.395377e-34, 3.439536e-34, 2.204501e-34, 3.287472e-33, 1.163844e-33, 
    2.336367e-31, 2.504481e-32, 7.238118e-30, 1.951952e-30, 9.868184e-30, 
    4.339491e-30, 1.761473e-29, 4.99948e-30, 4.35647e-29, 6.908819e-29, 
    5.043419e-29, 1.673547e-28, 4.658825e-30, 1.891616e-29, 2.177186e-34, 
    2.341478e-34, 3.282737e-34, 7.346344e-35, 6.696469e-35, 1.649919e-35, 
    5.7455e-35, 9.71388e-35, 3.622751e-34, 7.805815e-34, 1.607061e-33, 
    7.663924e-33, 4.211172e-32, 4.248621e-31, 2.126847e-30, 6.11915e-30, 
    3.207639e-30, 5.67531e-30, 2.998001e-30, 2.21778e-30, 5.815232e-29, 
    9.495581e-30, 1.410535e-28, 1.218806e-28, 3.638857e-29, 1.239053e-28, 
    2.464062e-34, 1.620086e-34, 3.708576e-35, 1.17869e-34, 1.414228e-35, 
    4.669021e-35, 9.200585e-35, 1.189744e-33, 2.062548e-33, 3.423044e-33, 
    9.209077e-33, 3.212953e-32, 2.72315e-31, 1.653352e-30, 8.206112e-30, 
    7.307472e-30, 7.61228e-30, 1.083164e-29, 4.504598e-30, 1.249454e-29, 
    1.480398e-29, 9.49276e-30, 1.195157e-28, 5.861191e-29, 1.21502e-28, 
    7.648794e-29, 1.85713e-34, 3.75053e-34, 2.567546e-34, 5.227588e-34, 
    3.170325e-34, 2.854734e-33, 5.445593e-33, 1.033385e-31, 3.13571e-32, 
    2.071028e-31, 3.807724e-32, 5.156965e-32, 2.201207e-31, 4.177144e-32, 
    1.49903e-30, 1.352572e-31, 1.098063e-29, 1.073556e-30, 1.266629e-29, 
    8.150196e-30, 1.688156e-29, 3.216838e-29, 7.16706e-29, 3.054282e-28, 
    2.19048e-28, 7.208468e-28, 1.056073e-33, 2.568472e-33, 2.375906e-33, 
    5.956528e-33, 1.166387e-32, 4.89346e-32, 4.583766e-31, 1.994095e-31, 
    9.11453e-31, 1.231308e-30, 1.219609e-31, 5.094384e-31, 4.626498e-33, 
    1.011631e-32, 6.355435e-33, 1.133327e-33, 2.418426e-31, 1.626341e-32, 
    2.183515e-30, 5.387992e-31, 2.9356e-29, 4.153776e-30, 1.822685e-28, 
    8.53538e-28, 3.509498e-27, 1.749362e-26, 4.151708e-33, 2.281859e-33, 
    6.638933e-33, 2.833154e-32, 1.059067e-31, 5.873432e-31, 6.980316e-31, 
    9.565577e-31, 2.147467e-30, 4.204851e-30, 1.056547e-30, 4.970501e-30, 
    1.211687e-32, 3.041076e-31, 1.817559e-33, 8.849973e-33, 2.602973e-32, 
    1.62479e-32, 1.811835e-31, 3.158537e-31, 2.878798e-30, 9.273917e-31, 
    5.854659e-28, 3.683497e-29, 5.749327e-26, 8.141073e-27, 1.849082e-33, 
    4.142942e-33, 6.392664e-32, 1.762827e-32, 6.57399e-31, 1.554377e-30, 
    3.101526e-30, 7.418777e-30, 8.144464e-30, 1.356381e-29, 5.866818e-30, 
    1.31244e-29, 5.894636e-31, 2.404681e-30, 4.701019e-32, 1.252646e-31, 
    7.994366e-32, 4.86796e-32, 2.223835e-31, 1.08006e-30, 1.116454e-30, 
    1.837555e-30, 7.32781e-30, 6.668421e-31, 8.288337e-28, 1.126786e-29, 
    9.880553e-33, 4.468353e-32, 5.5266e-32, 3.098417e-32, 1.426662e-30, 
    3.656221e-31, 1.339654e-29, 5.166848e-30, 2.442044e-29, 1.134383e-29, 
    1.01253e-29, 3.72007e-30, 1.977874e-30, 3.894398e-31, 1.006103e-31, 
    3.370658e-32, 4.353509e-32, 1.439197e-31, 1.188129e-30, 8.214235e-30, 
    5.406193e-30, 2.173204e-29, 5.09068e-31, 2.5269e-30, 1.367062e-30, 
    6.698029e-30, 1.950286e-31, 4.01478e-30, 8.793588e-32, 1.240688e-31, 
    3.557678e-31, 2.813183e-30, 4.403424e-30, 7.081958e-30, 5.284292e-30, 
    1.252357e-30, 9.859483e-31, 3.468262e-31, 2.591545e-31, 1.151262e-31, 
    5.83628e-32, 1.086033e-31, 2.071971e-31, 1.253013e-30, 6.076324e-30, 
    3.246413e-29, 4.857163e-29, 3.203862e-28, 6.932762e-29, 8.481906e-28, 
    1.016512e-28, 3.803561e-27, 4.761474e-30, 9.534733e-29, 3.730593e-31, 
    6.94683e-31, 2.106739e-30, 2.493042e-29, 6.648807e-30, 3.109758e-29, 
    9.767187e-31, 1.499396e-31, 9.148169e-32, 3.604371e-32, 9.343632e-32, 
    8.65142e-32, 2.127538e-31, 1.59543e-31, 1.32901e-30, 4.293313e-31, 
    1.009697e-29, 3.072443e-29, 6.370551e-28, 3.777978e-27, 2.179006e-26, 
    4.636085e-26, 5.820647e-26, 6.399617e-26,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 F_N2O_DENIT =
  5.253709e-38, 4.494531e-37, 2.975312e-37, 1.622862e-36, 6.363179e-37, 
    1.918958e-36, 8.15815e-38, 4.888534e-37, 1.566469e-37, 6.388988e-38, 
    3.908295e-35, 1.748821e-36, 8.528004e-34, 1.306331e-34, 1.315443e-32, 
    6.392049e-34, 2.3785e-32, 1.207765e-32, 9.073259e-32, 5.12709e-32, 
    6.286719e-31, 1.178608e-31, 2.209143e-30, 4.233279e-31, 5.499984e-31, 
    1.11438e-31, 3.303852e-36, 2.674786e-35, 2.913186e-36, 3.942604e-36, 
    3.44241e-36, 6.488707e-37, 2.758064e-37, 4.446766e-38, 6.213666e-38, 
    2.369908e-37, 4.515348e-36, 1.682564e-36, 1.97235e-35, 1.867467e-35, 
    2.624352e-34, 8.073966e-35, 5.887745e-33, 1.790664e-33, 5.251256e-32, 
    2.284844e-32, 5.05143e-32, 3.975646e-32, 5.067176e-32, 1.488238e-32, 
    2.523358e-32, 8.488663e-33, 1.008488e-34, 3.831191e-34, 6.599496e-36, 
    5.096627e-37, 8.832932e-38, 2.483534e-38, 2.975291e-38, 4.1938e-38, 
    2.388393e-37, 1.181823e-36, 3.905675e-36, 8.593241e-36, 1.852855e-35, 
    1.802324e-34, 5.824286e-34, 7.470126e-33, 4.74877e-33, 1.020915e-32, 
    2.101955e-32, 6.933751e-32, 5.706293e-32, 9.598667e-32, 1.000511e-32, 
    4.53941e-32, 3.663381e-33, 7.368165e-33, 2.28151e-35, 2.198892e-36, 
    7.948208e-37, 3.221505e-37, 3.417725e-38, 1.620696e-37, 8.808444e-38, 
    3.726462e-37, 9.185549e-37, 5.887291e-37, 8.779453e-36, 3.108136e-36, 
    6.239453e-34, 6.688413e-35, 1.932997e-32, 5.212843e-33, 2.635376e-32, 
    1.158895e-32, 4.704154e-32, 1.335151e-32, 1.16343e-31, 1.845055e-31, 
    1.346885e-31, 4.469338e-31, 1.244176e-32, 5.051712e-32, 5.814343e-37, 
    6.253098e-37, 8.766805e-37, 1.961898e-37, 1.788343e-37, 4.406233e-38, 
    1.53438e-37, 2.594166e-37, 9.674838e-37, 2.084604e-36, 4.291782e-36, 
    2.046711e-35, 1.124627e-34, 1.134628e-33, 5.679912e-33, 1.634167e-32, 
    8.566253e-33, 1.515637e-32, 8.0064e-33, 5.922758e-33, 1.553004e-31, 
    2.53587e-32, 3.766944e-31, 3.254917e-31, 9.717855e-32, 3.308989e-31, 
    6.580469e-37, 4.326564e-37, 9.904037e-38, 3.147784e-37, 3.776805e-38, 
    1.246898e-37, 2.457087e-37, 3.177304e-36, 5.508195e-36, 9.141507e-36, 
    2.459356e-35, 8.580444e-35, 7.272386e-34, 4.415408e-33, 2.191507e-32, 
    1.951518e-32, 2.03292e-32, 2.892674e-32, 1.202989e-32, 3.336765e-32, 
    3.95352e-32, 2.535116e-32, 3.19176e-31, 1.565277e-31, 3.244807e-31, 
    2.042671e-31, 4.959609e-37, 1.001608e-36, 6.856829e-37, 1.396068e-36, 
    8.466599e-37, 7.62379e-36, 1.454288e-35, 2.759736e-34, 8.374161e-35, 
    5.530843e-34, 1.016883e-34, 1.377208e-34, 5.878496e-34, 1.115539e-34, 
    4.003278e-33, 3.612152e-34, 2.932463e-32, 2.867017e-33, 3.382632e-32, 
    2.176574e-32, 4.508353e-32, 8.59082e-32, 1.91402e-31, 8.156699e-31, 
    5.84985e-31, 1.925078e-30, 2.820324e-36, 6.859304e-36, 6.345043e-36, 
    1.590738e-35, 3.114929e-35, 1.306837e-34, 1.224131e-33, 5.325388e-34, 
    2.434108e-33, 3.288306e-33, 3.257063e-34, 1.360496e-33, 1.235543e-35, 
    2.701639e-35, 1.697269e-35, 3.026638e-36, 6.458599e-34, 4.343273e-35, 
    5.831251e-33, 1.438906e-33, 7.839752e-32, 1.109299e-32, 4.867623e-31, 
    2.279439e-30, 9.372386e-30, 4.671804e-29, 1.108746e-35, 6.093882e-36, 
    1.772979e-35, 7.566161e-35, 2.828322e-34, 1.568547e-33, 1.864149e-33, 
    2.554563e-33, 5.734982e-33, 1.122939e-32, 2.821592e-33, 1.327412e-32, 
    3.235905e-35, 8.121434e-34, 4.853933e-36, 2.363455e-35, 6.951444e-35, 
    4.339131e-35, 4.83865e-34, 8.435124e-34, 7.688059e-33, 2.476673e-33, 
    1.563532e-30, 9.837068e-32, 1.535401e-28, 2.174136e-29, 4.938117e-36, 
    1.106405e-35, 1.707212e-34, 4.707769e-35, 1.755636e-33, 4.151088e-33, 
    8.282872e-33, 1.981243e-32, 2.175043e-32, 3.622322e-32, 1.56678e-32, 
    3.504974e-32, 1.574209e-33, 6.421891e-33, 1.255444e-34, 3.345289e-34, 
    2.134959e-34, 1.300027e-34, 5.938927e-34, 2.884385e-33, 2.981579e-33, 
    4.907336e-33, 1.95695e-32, 1.780855e-33, 2.213465e-30, 3.009171e-32, 
    2.638679e-35, 1.193309e-34, 1.475922e-34, 8.274568e-35, 3.810015e-33, 
    9.764229e-34, 3.577651e-32, 1.379848e-32, 6.521672e-32, 3.029459e-32, 
    2.70404e-32, 9.934743e-33, 5.282069e-33, 1.04003e-33, 2.686879e-34, 
    9.001609e-35, 1.162639e-34, 3.843491e-34, 3.172992e-33, 2.193676e-32, 
    1.443767e-32, 5.803712e-32, 1.359507e-33, 6.748286e-33, 3.650846e-33, 
    1.788762e-32, 5.208393e-34, 1.072179e-32, 2.348397e-34, 3.313355e-34, 
    9.50106e-34, 7.512829e-33, 1.175969e-32, 1.891293e-32, 1.411212e-32, 
    3.344518e-33, 2.633053e-33, 9.262268e-34, 6.920925e-34, 3.074536e-34, 
    1.558625e-34, 2.900336e-34, 5.533361e-34, 3.34627e-33, 1.62273e-32, 
    8.669803e-32, 1.297144e-31, 8.556164e-31, 1.851449e-31, 2.265159e-30, 
    2.714675e-31, 1.01577e-29, 1.271589e-32, 2.546326e-31, 9.962843e-34, 
    1.855206e-33, 5.626213e-33, 6.657865e-32, 1.775616e-32, 8.304854e-32, 
    2.608405e-33, 4.004256e-34, 2.443091e-34, 9.625758e-35, 2.495291e-34, 
    2.31043e-34, 5.681759e-34, 4.260722e-34, 3.549227e-33, 1.146563e-33, 
    2.696476e-32, 8.205202e-32, 1.701305e-30, 1.008938e-29, 5.819199e-29, 
    1.238101e-28, 1.554447e-28, 1.709065e-28 ;

 F_N2O_NIT =
  3.450677e-14, 3.469339e-14, 3.465707e-14, 3.480784e-14, 3.472418e-14, 
    3.482294e-14, 3.454457e-14, 3.470077e-14, 3.460102e-14, 3.452355e-14, 
    3.510123e-14, 3.481456e-14, 3.540027e-14, 3.521658e-14, 3.567887e-14, 
    3.537164e-14, 3.574098e-14, 3.567002e-14, 3.588384e-14, 3.582252e-14, 
    3.609659e-14, 3.591215e-14, 3.623908e-14, 3.605252e-14, 3.608166e-14, 
    3.590606e-14, 3.487221e-14, 3.506549e-14, 3.486076e-14, 3.488829e-14, 
    3.487594e-14, 3.472588e-14, 3.465036e-14, 3.449252e-14, 3.452115e-14, 
    3.46371e-14, 3.490065e-14, 3.48111e-14, 3.503704e-14, 3.503193e-14, 
    3.528422e-14, 3.517036e-14, 3.559567e-14, 3.547456e-14, 3.582508e-14, 
    3.573677e-14, 3.582091e-14, 3.579539e-14, 3.582124e-14, 3.569178e-14, 
    3.574721e-14, 3.563339e-14, 3.51917e-14, 3.532125e-14, 3.493548e-14, 
    3.470442e-14, 3.455139e-14, 3.444298e-14, 3.445829e-14, 3.448749e-14, 
    3.463777e-14, 3.477936e-14, 3.488744e-14, 3.495981e-14, 3.503119e-14, 
    3.52476e-14, 3.536244e-14, 3.562016e-14, 3.557362e-14, 3.56525e-14, 
    3.572799e-14, 3.585484e-14, 3.583395e-14, 3.588988e-14, 3.565043e-14, 
    3.580947e-14, 3.554708e-14, 3.561875e-14, 3.505054e-14, 3.483527e-14, 
    3.474387e-14, 3.466402e-14, 3.447006e-14, 3.460395e-14, 3.455113e-14, 
    3.467684e-14, 3.475682e-14, 3.471725e-14, 3.496178e-14, 3.486662e-14, 
    3.536925e-14, 3.515235e-14, 3.571918e-14, 3.558316e-14, 3.575181e-14, 
    3.566571e-14, 3.581328e-14, 3.568045e-14, 3.591071e-14, 3.596093e-14, 
    3.59266e-14, 3.605856e-14, 3.567308e-14, 3.582087e-14, 3.471616e-14, 
    3.472261e-14, 3.475267e-14, 3.462058e-14, 3.461251e-14, 3.449171e-14, 
    3.45992e-14, 3.464501e-14, 3.476146e-14, 3.483041e-14, 3.489602e-14, 
    3.504047e-14, 3.520211e-14, 3.542873e-14, 3.559197e-14, 3.570157e-14, 
    3.563435e-14, 3.569369e-14, 3.562735e-14, 3.559627e-14, 3.594209e-14, 
    3.574771e-14, 3.603955e-14, 3.602338e-14, 3.589118e-14, 3.602519e-14, 
    3.472713e-14, 3.469001e-14, 3.456126e-14, 3.4662e-14, 3.447856e-14, 
    3.458117e-14, 3.464023e-14, 3.486858e-14, 3.491886e-14, 3.496549e-14, 
    3.505769e-14, 3.517616e-14, 3.538444e-14, 3.556612e-14, 3.573237e-14, 
    3.572017e-14, 3.572446e-14, 3.576163e-14, 3.566957e-14, 3.577675e-14, 
    3.579474e-14, 3.574769e-14, 3.60212e-14, 3.594297e-14, 3.602302e-14, 
    3.597207e-14, 3.470208e-14, 3.476455e-14, 3.473078e-14, 3.479429e-14, 
    3.474953e-14, 3.49487e-14, 3.500852e-14, 3.528907e-14, 3.517383e-14, 
    3.535734e-14, 3.519245e-14, 3.522164e-14, 3.536329e-14, 3.520135e-14, 
    3.555606e-14, 3.531536e-14, 3.576307e-14, 3.552203e-14, 3.57782e-14, 
    3.573163e-14, 3.580874e-14, 3.587787e-14, 3.596494e-14, 3.612582e-14, 
    3.608854e-14, 3.622328e-14, 3.485779e-14, 3.493899e-14, 3.493186e-14, 
    3.501693e-14, 3.50799e-14, 3.52166e-14, 3.543634e-14, 3.535364e-14, 
    3.550554e-14, 3.553606e-14, 3.530531e-14, 3.544689e-14, 3.499337e-14, 
    3.506644e-14, 3.502294e-14, 3.486414e-14, 3.537263e-14, 3.511124e-14, 
    3.559463e-14, 3.545251e-14, 3.5868e-14, 3.566107e-14, 3.606801e-14, 
    3.624258e-14, 3.640731e-14, 3.660014e-14, 3.498336e-14, 3.492814e-14, 
    3.502706e-14, 3.516409e-14, 3.529151e-14, 3.54612e-14, 3.547859e-14, 
    3.551042e-14, 3.559295e-14, 3.566241e-14, 3.552046e-14, 3.567983e-14, 
    3.508336e-14, 3.539537e-14, 3.490722e-14, 3.505386e-14, 3.515597e-14, 
    3.511118e-14, 3.534416e-14, 3.539916e-14, 3.562308e-14, 3.550726e-14, 
    3.619943e-14, 3.589244e-14, 3.674734e-14, 3.650749e-14, 3.490885e-14, 
    3.498317e-14, 3.524239e-14, 3.511894e-14, 3.547254e-14, 3.555982e-14, 
    3.563085e-14, 3.572173e-14, 3.573156e-14, 3.578546e-14, 3.569714e-14, 
    3.578197e-14, 3.546153e-14, 3.560456e-14, 3.52127e-14, 3.530788e-14, 
    3.526409e-14, 3.521606e-14, 3.536436e-14, 3.552265e-14, 3.552607e-14, 
    3.557688e-14, 3.572023e-14, 3.547393e-14, 3.623907e-14, 3.576561e-14, 
    3.50643e-14, 3.520777e-14, 3.522832e-14, 3.517269e-14, 3.555106e-14, 
    3.541374e-14, 3.578415e-14, 3.568387e-14, 3.584824e-14, 3.576651e-14, 
    3.575449e-14, 3.564967e-14, 3.558447e-14, 3.542e-14, 3.528645e-14, 
    3.518072e-14, 3.520529e-14, 3.532147e-14, 3.553235e-14, 3.573239e-14, 
    3.568852e-14, 3.58357e-14, 3.544679e-14, 3.560961e-14, 3.554663e-14, 
    3.571096e-14, 3.535142e-14, 3.565745e-14, 3.527338e-14, 3.530698e-14, 
    3.541101e-14, 3.562069e-14, 3.56672e-14, 3.571683e-14, 3.56862e-14, 
    3.553774e-14, 3.551345e-14, 3.540847e-14, 3.537949e-14, 3.529964e-14, 
    3.523357e-14, 3.529392e-14, 3.535734e-14, 3.553779e-14, 3.570075e-14, 
    3.587881e-14, 3.592247e-14, 3.613108e-14, 3.596118e-14, 3.62417e-14, 
    3.600308e-14, 3.641664e-14, 3.567526e-14, 3.599618e-14, 3.541576e-14, 
    3.547808e-14, 3.559092e-14, 3.585038e-14, 3.571022e-14, 3.587417e-14, 
    3.55125e-14, 3.532548e-14, 3.527719e-14, 3.518714e-14, 3.527925e-14, 
    3.527175e-14, 3.535998e-14, 3.533161e-14, 3.554378e-14, 3.542974e-14, 
    3.575414e-14, 3.587285e-14, 3.620911e-14, 3.641593e-14, 3.662707e-14, 
    3.672044e-14, 3.674888e-14, 3.676077e-14 ;

 F_NIT =
  5.751129e-11, 5.782231e-11, 5.77618e-11, 5.801307e-11, 5.787363e-11, 
    5.803824e-11, 5.757428e-11, 5.783463e-11, 5.766837e-11, 5.753924e-11, 
    5.850205e-11, 5.802427e-11, 5.900044e-11, 5.86943e-11, 5.946479e-11, 
    5.895273e-11, 5.956829e-11, 5.945003e-11, 5.98064e-11, 5.97042e-11, 
    6.016099e-11, 5.985359e-11, 6.039847e-11, 6.008753e-11, 6.013609e-11, 
    5.984342e-11, 5.812035e-11, 5.844249e-11, 5.810127e-11, 5.814715e-11, 
    5.812656e-11, 5.787647e-11, 5.77506e-11, 5.748753e-11, 5.753525e-11, 
    5.77285e-11, 5.816776e-11, 5.80185e-11, 5.839507e-11, 5.838655e-11, 
    5.880704e-11, 5.861727e-11, 5.932612e-11, 5.912426e-11, 5.970846e-11, 
    5.956128e-11, 5.970153e-11, 5.965898e-11, 5.970206e-11, 5.948629e-11, 
    5.957868e-11, 5.938899e-11, 5.865284e-11, 5.886876e-11, 5.822581e-11, 
    5.784069e-11, 5.758565e-11, 5.740496e-11, 5.743048e-11, 5.747915e-11, 
    5.772962e-11, 5.79656e-11, 5.814573e-11, 5.826634e-11, 5.838532e-11, 
    5.874599e-11, 5.89374e-11, 5.936694e-11, 5.928936e-11, 5.942084e-11, 
    5.954665e-11, 5.975806e-11, 5.972325e-11, 5.981646e-11, 5.941738e-11, 
    5.968245e-11, 5.924514e-11, 5.936459e-11, 5.841757e-11, 5.805878e-11, 
    5.790644e-11, 5.777337e-11, 5.745011e-11, 5.767324e-11, 5.758522e-11, 
    5.779474e-11, 5.792804e-11, 5.786209e-11, 5.826964e-11, 5.811103e-11, 
    5.894874e-11, 5.858724e-11, 5.953196e-11, 5.930527e-11, 5.958635e-11, 
    5.944285e-11, 5.968881e-11, 5.946742e-11, 5.985118e-11, 5.993488e-11, 
    5.987766e-11, 6.009759e-11, 5.945513e-11, 5.970146e-11, 5.786027e-11, 
    5.787102e-11, 5.792112e-11, 5.770098e-11, 5.768752e-11, 5.748619e-11, 
    5.766532e-11, 5.774168e-11, 5.793577e-11, 5.805068e-11, 5.816003e-11, 
    5.840078e-11, 5.867018e-11, 5.904788e-11, 5.931994e-11, 5.950262e-11, 
    5.939058e-11, 5.948948e-11, 5.937891e-11, 5.932712e-11, 5.990348e-11, 
    5.957952e-11, 6.006592e-11, 6.003897e-11, 5.981864e-11, 6.004199e-11, 
    5.787856e-11, 5.781669e-11, 5.76021e-11, 5.777e-11, 5.746427e-11, 
    5.763529e-11, 5.773371e-11, 5.81143e-11, 5.819811e-11, 5.827582e-11, 
    5.842948e-11, 5.862694e-11, 5.897407e-11, 5.927687e-11, 5.955395e-11, 
    5.953362e-11, 5.954078e-11, 5.960272e-11, 5.944929e-11, 5.962792e-11, 
    5.96579e-11, 5.957948e-11, 6.003534e-11, 5.990495e-11, 6.003838e-11, 
    5.995345e-11, 5.78368e-11, 5.794092e-11, 5.788463e-11, 5.799048e-11, 
    5.791588e-11, 5.824784e-11, 5.834754e-11, 5.881512e-11, 5.862304e-11, 
    5.89289e-11, 5.865408e-11, 5.870273e-11, 5.893881e-11, 5.866892e-11, 
    5.926011e-11, 5.885894e-11, 5.960512e-11, 5.920338e-11, 5.963033e-11, 
    5.955271e-11, 5.968125e-11, 5.979645e-11, 5.994157e-11, 6.02097e-11, 
    6.014756e-11, 6.037214e-11, 5.809632e-11, 5.823166e-11, 5.821976e-11, 
    5.836154e-11, 5.846651e-11, 5.869434e-11, 5.906056e-11, 5.892273e-11, 
    5.91759e-11, 5.922678e-11, 5.884219e-11, 5.907815e-11, 5.832228e-11, 
    5.844406e-11, 5.837156e-11, 5.81069e-11, 5.895439e-11, 5.851873e-11, 
    5.932438e-11, 5.908751e-11, 5.978e-11, 5.943512e-11, 6.011336e-11, 
    6.04043e-11, 6.067884e-11, 6.100024e-11, 5.83056e-11, 5.821357e-11, 
    5.837842e-11, 5.860681e-11, 5.881918e-11, 5.910199e-11, 5.913098e-11, 
    5.918403e-11, 5.932159e-11, 5.943736e-11, 5.920077e-11, 5.946638e-11, 
    5.847227e-11, 5.899228e-11, 5.81787e-11, 5.84231e-11, 5.859329e-11, 
    5.851863e-11, 5.890693e-11, 5.89986e-11, 5.937181e-11, 5.917876e-11, 
    6.033238e-11, 5.982073e-11, 6.124556e-11, 6.084582e-11, 5.818141e-11, 
    5.830528e-11, 5.873731e-11, 5.853158e-11, 5.91209e-11, 5.926637e-11, 
    5.938476e-11, 5.953622e-11, 5.955259e-11, 5.964243e-11, 5.949524e-11, 
    5.963662e-11, 5.910255e-11, 5.934093e-11, 5.868784e-11, 5.884647e-11, 
    5.877347e-11, 5.869343e-11, 5.894061e-11, 5.920443e-11, 5.921012e-11, 
    5.929481e-11, 5.953371e-11, 5.912321e-11, 6.039846e-11, 5.960935e-11, 
    5.84405e-11, 5.867962e-11, 5.871387e-11, 5.862115e-11, 5.925176e-11, 
    5.90229e-11, 5.964024e-11, 5.947311e-11, 5.974706e-11, 5.961086e-11, 
    5.959081e-11, 5.941612e-11, 5.930744e-11, 5.903334e-11, 5.881075e-11, 
    5.863454e-11, 5.867549e-11, 5.886912e-11, 5.922059e-11, 5.955399e-11, 
    5.948087e-11, 5.972616e-11, 5.907799e-11, 5.934936e-11, 5.924438e-11, 
    5.951827e-11, 5.891904e-11, 5.942908e-11, 5.878897e-11, 5.884496e-11, 
    5.901835e-11, 5.936782e-11, 5.944533e-11, 5.952806e-11, 5.9477e-11, 
    5.922957e-11, 5.918908e-11, 5.901411e-11, 5.896582e-11, 5.883273e-11, 
    5.872262e-11, 5.88232e-11, 5.89289e-11, 5.922964e-11, 5.950125e-11, 
    5.979802e-11, 5.987078e-11, 6.021847e-11, 5.99353e-11, 6.040284e-11, 
    6.000513e-11, 6.069439e-11, 5.945876e-11, 5.999364e-11, 5.902626e-11, 
    5.913014e-11, 5.93182e-11, 5.975063e-11, 5.951704e-11, 5.979029e-11, 
    5.91875e-11, 5.887579e-11, 5.879532e-11, 5.864523e-11, 5.879874e-11, 
    5.878625e-11, 5.89333e-11, 5.888603e-11, 5.923963e-11, 5.904957e-11, 
    5.959024e-11, 5.978808e-11, 6.034851e-11, 6.069321e-11, 6.104511e-11, 
    6.120073e-11, 6.124814e-11, 6.126796e-11 ;

 F_NIT_vr =
  2.589009e-10, 2.599879e-10, 2.597761e-10, 2.606531e-10, 2.601664e-10, 
    2.607402e-10, 2.5912e-10, 2.600291e-10, 2.594484e-10, 2.589967e-10, 
    2.623539e-10, 2.606901e-10, 2.640862e-10, 2.630227e-10, 2.656951e-10, 
    2.639197e-10, 2.660532e-10, 2.656436e-10, 2.668764e-10, 2.665227e-10, 
    2.680994e-10, 2.670387e-10, 2.689177e-10, 2.678457e-10, 2.680129e-10, 
    2.670023e-10, 2.610272e-10, 2.621486e-10, 2.609601e-10, 2.6112e-10, 
    2.61048e-10, 2.601751e-10, 2.597352e-10, 2.588157e-10, 2.589822e-10, 
    2.596575e-10, 2.611899e-10, 2.606693e-10, 2.619813e-10, 2.619517e-10, 
    2.634134e-10, 2.62754e-10, 2.652141e-10, 2.64514e-10, 2.665371e-10, 
    2.660275e-10, 2.665125e-10, 2.66365e-10, 2.665136e-10, 2.657671e-10, 
    2.660863e-10, 2.654297e-10, 2.628806e-10, 2.636305e-10, 2.613937e-10, 
    2.600496e-10, 2.591586e-10, 2.585268e-10, 2.586155e-10, 2.587858e-10, 
    2.596609e-10, 2.604846e-10, 2.611127e-10, 2.615326e-10, 2.619467e-10, 
    2.632007e-10, 2.638655e-10, 2.653548e-10, 2.650861e-10, 2.65541e-10, 
    2.659766e-10, 2.667074e-10, 2.665869e-10, 2.669087e-10, 2.655278e-10, 
    2.664451e-10, 2.649306e-10, 2.653445e-10, 2.620606e-10, 2.608109e-10, 
    2.602789e-10, 2.598142e-10, 2.58684e-10, 2.594641e-10, 2.591561e-10, 
    2.59888e-10, 2.603532e-10, 2.601226e-10, 2.615438e-10, 2.609906e-10, 
    2.639045e-10, 2.626485e-10, 2.659261e-10, 2.651406e-10, 2.661136e-10, 
    2.65617e-10, 2.664673e-10, 2.657015e-10, 2.670281e-10, 2.673172e-10, 
    2.671191e-10, 2.678786e-10, 2.656573e-10, 2.665096e-10, 2.601178e-10, 
    2.601553e-10, 2.603299e-10, 2.595606e-10, 2.595135e-10, 2.588093e-10, 
    2.594353e-10, 2.59702e-10, 2.603795e-10, 2.607799e-10, 2.611608e-10, 
    2.619996e-10, 2.629363e-10, 2.642478e-10, 2.651912e-10, 2.658235e-10, 
    2.654355e-10, 2.657775e-10, 2.653945e-10, 2.652147e-10, 2.67208e-10, 
    2.660881e-10, 2.677685e-10, 2.676755e-10, 2.669141e-10, 2.676852e-10, 
    2.601812e-10, 2.599648e-10, 2.592148e-10, 2.598012e-10, 2.587322e-10, 
    2.593301e-10, 2.596735e-10, 2.610014e-10, 2.612935e-10, 2.615642e-10, 
    2.62099e-10, 2.627856e-10, 2.639913e-10, 2.650412e-10, 2.660009e-10, 
    2.659301e-10, 2.659547e-10, 2.661686e-10, 2.656375e-10, 2.662553e-10, 
    2.663585e-10, 2.660874e-10, 2.676623e-10, 2.672121e-10, 2.676724e-10, 
    2.673789e-10, 2.600347e-10, 2.603977e-10, 2.602009e-10, 2.605703e-10, 
    2.603094e-10, 2.614668e-10, 2.618137e-10, 2.634397e-10, 2.627719e-10, 
    2.638347e-10, 2.628794e-10, 2.630485e-10, 2.638678e-10, 2.629304e-10, 
    2.649821e-10, 2.635897e-10, 2.661766e-10, 2.647843e-10, 2.662633e-10, 
    2.659944e-10, 2.664387e-10, 2.66837e-10, 2.673378e-10, 2.68263e-10, 
    2.680481e-10, 2.688225e-10, 2.609395e-10, 2.614107e-10, 2.613693e-10, 
    2.618628e-10, 2.622277e-10, 2.630204e-10, 2.642918e-10, 2.638131e-10, 
    2.646912e-10, 2.648676e-10, 2.635325e-10, 2.643515e-10, 2.617238e-10, 
    2.621471e-10, 2.618949e-10, 2.609723e-10, 2.639205e-10, 2.62406e-10, 
    2.652034e-10, 2.643818e-10, 2.667793e-10, 2.655861e-10, 2.6793e-10, 
    2.689326e-10, 2.698779e-10, 2.709816e-10, 2.616681e-10, 2.613471e-10, 
    2.619211e-10, 2.627155e-10, 2.634533e-10, 2.644351e-10, 2.645354e-10, 
    2.647189e-10, 2.651955e-10, 2.655965e-10, 2.647761e-10, 2.656962e-10, 
    2.622445e-10, 2.640521e-10, 2.61222e-10, 2.620731e-10, 2.626649e-10, 
    2.624054e-10, 2.637549e-10, 2.640727e-10, 2.653661e-10, 2.646973e-10, 
    2.68684e-10, 2.669186e-10, 2.718233e-10, 2.704508e-10, 2.612348e-10, 
    2.61666e-10, 2.631686e-10, 2.624534e-10, 2.645001e-10, 2.650044e-10, 
    2.654141e-10, 2.659384e-10, 2.659946e-10, 2.663054e-10, 2.657956e-10, 
    2.662849e-10, 2.644342e-10, 2.652608e-10, 2.62994e-10, 2.635447e-10, 
    2.632911e-10, 2.630125e-10, 2.638708e-10, 2.647858e-10, 2.648055e-10, 
    2.650985e-10, 2.659247e-10, 2.645032e-10, 2.689101e-10, 2.661856e-10, 
    2.621365e-10, 2.629675e-10, 2.630866e-10, 2.627643e-10, 2.64953e-10, 
    2.641594e-10, 2.662979e-10, 2.657192e-10, 2.666666e-10, 2.661956e-10, 
    2.661256e-10, 2.65521e-10, 2.651439e-10, 2.641934e-10, 2.6342e-10, 
    2.628078e-10, 2.629496e-10, 2.636223e-10, 2.648411e-10, 2.659961e-10, 
    2.657426e-10, 2.66591e-10, 2.643458e-10, 2.652865e-10, 2.649221e-10, 
    2.65871e-10, 2.637991e-10, 2.655668e-10, 2.633471e-10, 2.635412e-10, 
    2.641428e-10, 2.653542e-10, 2.656224e-10, 2.659088e-10, 2.657316e-10, 
    2.648743e-10, 2.647337e-10, 2.641264e-10, 2.639584e-10, 2.634964e-10, 
    2.631133e-10, 2.634627e-10, 2.638291e-10, 2.648726e-10, 2.65813e-10, 
    2.668391e-10, 2.670905e-10, 2.682894e-10, 2.673123e-10, 2.689238e-10, 
    2.675521e-10, 2.699272e-10, 2.656692e-10, 2.675185e-10, 2.641704e-10, 
    2.645304e-10, 2.651818e-10, 2.66678e-10, 2.658699e-10, 2.668148e-10, 
    2.64728e-10, 2.636457e-10, 2.633662e-10, 2.628446e-10, 2.633776e-10, 
    2.633343e-10, 2.638447e-10, 2.636801e-10, 2.649065e-10, 2.642475e-10, 
    2.6612e-10, 2.668042e-10, 2.687379e-10, 2.699241e-10, 2.711335e-10, 
    2.716671e-10, 2.718296e-10, 2.718972e-10,
  1.73745e-10, 1.746601e-10, 1.744822e-10, 1.752209e-10, 1.748111e-10, 
    1.752949e-10, 1.739305e-10, 1.746963e-10, 1.742074e-10, 1.738275e-10, 
    1.766566e-10, 1.752539e-10, 1.781183e-10, 1.772211e-10, 1.794777e-10, 
    1.779784e-10, 1.797805e-10, 1.794347e-10, 1.804767e-10, 1.80178e-10, 
    1.815118e-10, 1.806146e-10, 1.822047e-10, 1.812976e-10, 1.814393e-10, 
    1.805849e-10, 1.755363e-10, 1.764817e-10, 1.754802e-10, 1.75615e-10, 
    1.755546e-10, 1.748195e-10, 1.744491e-10, 1.736753e-10, 1.738158e-10, 
    1.743843e-10, 1.756756e-10, 1.752372e-10, 1.763433e-10, 1.763183e-10, 
    1.775518e-10, 1.769953e-10, 1.790722e-10, 1.784813e-10, 1.801905e-10, 
    1.797602e-10, 1.801702e-10, 1.800459e-10, 1.801718e-10, 1.795409e-10, 
    1.798111e-10, 1.792563e-10, 1.770994e-10, 1.777325e-10, 1.758461e-10, 
    1.74714e-10, 1.73964e-10, 1.734322e-10, 1.735073e-10, 1.736506e-10, 
    1.743876e-10, 1.750817e-10, 1.756111e-10, 1.759654e-10, 1.763147e-10, 
    1.773724e-10, 1.779337e-10, 1.791916e-10, 1.789647e-10, 1.793493e-10, 
    1.797174e-10, 1.803355e-10, 1.802338e-10, 1.805061e-10, 1.793394e-10, 
    1.801145e-10, 1.788354e-10, 1.79185e-10, 1.764085e-10, 1.753555e-10, 
    1.749074e-10, 1.745163e-10, 1.735651e-10, 1.742218e-10, 1.739628e-10, 
    1.745794e-10, 1.749713e-10, 1.747775e-10, 1.759751e-10, 1.755091e-10, 
    1.779669e-10, 1.769071e-10, 1.796745e-10, 1.790113e-10, 1.798336e-10, 
    1.794139e-10, 1.801331e-10, 1.794858e-10, 1.806076e-10, 1.80852e-10, 
    1.80685e-10, 1.813272e-10, 1.794499e-10, 1.801701e-10, 1.74772e-10, 
    1.748036e-10, 1.749509e-10, 1.743034e-10, 1.742638e-10, 1.736714e-10, 
    1.741986e-10, 1.744232e-10, 1.749941e-10, 1.753318e-10, 1.756531e-10, 
    1.763601e-10, 1.771504e-10, 1.782575e-10, 1.790542e-10, 1.795888e-10, 
    1.79261e-10, 1.795503e-10, 1.792269e-10, 1.790754e-10, 1.807603e-10, 
    1.798136e-10, 1.812348e-10, 1.811561e-10, 1.805126e-10, 1.81165e-10, 
    1.748258e-10, 1.746439e-10, 1.740125e-10, 1.745066e-10, 1.736069e-10, 
    1.741102e-10, 1.743997e-10, 1.755186e-10, 1.75765e-10, 1.759932e-10, 
    1.764444e-10, 1.770238e-10, 1.780413e-10, 1.789281e-10, 1.797389e-10, 
    1.796795e-10, 1.797004e-10, 1.798815e-10, 1.794328e-10, 1.799552e-10, 
    1.800428e-10, 1.798136e-10, 1.811456e-10, 1.807648e-10, 1.811545e-10, 
    1.809065e-10, 1.74703e-10, 1.750092e-10, 1.748437e-10, 1.751548e-10, 
    1.749355e-10, 1.759108e-10, 1.762036e-10, 1.775753e-10, 1.770123e-10, 
    1.77909e-10, 1.771034e-10, 1.77246e-10, 1.779377e-10, 1.77147e-10, 
    1.78879e-10, 1.777038e-10, 1.798885e-10, 1.787128e-10, 1.799623e-10, 
    1.797354e-10, 1.801112e-10, 1.804478e-10, 1.808718e-10, 1.816544e-10, 
    1.814731e-10, 1.821283e-10, 1.754659e-10, 1.758634e-10, 1.758286e-10, 
    1.762449e-10, 1.76553e-10, 1.772215e-10, 1.782948e-10, 1.77891e-10, 
    1.786327e-10, 1.787816e-10, 1.776551e-10, 1.783463e-10, 1.761297e-10, 
    1.764871e-10, 1.762744e-10, 1.754971e-10, 1.779837e-10, 1.767063e-10, 
    1.790674e-10, 1.783739e-10, 1.803998e-10, 1.793913e-10, 1.813733e-10, 
    1.822218e-10, 1.830223e-10, 1.839576e-10, 1.760807e-10, 1.758104e-10, 
    1.762945e-10, 1.769645e-10, 1.775875e-10, 1.784161e-10, 1.785011e-10, 
    1.786564e-10, 1.790592e-10, 1.793979e-10, 1.787053e-10, 1.794829e-10, 
    1.765696e-10, 1.780948e-10, 1.757081e-10, 1.764256e-10, 1.769251e-10, 
    1.767062e-10, 1.77845e-10, 1.781136e-10, 1.792061e-10, 1.786412e-10, 
    1.820121e-10, 1.805186e-10, 1.846714e-10, 1.835083e-10, 1.75716e-10, 
    1.760798e-10, 1.773474e-10, 1.76744e-10, 1.784716e-10, 1.788975e-10, 
    1.792441e-10, 1.79687e-10, 1.79735e-10, 1.799976e-10, 1.795673e-10, 
    1.799807e-10, 1.784179e-10, 1.791159e-10, 1.772027e-10, 1.776677e-10, 
    1.774538e-10, 1.772191e-10, 1.779437e-10, 1.787162e-10, 1.787331e-10, 
    1.789809e-10, 1.796791e-10, 1.784786e-10, 1.822044e-10, 1.799005e-10, 
    1.764768e-10, 1.771781e-10, 1.772788e-10, 1.770069e-10, 1.788548e-10, 
    1.781846e-10, 1.799912e-10, 1.795026e-10, 1.803035e-10, 1.799054e-10, 
    1.798468e-10, 1.793359e-10, 1.790179e-10, 1.782152e-10, 1.77563e-10, 
    1.770464e-10, 1.771665e-10, 1.777341e-10, 1.787636e-10, 1.797392e-10, 
    1.795253e-10, 1.802426e-10, 1.783462e-10, 1.791406e-10, 1.788333e-10, 
    1.796348e-10, 1.778802e-10, 1.79373e-10, 1.774991e-10, 1.776632e-10, 
    1.781713e-10, 1.791942e-10, 1.794213e-10, 1.796632e-10, 1.79514e-10, 
    1.787898e-10, 1.786714e-10, 1.78159e-10, 1.780174e-10, 1.776275e-10, 
    1.773047e-10, 1.775996e-10, 1.779093e-10, 1.787902e-10, 1.795849e-10, 
    1.804526e-10, 1.806652e-10, 1.816798e-10, 1.808533e-10, 1.822172e-10, 
    1.810567e-10, 1.830671e-10, 1.794602e-10, 1.810233e-10, 1.781945e-10, 
    1.784988e-10, 1.790491e-10, 1.803137e-10, 1.796311e-10, 1.804297e-10, 
    1.786667e-10, 1.777535e-10, 1.775178e-10, 1.770777e-10, 1.775279e-10, 
    1.774913e-10, 1.779223e-10, 1.777838e-10, 1.788195e-10, 1.78263e-10, 
    1.798452e-10, 1.804235e-10, 1.820595e-10, 1.83064e-10, 1.840887e-10, 
    1.845413e-10, 1.846791e-10, 1.847368e-10,
  1.861917e-10, 1.871851e-10, 1.869919e-10, 1.87794e-10, 1.87349e-10, 
    1.878744e-10, 1.863931e-10, 1.872245e-10, 1.866936e-10, 1.862812e-10, 
    1.893535e-10, 1.878299e-10, 1.909416e-10, 1.899666e-10, 1.924192e-10, 
    1.907896e-10, 1.927484e-10, 1.923725e-10, 1.935054e-10, 1.931807e-10, 
    1.946315e-10, 1.936554e-10, 1.953854e-10, 1.943985e-10, 1.945526e-10, 
    1.936232e-10, 1.881364e-10, 1.891635e-10, 1.880756e-10, 1.882219e-10, 
    1.881563e-10, 1.873581e-10, 1.869561e-10, 1.86116e-10, 1.862685e-10, 
    1.868857e-10, 1.882877e-10, 1.878116e-10, 1.890129e-10, 1.889857e-10, 
    1.903258e-10, 1.897212e-10, 1.919783e-10, 1.91336e-10, 1.931942e-10, 
    1.927263e-10, 1.931722e-10, 1.93037e-10, 1.931739e-10, 1.924879e-10, 
    1.927817e-10, 1.921785e-10, 1.898343e-10, 1.905222e-10, 1.884729e-10, 
    1.872437e-10, 1.864295e-10, 1.858522e-10, 1.859337e-10, 1.860892e-10, 
    1.868893e-10, 1.876428e-10, 1.882176e-10, 1.886024e-10, 1.889818e-10, 
    1.901311e-10, 1.907409e-10, 1.921081e-10, 1.918614e-10, 1.922796e-10, 
    1.926798e-10, 1.933519e-10, 1.932413e-10, 1.935375e-10, 1.922688e-10, 
    1.931116e-10, 1.917209e-10, 1.921009e-10, 1.890841e-10, 1.879401e-10, 
    1.874537e-10, 1.87029e-10, 1.859965e-10, 1.867092e-10, 1.864281e-10, 
    1.870974e-10, 1.875229e-10, 1.873124e-10, 1.886129e-10, 1.881069e-10, 
    1.907771e-10, 1.896255e-10, 1.926331e-10, 1.919121e-10, 1.928061e-10, 
    1.923498e-10, 1.931318e-10, 1.92428e-10, 1.936479e-10, 1.939137e-10, 
    1.93732e-10, 1.944306e-10, 1.923889e-10, 1.931721e-10, 1.873065e-10, 
    1.873408e-10, 1.875008e-10, 1.867978e-10, 1.867549e-10, 1.861118e-10, 
    1.866841e-10, 1.869279e-10, 1.875476e-10, 1.879144e-10, 1.882633e-10, 
    1.890311e-10, 1.898898e-10, 1.910928e-10, 1.919588e-10, 1.925399e-10, 
    1.921836e-10, 1.924981e-10, 1.921465e-10, 1.919817e-10, 1.93814e-10, 
    1.927844e-10, 1.943301e-10, 1.942445e-10, 1.935445e-10, 1.942541e-10, 
    1.873649e-10, 1.871675e-10, 1.864821e-10, 1.870184e-10, 1.860418e-10, 
    1.865881e-10, 1.869024e-10, 1.881173e-10, 1.883848e-10, 1.886327e-10, 
    1.891227e-10, 1.897521e-10, 1.908579e-10, 1.918217e-10, 1.927031e-10, 
    1.926385e-10, 1.926613e-10, 1.928582e-10, 1.923703e-10, 1.929384e-10, 
    1.930337e-10, 1.927844e-10, 1.94233e-10, 1.938188e-10, 1.942427e-10, 
    1.93973e-10, 1.872317e-10, 1.87564e-10, 1.873844e-10, 1.877222e-10, 
    1.874841e-10, 1.885433e-10, 1.888612e-10, 1.903515e-10, 1.897397e-10, 
    1.90714e-10, 1.898386e-10, 1.899936e-10, 1.907454e-10, 1.89886e-10, 
    1.917684e-10, 1.904912e-10, 1.928659e-10, 1.915878e-10, 1.92946e-10, 
    1.926993e-10, 1.93108e-10, 1.934741e-10, 1.939352e-10, 1.947866e-10, 
    1.945894e-10, 1.953022e-10, 1.8806e-10, 1.884917e-10, 1.884539e-10, 
    1.889061e-10, 1.892407e-10, 1.899669e-10, 1.911333e-10, 1.906945e-10, 
    1.915005e-10, 1.916624e-10, 1.90438e-10, 1.911893e-10, 1.887809e-10, 
    1.891692e-10, 1.889381e-10, 1.88094e-10, 1.907953e-10, 1.894073e-10, 
    1.919731e-10, 1.912193e-10, 1.934218e-10, 1.923253e-10, 1.944808e-10, 
    1.954041e-10, 1.962751e-10, 1.972936e-10, 1.887276e-10, 1.884341e-10, 
    1.889599e-10, 1.896879e-10, 1.903646e-10, 1.912652e-10, 1.913575e-10, 
    1.915264e-10, 1.919641e-10, 1.923324e-10, 1.915796e-10, 1.924247e-10, 
    1.892589e-10, 1.90916e-10, 1.883231e-10, 1.891024e-10, 1.89645e-10, 
    1.894071e-10, 1.906444e-10, 1.909363e-10, 1.92124e-10, 1.915098e-10, 
    1.951759e-10, 1.935512e-10, 1.980708e-10, 1.968044e-10, 1.883316e-10, 
    1.887267e-10, 1.901038e-10, 1.894482e-10, 1.913255e-10, 1.917884e-10, 
    1.921651e-10, 1.926467e-10, 1.926989e-10, 1.929845e-10, 1.925165e-10, 
    1.92966e-10, 1.912671e-10, 1.920258e-10, 1.899464e-10, 1.904518e-10, 
    1.902193e-10, 1.899643e-10, 1.907517e-10, 1.915914e-10, 1.916096e-10, 
    1.918791e-10, 1.926385e-10, 1.913331e-10, 1.953854e-10, 1.928791e-10, 
    1.891579e-10, 1.899199e-10, 1.900292e-10, 1.897338e-10, 1.917419e-10, 
    1.910135e-10, 1.929776e-10, 1.924462e-10, 1.933172e-10, 1.928842e-10, 
    1.928205e-10, 1.922649e-10, 1.919192e-10, 1.910468e-10, 1.90338e-10, 
    1.897767e-10, 1.899072e-10, 1.905239e-10, 1.916429e-10, 1.927035e-10, 
    1.92471e-10, 1.932509e-10, 1.911891e-10, 1.920527e-10, 1.917187e-10, 
    1.9259e-10, 1.906827e-10, 1.923056e-10, 1.902685e-10, 1.904469e-10, 
    1.90999e-10, 1.921111e-10, 1.923578e-10, 1.926209e-10, 1.924586e-10, 
    1.916713e-10, 1.915426e-10, 1.909857e-10, 1.908319e-10, 1.904081e-10, 
    1.900573e-10, 1.903777e-10, 1.907143e-10, 1.916718e-10, 1.925358e-10, 
    1.934793e-10, 1.937105e-10, 1.948144e-10, 1.939152e-10, 1.953993e-10, 
    1.941368e-10, 1.963243e-10, 1.924002e-10, 1.941002e-10, 1.910243e-10, 
    1.91355e-10, 1.919533e-10, 1.933284e-10, 1.925859e-10, 1.934544e-10, 
    1.915375e-10, 1.905451e-10, 1.902889e-10, 1.898107e-10, 1.902999e-10, 
    1.902601e-10, 1.907285e-10, 1.905779e-10, 1.917036e-10, 1.910987e-10, 
    1.928188e-10, 1.934476e-10, 1.952274e-10, 1.963207e-10, 1.974361e-10, 
    1.97929e-10, 1.980791e-10, 1.981419e-10,
  1.98294e-10, 1.993742e-10, 1.991641e-10, 2.000367e-10, 1.995525e-10, 
    2.001242e-10, 1.985128e-10, 1.994171e-10, 1.988397e-10, 1.983912e-10, 
    2.017346e-10, 2.000757e-10, 2.034645e-10, 2.02402e-10, 2.050756e-10, 
    2.032989e-10, 2.054347e-10, 2.050245e-10, 2.062606e-10, 2.059062e-10, 
    2.074903e-10, 2.064243e-10, 2.083137e-10, 2.072357e-10, 2.074041e-10, 
    2.063892e-10, 2.004093e-10, 2.015277e-10, 2.00343e-10, 2.005024e-10, 
    2.004309e-10, 1.995625e-10, 1.991253e-10, 1.982116e-10, 1.983774e-10, 
    1.990486e-10, 2.00574e-10, 2.000558e-10, 2.013633e-10, 2.013337e-10, 
    2.027934e-10, 2.021347e-10, 2.045946e-10, 2.038943e-10, 2.05921e-10, 
    2.054105e-10, 2.05897e-10, 2.057494e-10, 2.058989e-10, 2.051504e-10, 
    2.054709e-10, 2.048129e-10, 2.022579e-10, 2.030074e-10, 2.007755e-10, 
    1.994382e-10, 1.985524e-10, 1.979248e-10, 1.980134e-10, 1.981825e-10, 
    1.990525e-10, 1.998721e-10, 2.004976e-10, 2.009164e-10, 2.013295e-10, 
    2.025815e-10, 2.032458e-10, 2.047363e-10, 2.044671e-10, 2.049233e-10, 
    2.053598e-10, 2.060931e-10, 2.059724e-10, 2.062957e-10, 2.049114e-10, 
    2.058309e-10, 2.043138e-10, 2.047283e-10, 2.014413e-10, 2.001956e-10, 
    1.996666e-10, 1.992045e-10, 1.980816e-10, 1.988567e-10, 1.98551e-10, 
    1.992787e-10, 1.997417e-10, 1.995127e-10, 2.009279e-10, 2.003772e-10, 
    2.032852e-10, 2.020305e-10, 2.053088e-10, 2.045224e-10, 2.054975e-10, 
    2.049997e-10, 2.058529e-10, 2.05085e-10, 2.064161e-10, 2.067064e-10, 
    2.06508e-10, 2.072707e-10, 2.050424e-10, 2.058969e-10, 1.995062e-10, 
    1.995436e-10, 1.997176e-10, 1.98953e-10, 1.989063e-10, 1.98207e-10, 
    1.988293e-10, 1.990945e-10, 1.997686e-10, 2.001676e-10, 2.005473e-10, 
    2.013832e-10, 2.023184e-10, 2.036293e-10, 2.045733e-10, 2.052071e-10, 
    2.048184e-10, 2.051615e-10, 2.04778e-10, 2.045983e-10, 2.065976e-10, 
    2.054739e-10, 2.071609e-10, 2.070675e-10, 2.063034e-10, 2.07078e-10, 
    1.995698e-10, 1.99355e-10, 1.986097e-10, 1.991928e-10, 1.981309e-10, 
    1.98725e-10, 1.990668e-10, 2.003885e-10, 2.006796e-10, 2.009494e-10, 
    2.014829e-10, 2.021684e-10, 2.033732e-10, 2.044239e-10, 2.053852e-10, 
    2.053147e-10, 2.053395e-10, 2.055544e-10, 2.050222e-10, 2.056418e-10, 
    2.057459e-10, 2.054738e-10, 2.070549e-10, 2.066027e-10, 2.070655e-10, 
    2.06771e-10, 1.994248e-10, 1.997864e-10, 1.99591e-10, 1.999585e-10, 
    1.996995e-10, 2.008522e-10, 2.011984e-10, 2.028215e-10, 2.021548e-10, 
    2.032164e-10, 2.022626e-10, 2.024315e-10, 2.032508e-10, 2.023142e-10, 
    2.043658e-10, 2.029737e-10, 2.055627e-10, 2.04169e-10, 2.056502e-10, 
    2.05381e-10, 2.058269e-10, 2.062265e-10, 2.067298e-10, 2.076595e-10, 
    2.074441e-10, 2.082228e-10, 2.003261e-10, 2.00796e-10, 2.007547e-10, 
    2.01247e-10, 2.016114e-10, 2.024023e-10, 2.036733e-10, 2.03195e-10, 
    2.040736e-10, 2.042501e-10, 2.029156e-10, 2.037344e-10, 2.011109e-10, 
    2.015337e-10, 2.01282e-10, 2.003631e-10, 2.03305e-10, 2.017929e-10, 
    2.045889e-10, 2.037671e-10, 2.061695e-10, 2.049731e-10, 2.073255e-10, 
    2.083342e-10, 2.09286e-10, 2.103998e-10, 2.010528e-10, 2.007333e-10, 
    2.013057e-10, 2.020985e-10, 2.028356e-10, 2.038171e-10, 2.039177e-10, 
    2.041018e-10, 2.045791e-10, 2.049808e-10, 2.041599e-10, 2.050815e-10, 
    2.016316e-10, 2.034365e-10, 2.006124e-10, 2.014609e-10, 2.020518e-10, 
    2.017926e-10, 2.031404e-10, 2.034586e-10, 2.047535e-10, 2.040837e-10, 
    2.08085e-10, 2.063108e-10, 2.112499e-10, 2.098647e-10, 2.006216e-10, 
    2.010518e-10, 2.025515e-10, 2.018374e-10, 2.038828e-10, 2.043875e-10, 
    2.047983e-10, 2.053237e-10, 2.053806e-10, 2.056922e-10, 2.051816e-10, 
    2.05672e-10, 2.038192e-10, 2.046464e-10, 2.0238e-10, 2.029306e-10, 
    2.026772e-10, 2.023994e-10, 2.032574e-10, 2.041728e-10, 2.041926e-10, 
    2.044865e-10, 2.053152e-10, 2.038911e-10, 2.083141e-10, 2.055777e-10, 
    2.015212e-10, 2.023513e-10, 2.024702e-10, 2.021483e-10, 2.043369e-10, 
    2.035428e-10, 2.056846e-10, 2.051049e-10, 2.060551e-10, 2.055827e-10, 
    2.055132e-10, 2.049072e-10, 2.045302e-10, 2.035791e-10, 2.028066e-10, 
    2.02195e-10, 2.023372e-10, 2.030092e-10, 2.042289e-10, 2.053856e-10, 
    2.05132e-10, 2.059829e-10, 2.037342e-10, 2.046758e-10, 2.043116e-10, 
    2.052618e-10, 2.031823e-10, 2.04952e-10, 2.027309e-10, 2.029252e-10, 
    2.03527e-10, 2.047396e-10, 2.050085e-10, 2.052955e-10, 2.051184e-10, 
    2.0426e-10, 2.041195e-10, 2.035124e-10, 2.033448e-10, 2.028829e-10, 
    2.025008e-10, 2.028499e-10, 2.032167e-10, 2.042604e-10, 2.052027e-10, 
    2.062321e-10, 2.064845e-10, 2.076901e-10, 2.067082e-10, 2.083294e-10, 
    2.069504e-10, 2.0934e-10, 2.05055e-10, 2.069102e-10, 2.035545e-10, 
    2.039149e-10, 2.045674e-10, 2.060676e-10, 2.052573e-10, 2.062051e-10, 
    2.04114e-10, 2.030324e-10, 2.027531e-10, 2.022322e-10, 2.02765e-10, 
    2.027217e-10, 2.032321e-10, 2.03068e-10, 2.042951e-10, 2.036356e-10, 
    2.055114e-10, 2.061977e-10, 2.08141e-10, 2.09336e-10, 2.105555e-10, 
    2.110947e-10, 2.11259e-10, 2.113276e-10,
  2.010817e-10, 2.022192e-10, 2.019978e-10, 2.029173e-10, 2.024069e-10, 
    2.030095e-10, 2.01312e-10, 2.022644e-10, 2.016561e-10, 2.011839e-10, 
    2.047086e-10, 2.029584e-10, 2.065359e-10, 2.05413e-10, 2.082406e-10, 
    2.063609e-10, 2.086208e-10, 2.081863e-10, 2.094958e-10, 2.091202e-10, 
    2.108003e-10, 2.096693e-10, 2.116743e-10, 2.105299e-10, 2.107086e-10, 
    2.096321e-10, 2.0331e-10, 2.044902e-10, 2.032401e-10, 2.034082e-10, 
    2.033328e-10, 2.024175e-10, 2.019571e-10, 2.009949e-10, 2.011694e-10, 
    2.018762e-10, 2.034838e-10, 2.029373e-10, 2.043162e-10, 2.042851e-10, 
    2.058264e-10, 2.051306e-10, 2.077312e-10, 2.069902e-10, 2.091358e-10, 
    2.08595e-10, 2.091104e-10, 2.08954e-10, 2.091124e-10, 2.083196e-10, 
    2.086591e-10, 2.079622e-10, 2.052608e-10, 2.060526e-10, 2.036962e-10, 
    2.022868e-10, 2.013537e-10, 2.006931e-10, 2.007864e-10, 2.009644e-10, 
    2.018803e-10, 2.027437e-10, 2.03403e-10, 2.038448e-10, 2.042806e-10, 
    2.056028e-10, 2.063047e-10, 2.078813e-10, 2.075963e-10, 2.080792e-10, 
    2.085413e-10, 2.093183e-10, 2.091903e-10, 2.09533e-10, 2.080665e-10, 
    2.090405e-10, 2.07434e-10, 2.078727e-10, 2.04399e-10, 2.030846e-10, 
    2.025273e-10, 2.020403e-10, 2.008582e-10, 2.016741e-10, 2.013522e-10, 
    2.021185e-10, 2.026062e-10, 2.023649e-10, 2.038569e-10, 2.032761e-10, 
    2.063464e-10, 2.050207e-10, 2.084873e-10, 2.076548e-10, 2.086872e-10, 
    2.0816e-10, 2.090638e-10, 2.082503e-10, 2.096606e-10, 2.099685e-10, 
    2.097581e-10, 2.105669e-10, 2.082052e-10, 2.091104e-10, 2.023582e-10, 
    2.023975e-10, 2.025808e-10, 2.017756e-10, 2.017263e-10, 2.009901e-10, 
    2.016452e-10, 2.019245e-10, 2.026345e-10, 2.030552e-10, 2.034555e-10, 
    2.043373e-10, 2.053248e-10, 2.067101e-10, 2.077087e-10, 2.083796e-10, 
    2.07968e-10, 2.083313e-10, 2.079252e-10, 2.077351e-10, 2.098531e-10, 
    2.086623e-10, 2.104505e-10, 2.103513e-10, 2.095412e-10, 2.103625e-10, 
    2.024251e-10, 2.021988e-10, 2.014139e-10, 2.02028e-10, 2.0091e-10, 
    2.015353e-10, 2.018954e-10, 2.032882e-10, 2.03595e-10, 2.038796e-10, 
    2.044425e-10, 2.051662e-10, 2.064393e-10, 2.075506e-10, 2.085682e-10, 
    2.084935e-10, 2.085198e-10, 2.087474e-10, 2.081838e-10, 2.088401e-10, 
    2.089503e-10, 2.086621e-10, 2.10338e-10, 2.098585e-10, 2.103492e-10, 
    2.100369e-10, 2.022723e-10, 2.026534e-10, 2.024474e-10, 2.028348e-10, 
    2.025619e-10, 2.037772e-10, 2.041424e-10, 2.058563e-10, 2.051519e-10, 
    2.062736e-10, 2.052657e-10, 2.054441e-10, 2.063102e-10, 2.053201e-10, 
    2.074892e-10, 2.060172e-10, 2.087563e-10, 2.072811e-10, 2.088489e-10, 
    2.085637e-10, 2.090361e-10, 2.094596e-10, 2.099932e-10, 2.109797e-10, 
    2.10751e-10, 2.115776e-10, 2.032222e-10, 2.037179e-10, 2.036742e-10, 
    2.041936e-10, 2.045782e-10, 2.054132e-10, 2.067566e-10, 2.062508e-10, 
    2.071798e-10, 2.073666e-10, 2.059555e-10, 2.068212e-10, 2.0405e-10, 
    2.044963e-10, 2.042305e-10, 2.032613e-10, 2.063673e-10, 2.047699e-10, 
    2.077252e-10, 2.068557e-10, 2.093992e-10, 2.08132e-10, 2.106252e-10, 
    2.116962e-10, 2.127072e-10, 2.138922e-10, 2.039887e-10, 2.036516e-10, 
    2.042554e-10, 2.050925e-10, 2.058711e-10, 2.069086e-10, 2.07015e-10, 
    2.072097e-10, 2.077148e-10, 2.081399e-10, 2.072714e-10, 2.082466e-10, 
    2.045998e-10, 2.065063e-10, 2.035242e-10, 2.044195e-10, 2.050431e-10, 
    2.047695e-10, 2.061931e-10, 2.065294e-10, 2.078995e-10, 2.071906e-10, 
    2.114316e-10, 2.095491e-10, 2.14797e-10, 2.133228e-10, 2.035339e-10, 
    2.039875e-10, 2.055709e-10, 2.048167e-10, 2.06978e-10, 2.07512e-10, 
    2.079467e-10, 2.085031e-10, 2.085633e-10, 2.088934e-10, 2.083526e-10, 
    2.08872e-10, 2.069109e-10, 2.077859e-10, 2.053896e-10, 2.059714e-10, 
    2.057036e-10, 2.054102e-10, 2.063167e-10, 2.07285e-10, 2.073057e-10, 
    2.076168e-10, 2.084947e-10, 2.069868e-10, 2.116752e-10, 2.087726e-10, 
    2.044829e-10, 2.053595e-10, 2.05485e-10, 2.05145e-10, 2.074584e-10, 
    2.066185e-10, 2.088854e-10, 2.082713e-10, 2.09278e-10, 2.087774e-10, 
    2.087038e-10, 2.08062e-10, 2.07663e-10, 2.06657e-10, 2.058404e-10, 
    2.051943e-10, 2.053444e-10, 2.060546e-10, 2.073443e-10, 2.085687e-10, 
    2.083002e-10, 2.092014e-10, 2.068209e-10, 2.078172e-10, 2.074318e-10, 
    2.084375e-10, 2.062374e-10, 2.0811e-10, 2.057603e-10, 2.059657e-10, 
    2.066018e-10, 2.078848e-10, 2.081693e-10, 2.084733e-10, 2.082857e-10, 
    2.073771e-10, 2.072285e-10, 2.065864e-10, 2.064093e-10, 2.05921e-10, 
    2.055172e-10, 2.058861e-10, 2.062739e-10, 2.073775e-10, 2.08375e-10, 
    2.094656e-10, 2.097331e-10, 2.110124e-10, 2.099706e-10, 2.116914e-10, 
    2.102279e-10, 2.127652e-10, 2.082189e-10, 2.101849e-10, 2.066308e-10, 
    2.07012e-10, 2.077026e-10, 2.092914e-10, 2.084328e-10, 2.094371e-10, 
    2.072227e-10, 2.060791e-10, 2.057838e-10, 2.052336e-10, 2.057964e-10, 
    2.057506e-10, 2.0629e-10, 2.061166e-10, 2.074142e-10, 2.067166e-10, 
    2.08702e-10, 2.094292e-10, 2.114909e-10, 2.127605e-10, 2.140576e-10, 
    2.146317e-10, 2.148066e-10, 2.148798e-10,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GC_HEAT1 =
  24786.36, 24802.14, 24799.05, 24811.94, 24804.77, 24813.23, 24789.54, 
    24802.78, 24794.31, 24787.77, 24837.41, 24812.51, 24863.89, 24847.57, 
    24889.16, 24861.33, 24894.82, 24888.34, 24907.9, 24902.26, 24927.74, 
    24910.52, 24941.26, 24923.59, 24926.33, 24909.96, 24817.47, 24834.27, 
    24816.48, 24818.86, 24817.79, 24804.92, 24798.49, 24785.16, 24787.57, 
    24797.36, 24819.93, 24812.21, 24831.77, 24831.32, 24853.55, 24843.49, 
    24881.54, 24870.56, 24902.5, 24894.44, 24902.12, 24899.78, 24902.15, 
    24890.35, 24895.39, 24884.99, 24845.37, 24856.83, 24822.94, 24803.09, 
    24790.12, 24781.01, 24782.29, 24784.74, 24797.42, 24809.49, 24818.78, 
    24825.04, 24831.26, 24850.32, 24860.51, 24883.78, 24879.53, 24886.74, 
    24893.64, 24905.23, 24903.31, 24908.46, 24886.55, 24901.07, 24877.12, 
    24883.65, 24832.96, 24814.29, 24806.46, 24799.65, 24783.28, 24794.56, 
    24790.1, 24800.74, 24807.56, 24804.18, 24825.22, 24816.99, 24861.12, 
    24841.9, 24892.84, 24880.4, 24895.81, 24887.95, 24901.42, 24889.3, 
    24910.39, 24915.04, 24911.86, 24924.16, 24888.63, 24902.12, 24804.09, 
    24804.64, 24807.21, 24795.96, 24795.28, 24785.1, 24794.15, 24798.04, 
    24807.96, 24813.88, 24819.52, 24832.07, 24846.29, 24866.44, 24881.21, 
    24891.24, 24885.08, 24890.52, 24884.44, 24881.6, 24913.29, 24895.44, 
    24922.38, 24920.86, 24908.59, 24921.03, 24805.02, 24801.86, 24790.95, 
    24799.48, 24783.99, 24792.63, 24797.63, 24817.16, 24821.5, 24825.54, 
    24833.58, 24844, 24862.47, 24878.86, 24894.04, 24892.93, 24893.32, 
    24896.7, 24888.31, 24898.08, 24899.73, 24895.43, 24920.66, 24913.38, 
    24920.83, 24916.08, 24802.89, 24808.23, 24805.34, 24810.78, 24806.94, 
    24824.09, 24829.29, 24853.98, 24843.79, 24860.05, 24845.44, 24848.02, 
    24860.59, 24846.23, 24877.95, 24856.32, 24896.84, 24874.86, 24898.21, 
    24893.97, 24901.01, 24907.36, 24915.42, 24930.5, 24926.98, 24939.75, 
    24816.23, 24823.24, 24822.62, 24830.02, 24835.53, 24847.57, 24867.12, 
    24859.72, 24873.36, 24876.12, 24855.42, 24868.07, 24827.97, 24834.35, 
    24830.54, 24816.78, 24861.42, 24838.29, 24881.45, 24868.58, 24906.45, 
    24887.53, 24925.05, 24941.6, 24957.49, 24976.47, 24827.09, 24822.3, 
    24830.9, 24842.94, 24854.2, 24869.36, 24870.93, 24873.8, 24881.3, 
    24887.65, 24874.71, 24889.25, 24835.84, 24863.45, 24820.5, 24833.25, 
    24842.22, 24838.28, 24858.88, 24863.79, 24884.05, 24873.52, 24937.49, 
    24908.71, 24991.23, 24967.3, 24820.63, 24827.08, 24849.85, 24838.96, 
    24870.38, 24878.28, 24884.76, 24893.08, 24893.97, 24898.88, 24890.84, 
    24898.56, 24869.39, 24882.36, 24847.23, 24855.65, 24851.77, 24847.53, 
    24860.68, 24874.92, 24875.22, 24879.84, 24892.96, 24870.51, 24941.28, 
    24897.08, 24834.16, 24846.8, 24848.61, 24843.69, 24877.49, 24865.1, 
    24898.76, 24889.62, 24904.63, 24897.15, 24896.05, 24886.48, 24880.53, 
    24865.66, 24853.75, 24844.41, 24846.58, 24856.86, 24875.79, 24894.05, 
    24890.05, 24903.48, 24868.07, 24882.82, 24877.09, 24892.1, 24859.53, 
    24887.21, 24852.59, 24855.57, 24864.85, 24883.84, 24888.09, 24892.63, 
    24889.84, 24876.28, 24874.08, 24864.62, 24862.03, 24854.92, 24849.07, 
    24854.41, 24860.06, 24876.29, 24891.18, 24907.45, 24911.48, 24931.01, 
    24915.08, 24941.54, 24918.99, 24958.42, 24888.84, 24918.33, 24865.28, 
    24870.88, 24881.12, 24904.83, 24892.03, 24907.02, 24873.99, 24857.22, 
    24852.93, 24844.97, 24853.11, 24852.45, 24860.29, 24857.76, 24876.83, 
    24866.54, 24896.03, 24906.9, 24938.4, 24958.34, 24979.15, 24988.52, 
    24991.39, 24992.59 ;

 GC_ICE1 =
  17951.59, 17976.47, 17971.61, 17991.91, 17980.61, 17993.95, 17956.6, 
    17977.47, 17964.12, 17953.81, 18032.04, 17992.82, 18073.72, 18048.04, 
    18113.48, 18069.69, 18122.37, 18112.19, 18142.89, 18134.04, 18174.01, 
    18146.99, 18195.22, 18167.51, 18171.8, 18146.11, 18000.62, 18027.09, 
    17999.07, 18002.81, 18001.13, 17980.85, 17970.71, 17949.7, 17953.49, 
    17968.94, 18004.49, 17992.35, 18023.15, 18022.45, 18057.45, 18041.61, 
    18101.49, 18084.21, 18134.41, 18121.76, 18133.81, 18130.15, 18133.86, 
    18115.34, 18123.26, 18106.91, 18044.57, 18062.62, 18009.24, 17977.97, 
    17957.51, 17943.16, 17945.18, 17949.04, 17969.03, 17988.06, 18002.69, 
    18012.56, 18022.35, 18052.36, 18068.4, 18105.01, 18098.33, 18109.67, 
    18120.51, 18138.7, 18135.69, 18143.77, 18109.37, 18132.18, 18094.54, 
    18104.81, 18025.04, 17995.61, 17983.28, 17972.54, 17946.73, 17964.51, 
    17957.48, 17974.26, 17985.02, 17979.68, 18012.83, 17999.87, 18069.36, 
    18039.11, 18119.25, 18099.7, 18123.91, 18111.57, 18132.72, 18113.7, 
    18146.79, 18154.09, 18149.1, 18168.39, 18112.64, 18133.82, 17979.54, 
    17980.4, 17984.45, 17966.73, 17965.66, 17949.6, 17963.88, 17970, 
    17985.64, 17994.96, 18003.86, 18023.63, 18046.03, 18077.73, 18100.96, 
    18116.75, 18107.05, 18115.62, 18106.04, 18101.58, 18151.35, 18123.33, 
    18165.6, 18163.23, 18143.96, 18163.49, 17981.01, 17976.02, 17958.82, 
    17972.27, 17947.86, 17961.48, 17969.36, 18000.14, 18006.97, 18013.34, 
    18026, 18042.42, 18071.49, 18097.26, 18121.13, 18119.4, 18120.01, 
    18125.32, 18112.13, 18127.48, 18130.06, 18123.32, 18162.91, 18151.48, 
    18163.18, 18155.72, 17977.64, 17986.06, 17981.51, 17990.08, 17984.04, 
    18011.05, 18019.25, 18058.13, 18042.09, 18067.68, 18044.69, 18048.75, 
    18068.53, 18045.92, 18095.83, 18061.81, 18125.52, 18090.98, 18127.69, 
    18121.03, 18132.07, 18142.04, 18154.68, 18178.34, 18172.82, 18192.86, 
    17998.67, 18009.72, 18008.74, 18020.39, 18029.07, 18048.05, 18078.8, 
    18067.16, 18088.62, 18092.96, 18060.39, 18080.3, 18017.17, 18027.22, 
    18021.22, 17999.54, 18069.84, 18033.42, 18101.35, 18081.1, 18140.61, 
    18110.91, 18169.79, 18195.76, 18220.68, 18250.46, 18015.79, 18008.24, 
    18021.79, 18040.75, 18058.47, 18082.32, 18084.79, 18089.31, 18101.1, 
    18111.1, 18090.75, 18113.61, 18029.57, 18073.03, 18005.39, 18025.49, 
    18039.62, 18033.4, 18065.83, 18073.56, 18105.44, 18088.87, 18189.31, 
    18144.15, 18273.6, 18236.08, 18005.61, 18015.76, 18051.63, 18034.47, 
    18083.93, 18096.36, 18106.55, 18119.62, 18121.02, 18128.73, 18116.12, 
    18128.23, 18082.38, 18102.77, 18047.51, 18060.76, 18054.65, 18047.98, 
    18068.67, 18091.07, 18091.54, 18098.81, 18119.44, 18084.13, 18195.26, 
    18125.92, 18026.92, 18046.83, 18049.68, 18041.94, 18095.11, 18075.62, 
    18128.54, 18114.2, 18137.75, 18126.02, 18124.3, 18109.26, 18099.89, 
    18076.5, 18057.77, 18043.06, 18046.48, 18062.66, 18092.45, 18121.15, 
    18114.88, 18135.95, 18080.29, 18103.5, 18094.49, 18118.1, 18066.85, 
    18110.4, 18055.94, 18060.63, 18075.23, 18105.1, 18111.79, 18118.93, 
    18114.54, 18093.21, 18089.75, 18074.88, 18070.8, 18059.61, 18050.41, 
    18058.81, 18067.69, 18093.22, 18116.64, 18142.18, 18148.5, 18179.14, 
    18154.15, 18195.66, 18160.29, 18222.14, 18112.96, 18159.26, 18075.9, 
    18084.72, 18100.82, 18138.07, 18117.99, 18141.51, 18089.61, 18063.22, 
    18056.47, 18043.95, 18056.76, 18055.72, 18068.05, 18064.08, 18094.08, 
    18077.88, 18124.26, 18141.32, 18190.75, 18222.02, 18254.65, 18269.34, 
    18273.84, 18275.73 ;

 GC_LIQ1 =
  5291.727, 5293.509, 5293.16, 5294.615, 5293.805, 5294.762, 5292.086, 
    5293.58, 5292.624, 5291.886, 5297.501, 5294.68, 5300.52, 5298.655, 
    5303.409, 5300.228, 5304.064, 5303.316, 5305.585, 5304.93, 5307.894, 
    5305.89, 5309.469, 5307.411, 5307.73, 5305.824, 5295.242, 5297.146, 
    5295.13, 5295.399, 5295.278, 5293.822, 5293.096, 5291.592, 5291.863, 
    5292.969, 5295.52, 5294.646, 5296.862, 5296.812, 5299.338, 5298.191, 
    5302.538, 5301.282, 5304.957, 5304.019, 5304.913, 5304.641, 5304.916, 
    5303.545, 5304.13, 5302.932, 5298.405, 5299.713, 5295.861, 5293.616, 
    5292.151, 5291.125, 5291.269, 5291.545, 5292.975, 5294.339, 5295.391, 
    5296.1, 5296.805, 5298.969, 5300.133, 5302.794, 5302.308, 5303.132, 
    5303.926, 5305.275, 5305.052, 5305.65, 5303.11, 5304.791, 5302.033, 
    5302.779, 5296.998, 5294.881, 5293.996, 5293.227, 5291.38, 5292.652, 
    5292.148, 5293.35, 5294.121, 5293.739, 5296.12, 5295.187, 5300.203, 
    5298.011, 5303.833, 5302.408, 5304.178, 5303.271, 5304.832, 5303.426, 
    5305.875, 5306.416, 5306.045, 5307.477, 5303.348, 5304.913, 5293.728, 
    5293.79, 5294.08, 5292.811, 5292.733, 5291.585, 5292.606, 5293.044, 
    5294.166, 5294.834, 5295.475, 5296.897, 5298.51, 5300.812, 5302.5, 
    5303.648, 5302.942, 5303.565, 5302.869, 5302.544, 5306.213, 5304.135, 
    5307.27, 5307.094, 5305.665, 5307.113, 5293.834, 5293.476, 5292.245, 
    5293.207, 5291.46, 5292.435, 5292.999, 5295.207, 5295.698, 5296.157, 
    5297.067, 5298.25, 5300.358, 5302.23, 5303.973, 5303.844, 5303.889, 
    5304.283, 5303.312, 5304.443, 5304.634, 5304.135, 5307.07, 5306.222, 
    5307.09, 5306.537, 5293.592, 5294.195, 5293.869, 5294.483, 5294.05, 
    5295.992, 5296.581, 5299.388, 5298.226, 5300.082, 5298.413, 5298.707, 
    5300.143, 5298.502, 5302.126, 5299.655, 5304.298, 5301.774, 5304.458, 
    5303.965, 5304.783, 5305.522, 5306.459, 5308.215, 5307.806, 5309.293, 
    5295.101, 5295.896, 5295.826, 5296.664, 5297.288, 5298.655, 5300.89, 
    5300.043, 5301.602, 5301.918, 5299.552, 5300.998, 5296.432, 5297.155, 
    5296.724, 5295.164, 5300.238, 5297.601, 5302.527, 5301.056, 5305.417, 
    5303.223, 5307.581, 5309.509, 5311.36, 5313.573, 5296.333, 5295.789, 
    5296.764, 5298.129, 5299.412, 5301.145, 5301.324, 5301.653, 5302.51, 
    5303.236, 5301.757, 5303.419, 5297.324, 5300.47, 5295.585, 5297.031, 
    5298.048, 5297.6, 5299.947, 5300.509, 5302.825, 5301.621, 5309.029, 
    5305.679, 5315.295, 5312.504, 5295.6, 5296.331, 5298.916, 5297.677, 
    5301.262, 5302.165, 5302.905, 5303.861, 5303.964, 5304.536, 5303.602, 
    5304.499, 5301.149, 5302.631, 5298.617, 5299.579, 5299.135, 5298.65, 
    5300.153, 5301.78, 5301.815, 5302.343, 5303.847, 5301.276, 5309.471, 
    5304.327, 5297.133, 5298.567, 5298.774, 5298.214, 5302.074, 5300.658, 
    5304.521, 5303.462, 5305.205, 5304.334, 5304.207, 5303.103, 5302.422, 
    5300.722, 5299.361, 5298.295, 5298.542, 5299.717, 5301.881, 5303.974, 
    5303.511, 5305.071, 5300.998, 5302.685, 5302.029, 5303.748, 5300.021, 
    5303.186, 5299.229, 5299.569, 5300.63, 5302.8, 5303.287, 5303.809, 
    5303.486, 5301.936, 5301.685, 5300.604, 5300.308, 5299.495, 5298.827, 
    5299.437, 5300.082, 5301.937, 5303.64, 5305.533, 5306.001, 5308.274, 
    5306.42, 5309.5, 5306.876, 5311.468, 5303.372, 5306.799, 5300.678, 
    5301.319, 5302.489, 5305.228, 5303.739, 5305.483, 5301.675, 5299.758, 
    5299.268, 5298.36, 5299.288, 5299.212, 5300.108, 5299.82, 5301.999, 
    5300.822, 5304.204, 5305.469, 5309.136, 5311.459, 5313.885, 5314.978, 
    5315.313, 5315.454 ;

 GPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GROSS_NMIN =
  1.074113e-08, 1.077053e-08, 1.076482e-08, 1.078852e-08, 1.077538e-08, 
    1.079089e-08, 1.074709e-08, 1.07717e-08, 1.075599e-08, 1.074378e-08, 
    1.08345e-08, 1.078958e-08, 1.088117e-08, 1.085253e-08, 1.092447e-08, 
    1.087671e-08, 1.09341e-08, 1.09231e-08, 1.095621e-08, 1.094673e-08, 
    1.098906e-08, 1.096059e-08, 1.101101e-08, 1.098227e-08, 1.098676e-08, 
    1.095965e-08, 1.079863e-08, 1.082891e-08, 1.079683e-08, 1.080115e-08, 
    1.079921e-08, 1.077565e-08, 1.076376e-08, 1.073889e-08, 1.074341e-08, 
    1.076168e-08, 1.080309e-08, 1.078904e-08, 1.082446e-08, 1.082367e-08, 
    1.086309e-08, 1.084531e-08, 1.091156e-08, 1.089274e-08, 1.094712e-08, 
    1.093345e-08, 1.094648e-08, 1.094253e-08, 1.094653e-08, 1.092647e-08, 
    1.093507e-08, 1.091742e-08, 1.084864e-08, 1.086886e-08, 1.080855e-08, 
    1.077227e-08, 1.074817e-08, 1.073107e-08, 1.073349e-08, 1.07381e-08, 
    1.076178e-08, 1.078405e-08, 1.080102e-08, 1.081237e-08, 1.082355e-08, 
    1.085737e-08, 1.087528e-08, 1.091536e-08, 1.090813e-08, 1.092038e-08, 
    1.093209e-08, 1.095173e-08, 1.09485e-08, 1.095715e-08, 1.092006e-08, 
    1.094471e-08, 1.090402e-08, 1.091515e-08, 1.082657e-08, 1.079283e-08, 
    1.077847e-08, 1.076592e-08, 1.073535e-08, 1.075646e-08, 1.074813e-08, 
    1.076793e-08, 1.078051e-08, 1.077429e-08, 1.081268e-08, 1.079776e-08, 
    1.087634e-08, 1.08425e-08, 1.093072e-08, 1.090962e-08, 1.093578e-08, 
    1.092243e-08, 1.09453e-08, 1.092472e-08, 1.096037e-08, 1.096813e-08, 
    1.096283e-08, 1.09832e-08, 1.092358e-08, 1.094648e-08, 1.077412e-08, 
    1.077513e-08, 1.077986e-08, 1.075908e-08, 1.075781e-08, 1.073876e-08, 
    1.075571e-08, 1.076292e-08, 1.078124e-08, 1.079207e-08, 1.080237e-08, 
    1.0825e-08, 1.085028e-08, 1.088561e-08, 1.091099e-08, 1.092799e-08, 
    1.091757e-08, 1.092677e-08, 1.091648e-08, 1.091166e-08, 1.096522e-08, 
    1.093515e-08, 1.098027e-08, 1.097778e-08, 1.095736e-08, 1.097806e-08, 
    1.077584e-08, 1.077001e-08, 1.074973e-08, 1.07656e-08, 1.073669e-08, 
    1.075287e-08, 1.076217e-08, 1.079806e-08, 1.080595e-08, 1.081326e-08, 
    1.08277e-08, 1.084622e-08, 1.087871e-08, 1.090697e-08, 1.093277e-08, 
    1.093088e-08, 1.093154e-08, 1.09373e-08, 1.092303e-08, 1.093965e-08, 
    1.094243e-08, 1.093515e-08, 1.097744e-08, 1.096536e-08, 1.097772e-08, 
    1.096986e-08, 1.07719e-08, 1.078173e-08, 1.077642e-08, 1.07864e-08, 
    1.077937e-08, 1.081063e-08, 1.082e-08, 1.086385e-08, 1.084586e-08, 
    1.087449e-08, 1.084877e-08, 1.085333e-08, 1.087542e-08, 1.085016e-08, 
    1.090541e-08, 1.086795e-08, 1.093753e-08, 1.090012e-08, 1.093987e-08, 
    1.093266e-08, 1.09446e-08, 1.09553e-08, 1.096876e-08, 1.099358e-08, 
    1.098783e-08, 1.100859e-08, 1.079637e-08, 1.080911e-08, 1.080799e-08, 
    1.082132e-08, 1.083118e-08, 1.085254e-08, 1.088679e-08, 1.087391e-08, 
    1.089756e-08, 1.09023e-08, 1.086638e-08, 1.088844e-08, 1.081763e-08, 
    1.082907e-08, 1.082226e-08, 1.079738e-08, 1.087688e-08, 1.083608e-08, 
    1.091141e-08, 1.088931e-08, 1.095377e-08, 1.092172e-08, 1.098467e-08, 
    1.101156e-08, 1.103688e-08, 1.106644e-08, 1.081606e-08, 1.080741e-08, 
    1.082291e-08, 1.084434e-08, 1.086423e-08, 1.089066e-08, 1.089337e-08, 
    1.089832e-08, 1.091114e-08, 1.092192e-08, 1.089988e-08, 1.092463e-08, 
    1.083172e-08, 1.088042e-08, 1.080413e-08, 1.082711e-08, 1.084308e-08, 
    1.083607e-08, 1.087244e-08, 1.088101e-08, 1.091582e-08, 1.089783e-08, 
    1.100492e-08, 1.095755e-08, 1.108895e-08, 1.105225e-08, 1.080438e-08, 
    1.081603e-08, 1.085657e-08, 1.083728e-08, 1.089243e-08, 1.0906e-08, 
    1.091703e-08, 1.093112e-08, 1.093265e-08, 1.094099e-08, 1.092731e-08, 
    1.094046e-08, 1.089072e-08, 1.091295e-08, 1.085194e-08, 1.086679e-08, 
    1.085996e-08, 1.085246e-08, 1.087559e-08, 1.090023e-08, 1.090076e-08, 
    1.090865e-08, 1.093089e-08, 1.089265e-08, 1.101102e-08, 1.093793e-08, 
    1.082874e-08, 1.085116e-08, 1.085437e-08, 1.084568e-08, 1.090463e-08, 
    1.088328e-08, 1.094079e-08, 1.092525e-08, 1.095071e-08, 1.093806e-08, 
    1.09362e-08, 1.091995e-08, 1.090983e-08, 1.088426e-08, 1.086345e-08, 
    1.084694e-08, 1.085078e-08, 1.086891e-08, 1.090173e-08, 1.093278e-08, 
    1.092598e-08, 1.094878e-08, 1.088843e-08, 1.091374e-08, 1.090396e-08, 
    1.092946e-08, 1.087357e-08, 1.092115e-08, 1.08614e-08, 1.086664e-08, 
    1.088285e-08, 1.091545e-08, 1.092267e-08, 1.093037e-08, 1.092562e-08, 
    1.090257e-08, 1.089879e-08, 1.088246e-08, 1.087795e-08, 1.08655e-08, 
    1.08552e-08, 1.086461e-08, 1.08745e-08, 1.090258e-08, 1.092788e-08, 
    1.095545e-08, 1.09622e-08, 1.099439e-08, 1.096818e-08, 1.101143e-08, 
    1.097465e-08, 1.103831e-08, 1.092392e-08, 1.097358e-08, 1.088359e-08, 
    1.089329e-08, 1.091083e-08, 1.095105e-08, 1.092934e-08, 1.095473e-08, 
    1.089865e-08, 1.086953e-08, 1.0862e-08, 1.084795e-08, 1.086233e-08, 
    1.086116e-08, 1.087491e-08, 1.087049e-08, 1.090351e-08, 1.088578e-08, 
    1.093615e-08, 1.095453e-08, 1.100641e-08, 1.103821e-08, 1.107056e-08, 
    1.108485e-08, 1.108919e-08, 1.109101e-08 ;

 H2OCAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO_TOP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSOI =
  6.431451, 6.459606, 6.454126, 6.476879, 6.464251, 6.479159, 6.437151, 
    6.460727, 6.44567, 6.43398, 6.521176, 6.477895, 6.5663, 6.538567, 
    6.60836, 6.561982, 6.617734, 6.607016, 6.639297, 6.630039, 6.671434, 
    6.643571, 6.692944, 6.664772, 6.669176, 6.642654, 6.486588, 6.515779, 
    6.484862, 6.489019, 6.487153, 6.464512, 6.453123, 6.429299, 6.43362, 
    6.451118, 6.490889, 6.47737, 6.511466, 6.510695, 6.548778, 6.531591, 
    6.595793, 6.577507, 6.630425, 6.617095, 6.629799, 6.625945, 6.629849, 
    6.610305, 6.618675, 6.60149, 6.534808, 6.554366, 6.49614, 6.461283, 
    6.438185, 6.421827, 6.424138, 6.428545, 6.451221, 6.472581, 6.488889, 
    6.499811, 6.510583, 6.543264, 6.560593, 6.599496, 6.592463, 6.604378, 
    6.615769, 6.634923, 6.631768, 6.640215, 6.604062, 6.628078, 6.588459, 
    6.599281, 6.513526, 6.481015, 6.467235, 6.45518, 6.425915, 6.446117, 
    6.438149, 6.457112, 6.469181, 6.46321, 6.50011, 6.48575, 6.561621, 
    6.528876, 6.61444, 6.593905, 6.619367, 6.606367, 6.628652, 6.608593, 
    6.643359, 6.650945, 6.645761, 6.665683, 6.607483, 6.6298, 6.463043, 
    6.464016, 6.468553, 6.448628, 6.44741, 6.429182, 6.445398, 6.452312, 
    6.46988, 6.480287, 6.490188, 6.511989, 6.536389, 6.570597, 6.595235, 
    6.611782, 6.601632, 6.610592, 6.600577, 6.595885, 6.648103, 6.618753, 
    6.662815, 6.660372, 6.640416, 6.660647, 6.4647, 6.459098, 6.439675, 
    6.454873, 6.427198, 6.442682, 6.451595, 6.486053, 6.493635, 6.500674, 
    6.514587, 6.53247, 6.563911, 6.591338, 6.616432, 6.614591, 6.615239, 
    6.620853, 6.606954, 6.623137, 6.625855, 6.618749, 6.660045, 6.648232, 
    6.66032, 6.652627, 6.460918, 6.470347, 6.465251, 6.474836, 6.468084, 
    6.498145, 6.507174, 6.54952, 6.532118, 6.559822, 6.534928, 6.539336, 
    6.560732, 6.536272, 6.589827, 6.553494, 6.621071, 6.584694, 6.623355, 
    6.616323, 6.627966, 6.638406, 6.651551, 6.675848, 6.670216, 6.690562, 
    6.484417, 6.496676, 6.495595, 6.508435, 6.517941, 6.538572, 6.571743, 
    6.559257, 6.582188, 6.586798, 6.551963, 6.57334, 6.504887, 6.51592, 
    6.509347, 6.485385, 6.562136, 6.522682, 6.595644, 6.574189, 6.636918, 
    6.60568, 6.667118, 6.693488, 6.718348, 6.747479, 6.50337, 6.495034, 
    6.509962, 6.530654, 6.549881, 6.575497, 6.578119, 6.582927, 6.595385, 
    6.605872, 6.584449, 6.608502, 6.518485, 6.565567, 6.491886, 6.514024, 
    6.529432, 6.522668, 6.55783, 6.566135, 6.599944, 6.582453, 6.686976, 
    6.640616, 6.7697, 6.733487, 6.492124, 6.50334, 6.54247, 6.523835, 
    6.577208, 6.590385, 6.601107, 6.614831, 6.616312, 6.624452, 6.611116, 
    6.623924, 6.575551, 6.597142, 6.537988, 6.552359, 6.545744, 6.538496, 
    6.560883, 6.584787, 6.585294, 6.592971, 6.614637, 6.577424, 6.69298, 
    6.621485, 6.515584, 6.537251, 6.540345, 6.531945, 6.589063, 6.568334, 
    6.624253, 6.609112, 6.633929, 6.621591, 6.619777, 6.603951, 6.59411, 
    6.569284, 6.549125, 6.533163, 6.536872, 6.554413, 6.58625, 6.616447, 
    6.609826, 6.632041, 6.573329, 6.597913, 6.588406, 6.613211, 6.558927, 
    6.605148, 6.547143, 6.552217, 6.567923, 6.599585, 6.606596, 6.614094, 
    6.609467, 6.587059, 6.58339, 6.56754, 6.56317, 6.551112, 6.54114, 
    6.550251, 6.559828, 6.587066, 6.611671, 6.638556, 6.645143, 6.676661, 
    6.651002, 6.69338, 6.657349, 6.719786, 6.607827, 6.656284, 6.568637, 
    6.578046, 6.595088, 6.634265, 6.613094, 6.637856, 6.583246, 6.55502, 
    6.547725, 6.534133, 6.548036, 6.546904, 6.560223, 6.555941, 6.587972, 
    6.570755, 6.619732, 6.637659, 6.688429, 6.719665, 6.751538, 6.765638, 
    6.769933, 6.771729,
  4.808921, 4.825948, 4.822634, 4.836389, 4.828754, 4.837767, 4.812368, 
    4.826627, 4.817521, 4.81045, 4.863151, 4.837003, 4.890371, 4.873639, 
    4.915723, 4.887769, 4.921369, 4.91491, 4.934351, 4.928777, 4.953697, 
    4.936924, 4.966632, 4.949686, 4.952337, 4.936372, 4.842254, 4.859892, 
    4.841211, 4.843724, 4.842595, 4.828914, 4.822031, 4.807618, 4.810232, 
    4.820817, 4.844853, 4.836683, 4.857279, 4.856813, 4.8798, 4.869429, 
    4.908148, 4.897126, 4.929009, 4.920981, 4.928633, 4.926311, 4.928663, 
    4.916892, 4.921934, 4.911581, 4.871371, 4.883172, 4.848025, 4.826966, 
    4.812994, 4.803097, 4.804495, 4.807163, 4.820879, 4.83379, 4.843643, 
    4.850241, 4.856746, 4.876479, 4.88693, 4.910381, 4.90614, 4.913322, 
    4.920183, 4.931718, 4.929818, 4.934905, 4.91313, 4.927598, 4.903727, 
    4.91025, 4.858532, 4.838886, 4.830563, 4.823272, 4.805571, 4.817792, 
    4.812973, 4.824439, 4.831735, 4.828125, 4.850421, 4.841747, 4.887549, 
    4.867792, 4.919383, 4.90701, 4.92235, 4.914518, 4.927943, 4.91586, 
    4.936797, 4.941365, 4.938244, 4.950232, 4.915191, 4.928635, 4.828024, 
    4.828613, 4.831355, 4.819311, 4.818573, 4.807547, 4.817356, 4.821538, 
    4.832156, 4.838446, 4.844429, 4.857595, 4.872327, 4.892962, 4.907812, 
    4.917781, 4.911665, 4.917064, 4.91103, 4.908202, 4.939654, 4.921982, 
    4.948507, 4.947037, 4.935027, 4.947202, 4.829026, 4.825639, 4.813895, 
    4.823085, 4.806347, 4.815714, 4.821106, 4.841932, 4.84651, 4.850763, 
    4.859164, 4.869959, 4.888929, 4.905464, 4.920582, 4.919473, 4.919863, 
    4.923245, 4.914873, 4.924621, 4.926259, 4.921978, 4.94684, 4.93973, 
    4.947005, 4.942375, 4.82674, 4.832439, 4.82936, 4.835153, 4.831072, 
    4.849238, 4.854692, 4.88025, 4.869748, 4.886463, 4.871443, 4.874104, 
    4.887016, 4.872252, 4.904555, 4.882649, 4.923377, 4.901464, 4.924752, 
    4.920516, 4.927529, 4.933816, 4.941728, 4.956349, 4.95296, 4.965199, 
    4.840942, 4.84835, 4.847694, 4.855449, 4.86119, 4.873641, 4.893651, 
    4.88612, 4.899947, 4.902726, 4.88172, 4.894615, 4.853308, 4.859972, 
    4.856001, 4.841528, 4.88786, 4.864054, 4.908058, 4.895125, 4.93292, 
    4.914108, 4.951097, 4.966962, 4.981902, 4.999408, 4.852391, 4.847355, 
    4.856371, 4.868865, 4.880465, 4.895914, 4.897494, 4.900393, 4.907901, 
    4.91422, 4.901313, 4.915805, 4.861525, 4.889927, 4.845455, 4.858828, 
    4.868127, 4.864043, 4.885259, 4.890268, 4.910651, 4.900106, 4.963047, 
    4.935149, 5.012747, 4.991002, 4.845597, 4.852372, 4.875996, 4.864748, 
    4.896945, 4.904889, 4.911349, 4.919619, 4.92051, 4.925413, 4.91738, 
    4.925095, 4.895947, 4.908961, 4.873288, 4.88196, 4.877968, 4.873595, 
    4.887101, 4.901516, 4.90182, 4.906448, 4.919512, 4.897075, 4.966663, 
    4.923635, 4.859766, 4.872848, 4.874712, 4.869642, 4.904092, 4.891595, 
    4.925293, 4.916173, 4.931119, 4.923689, 4.922597, 4.913063, 4.907134, 
    4.892169, 4.880009, 4.870376, 4.872615, 4.8832, 4.902398, 4.920593, 
    4.916605, 4.929983, 4.894606, 4.909427, 4.903697, 4.918643, 4.885921, 
    4.913794, 4.878812, 4.881873, 4.891347, 4.910436, 4.914657, 4.919175, 
    4.916386, 4.902885, 4.900672, 4.891116, 4.888481, 4.881206, 4.87519, 
    4.880688, 4.886467, 4.902888, 4.917716, 4.933906, 4.937871, 4.956844, 
    4.941403, 4.966904, 4.94523, 4.982774, 4.915404, 4.944583, 4.891777, 
    4.89745, 4.907726, 4.931326, 4.918572, 4.933487, 4.900585, 4.883568, 
    4.879163, 4.870963, 4.879351, 4.878668, 4.886702, 4.884119, 4.903434, 
    4.893054, 4.922571, 4.933368, 4.963917, 4.982696, 5.001841, 5.010307, 
    5.012885, 5.013963,
  4.269209, 4.283816, 4.280973, 4.292773, 4.286224, 4.293955, 4.272167, 
    4.284398, 4.276587, 4.270521, 4.315732, 4.2933, 4.339086, 4.32473, 
    4.360839, 4.336853, 4.365684, 4.360142, 4.376823, 4.37204, 4.393425, 
    4.379032, 4.404526, 4.389983, 4.392258, 4.378558, 4.297804, 4.312936, 
    4.29691, 4.299065, 4.298097, 4.28636, 4.280456, 4.268092, 4.270334, 
    4.279414, 4.300035, 4.293026, 4.310695, 4.310295, 4.330016, 4.321118, 
    4.354339, 4.344882, 4.37224, 4.365351, 4.371917, 4.369925, 4.371943, 
    4.361842, 4.366168, 4.357285, 4.322785, 4.332909, 4.302756, 4.284689, 
    4.272704, 4.264213, 4.265413, 4.267701, 4.279467, 4.290543, 4.298996, 
    4.304657, 4.310238, 4.327167, 4.336133, 4.356255, 4.352616, 4.358779, 
    4.364666, 4.374564, 4.372934, 4.377299, 4.358614, 4.371028, 4.350545, 
    4.356143, 4.311769, 4.294915, 4.287775, 4.28152, 4.266336, 4.276819, 
    4.272685, 4.282521, 4.28878, 4.285684, 4.304811, 4.29737, 4.336665, 
    4.319714, 4.363979, 4.353363, 4.366525, 4.359805, 4.371324, 4.360957, 
    4.378922, 4.382842, 4.380164, 4.390451, 4.360383, 4.371918, 4.285597, 
    4.286102, 4.288454, 4.278122, 4.27749, 4.268031, 4.276445, 4.280033, 
    4.289142, 4.294538, 4.29967, 4.310966, 4.323605, 4.341309, 4.354051, 
    4.362605, 4.357358, 4.36199, 4.356812, 4.354386, 4.381374, 4.36621, 
    4.388971, 4.387709, 4.377403, 4.387851, 4.286457, 4.283551, 4.273477, 
    4.28136, 4.267001, 4.275037, 4.279662, 4.297528, 4.301456, 4.305104, 
    4.312312, 4.321574, 4.337849, 4.352036, 4.365008, 4.364057, 4.364391, 
    4.367294, 4.360109, 4.368474, 4.36988, 4.366206, 4.38754, 4.381439, 
    4.387682, 4.383709, 4.284495, 4.289385, 4.286743, 4.291713, 4.288212, 
    4.303796, 4.308475, 4.330402, 4.321392, 4.335733, 4.322846, 4.325129, 
    4.336207, 4.323541, 4.351256, 4.33246, 4.367406, 4.348603, 4.368587, 
    4.364952, 4.370969, 4.376364, 4.383153, 4.395701, 4.392793, 4.403296, 
    4.296679, 4.303034, 4.302472, 4.309125, 4.31405, 4.324732, 4.3419, 
    4.335439, 4.347302, 4.349687, 4.331664, 4.342727, 4.307288, 4.313005, 
    4.309598, 4.297182, 4.336931, 4.316507, 4.354262, 4.343165, 4.375595, 
    4.359453, 4.391193, 4.404809, 4.417631, 4.432656, 4.306501, 4.302181, 
    4.309916, 4.320635, 4.330587, 4.343842, 4.345198, 4.347685, 4.354127, 
    4.35955, 4.348474, 4.360909, 4.314336, 4.338706, 4.300551, 4.312023, 
    4.320002, 4.316498, 4.3347, 4.338998, 4.356486, 4.347439, 4.401448, 
    4.377508, 4.444106, 4.425441, 4.300673, 4.306485, 4.326752, 4.317102, 
    4.344726, 4.351542, 4.357086, 4.364182, 4.364946, 4.369154, 4.36226, 
    4.36888, 4.34387, 4.355036, 4.32443, 4.33187, 4.328445, 4.324693, 
    4.33628, 4.348649, 4.348909, 4.35288, 4.364089, 4.344838, 4.404551, 
    4.367628, 4.312829, 4.324051, 4.325651, 4.321301, 4.350859, 4.340137, 
    4.369051, 4.361225, 4.374051, 4.367675, 4.366737, 4.358556, 4.353468, 
    4.340629, 4.330196, 4.321931, 4.323852, 4.332933, 4.349405, 4.365017, 
    4.361596, 4.373075, 4.34272, 4.355436, 4.35052, 4.363344, 4.335268, 
    4.359183, 4.329169, 4.331795, 4.339923, 4.356302, 4.359924, 4.363801, 
    4.361408, 4.349823, 4.347925, 4.339725, 4.337464, 4.331223, 4.326061, 
    4.330778, 4.335736, 4.349826, 4.362548, 4.376441, 4.379844, 4.396125, 
    4.382874, 4.404758, 4.386158, 4.418379, 4.360564, 4.385603, 4.340292, 
    4.34516, 4.353977, 4.374227, 4.363284, 4.376081, 4.34785, 4.333249, 
    4.32947, 4.322434, 4.329631, 4.329045, 4.335938, 4.333722, 4.350294, 
    4.341388, 4.366715, 4.375979, 4.402195, 4.418313, 4.434745, 4.442012, 
    4.444225, 4.44515,
  3.964825, 3.978192, 3.975628, 3.986269, 3.980363, 3.987335, 3.967578, 
    3.978716, 3.971674, 3.966046, 4.006982, 3.986744, 4.028073, 4.015109, 
    4.047731, 4.026055, 4.052112, 4.047101, 4.062187, 4.057861, 4.077207, 
    4.064185, 4.087257, 4.074093, 4.076151, 4.063756, 3.990808, 4.004459, 
    3.990001, 3.991945, 3.991072, 3.980486, 3.975161, 3.963785, 3.965872, 
    3.974222, 3.992819, 3.986497, 4.002439, 4.002078, 4.019882, 4.011847, 
    4.041857, 4.03331, 4.058042, 4.051812, 4.057749, 4.055948, 4.057773, 
    4.048639, 4.05255, 4.044519, 4.013352, 4.022494, 3.995275, 3.978978, 
    3.968078, 3.960174, 3.961291, 3.963421, 3.97427, 3.984258, 3.991883, 
    3.99699, 4.002027, 4.017307, 4.025405, 4.043588, 4.0403, 4.045869, 
    4.051192, 4.060143, 4.058669, 4.062617, 4.045721, 4.056945, 4.038428, 
    4.043487, 4.003407, 3.988202, 3.981761, 3.976121, 3.96215, 3.971883, 
    3.96806, 3.977025, 3.982668, 3.979876, 3.99713, 3.990416, 4.025886, 
    4.010579, 4.050571, 4.040974, 4.052874, 4.046798, 4.057213, 4.047839, 
    4.064086, 4.067631, 4.065208, 4.074518, 4.047319, 4.05775, 3.979798, 
    3.980253, 3.982374, 3.973058, 3.972488, 3.963728, 3.971547, 3.974781, 
    3.982995, 3.987861, 3.992491, 4.002684, 4.014091, 4.030081, 4.041596, 
    4.049328, 4.044585, 4.048773, 4.044092, 4.041899, 4.066303, 4.052588, 
    4.073178, 4.072036, 4.062711, 4.072165, 3.980573, 3.977953, 3.968798, 
    3.975977, 3.96277, 3.97025, 3.974446, 3.990558, 3.994102, 3.997394, 
    4.003898, 4.012259, 4.026956, 4.039775, 4.051502, 4.050642, 4.050944, 
    4.053568, 4.047072, 4.054635, 4.055906, 4.052585, 4.071883, 4.066363, 
    4.072012, 4.068417, 3.978804, 3.983214, 3.980831, 3.985313, 3.982156, 
    3.996212, 4.000434, 4.020229, 4.012094, 4.025044, 4.013408, 4.015468, 
    4.025472, 4.014035, 4.039069, 4.022088, 4.05367, 4.036672, 4.054738, 
    4.051451, 4.056892, 4.061771, 4.067914, 4.079268, 4.076636, 4.086143, 
    3.989793, 3.995525, 3.995018, 4.001022, 4.005467, 4.01511, 4.030616, 
    4.02478, 4.035498, 4.037652, 4.02137, 4.031363, 3.999364, 4.004523, 
    4.001449, 3.990246, 4.026127, 4.007684, 4.041787, 4.031759, 4.061076, 
    4.046478, 4.075189, 4.087512, 4.099127, 4.112741, 3.998654, 3.994756, 
    4.001736, 4.011411, 4.020397, 4.032371, 4.033596, 4.035843, 4.041666, 
    4.046566, 4.036556, 4.047796, 4.005724, 4.02773, 3.993285, 4.003637, 
    4.010839, 4.007677, 4.024113, 4.027994, 4.043797, 4.035621, 4.08447, 
    4.062805, 4.123122, 4.106202, 3.993396, 3.99864, 4.016934, 4.008222, 
    4.03317, 4.039329, 4.04434, 4.050754, 4.051446, 4.05525, 4.049017, 
    4.055003, 4.032396, 4.042487, 4.014837, 4.021555, 4.018463, 4.015075, 
    4.025539, 4.036714, 4.03695, 4.040538, 4.050668, 4.033271, 4.087278, 
    4.053868, 4.004364, 4.014495, 4.01594, 4.012013, 4.038712, 4.029023, 
    4.055157, 4.048081, 4.059679, 4.053913, 4.053065, 4.045669, 4.04107, 
    4.029467, 4.020044, 4.012582, 4.014316, 4.022516, 4.037397, 4.05151, 
    4.048416, 4.058796, 4.031357, 4.042848, 4.038405, 4.049997, 4.024625, 
    4.046233, 4.019117, 4.021489, 4.028831, 4.04363, 4.046906, 4.05041, 
    4.048246, 4.037775, 4.03606, 4.028651, 4.026609, 4.020972, 4.016311, 
    4.02057, 4.025047, 4.037778, 4.049277, 4.061841, 4.064919, 4.079651, 
    4.06766, 4.087465, 4.070629, 4.099803, 4.047483, 4.070128, 4.029164, 
    4.033562, 4.041528, 4.059838, 4.049942, 4.061515, 4.035992, 4.0228, 
    4.019389, 4.013036, 4.019534, 4.019005, 4.025231, 4.023229, 4.038201, 
    4.030154, 4.053045, 4.061423, 4.085148, 4.099744, 4.114635, 4.121224, 
    4.12323, 4.12407,
  3.777821, 3.791197, 3.788592, 3.79941, 3.793405, 3.800494, 3.780528, 
    3.79173, 3.784574, 3.779022, 3.820498, 3.799893, 3.841452, 3.828643, 
    3.860905, 3.839457, 3.865245, 3.860282, 3.875235, 3.870944, 3.890142, 
    3.877216, 3.900131, 3.88705, 3.889094, 3.876791, 3.804029, 3.817927, 
    3.803207, 3.805186, 3.804297, 3.793529, 3.788116, 3.776799, 3.778851, 
    3.787163, 3.806075, 3.799643, 3.815871, 3.815504, 3.833358, 3.825423, 
    3.855089, 3.846632, 3.871124, 3.864949, 3.870833, 3.869048, 3.870857, 
    3.861805, 3.86568, 3.857725, 3.826908, 3.835938, 3.808575, 3.791995, 
    3.781019, 3.773252, 3.774349, 3.776441, 3.787212, 3.797366, 3.805124, 
    3.810322, 3.815451, 3.830812, 3.838815, 3.856802, 3.853548, 3.859062, 
    3.864335, 3.873208, 3.871745, 3.87566, 3.858915, 3.870036, 3.851696, 
    3.856703, 3.816854, 3.801377, 3.794824, 3.789093, 3.775192, 3.784787, 
    3.781002, 3.790012, 3.795749, 3.79291, 3.810464, 3.80363, 3.83929, 
    3.824167, 3.863719, 3.854215, 3.866001, 3.859982, 3.870302, 3.861012, 
    3.877118, 3.880635, 3.878232, 3.887472, 3.860498, 3.870834, 3.792831, 
    3.793294, 3.79545, 3.78598, 3.785401, 3.776743, 3.784445, 3.787731, 
    3.796081, 3.801031, 3.805742, 3.816121, 3.827638, 3.843438, 3.854831, 
    3.862489, 3.85779, 3.861938, 3.857302, 3.855131, 3.879318, 3.865717, 
    3.886142, 3.885008, 3.875754, 3.885136, 3.793619, 3.790956, 3.781727, 
    3.788947, 3.775802, 3.783155, 3.78739, 3.803774, 3.807382, 3.810733, 
    3.817358, 3.825829, 3.840348, 3.853028, 3.864641, 3.863789, 3.864089, 
    3.866689, 3.860253, 3.867747, 3.869006, 3.865715, 3.884856, 3.879377, 
    3.884984, 3.881415, 3.791821, 3.796304, 3.793881, 3.798439, 3.795227, 
    3.809529, 3.813828, 3.8337, 3.825667, 3.838459, 3.826964, 3.828998, 
    3.838879, 3.827584, 3.852329, 3.835536, 3.86679, 3.849955, 3.867848, 
    3.864591, 3.869984, 3.874822, 3.880916, 3.89219, 3.889576, 3.899024, 
    3.802996, 3.80883, 3.808315, 3.814428, 3.818956, 3.828645, 3.843967, 
    3.838197, 3.848796, 3.850928, 3.834828, 3.844706, 3.812739, 3.817993, 
    3.814863, 3.803457, 3.839528, 3.821215, 3.85502, 3.845098, 3.874132, 
    3.859664, 3.888138, 3.900384, 3.911941, 3.925501, 3.812016, 3.808048, 
    3.815156, 3.824991, 3.833867, 3.845702, 3.846915, 3.849137, 3.8549, 
    3.859753, 3.849842, 3.86097, 3.819216, 3.841113, 3.80655, 3.817091, 
    3.824428, 3.821208, 3.837538, 3.841375, 3.85701, 3.848918, 3.897359, 
    3.875846, 3.935856, 3.918985, 3.806663, 3.812002, 3.830445, 3.821764, 
    3.846493, 3.852587, 3.857547, 3.8639, 3.864586, 3.868356, 3.86218, 
    3.868112, 3.845727, 3.855713, 3.828376, 3.835011, 3.831957, 3.82861, 
    3.838948, 3.849998, 3.850232, 3.853783, 3.863812, 3.846593, 3.900148, 
    3.866983, 3.817833, 3.828036, 3.829464, 3.825587, 3.851975, 3.842391, 
    3.868264, 3.861253, 3.872747, 3.867031, 3.866191, 3.858864, 3.85431, 
    3.842831, 3.833518, 3.826149, 3.827861, 3.83596, 3.850674, 3.864649, 
    3.861583, 3.871872, 3.8447, 3.85607, 3.851672, 3.86315, 3.838045, 
    3.859419, 3.832603, 3.834945, 3.842201, 3.856844, 3.860088, 3.863559, 
    3.861417, 3.851048, 3.849352, 3.842025, 3.840005, 3.834435, 3.829831, 
    3.834038, 3.838461, 3.851052, 3.862437, 3.874891, 3.877945, 3.892569, 
    3.880662, 3.900334, 3.883607, 3.91261, 3.860658, 3.883112, 3.842531, 
    3.846881, 3.854763, 3.872903, 3.863096, 3.874567, 3.849285, 3.836241, 
    3.832871, 3.826596, 3.833014, 3.832492, 3.838643, 3.836665, 3.85147, 
    3.84351, 3.86617, 3.874476, 3.898033, 3.912553, 3.927391, 3.933962, 
    3.935964, 3.936801,
  3.838219, 3.852606, 3.849802, 3.861416, 3.854983, 3.862548, 3.841128, 
    3.853179, 3.845479, 3.839509, 3.883466, 3.86192, 3.906037, 3.892152, 
    3.92718, 3.903872, 3.931905, 3.926502, 3.942796, 3.938117, 3.959078, 
    3.944958, 3.970011, 3.955697, 3.957932, 3.944494, 3.86624, 3.880774, 
    3.865382, 3.867448, 3.866521, 3.855117, 3.849289, 3.837121, 3.839326, 
    3.848264, 3.868378, 3.86166, 3.878623, 3.878239, 3.897259, 3.888666, 
    3.920852, 3.911661, 3.938312, 3.931583, 3.937996, 3.936049, 3.938021, 
    3.928159, 3.93238, 3.923719, 3.890273, 3.900057, 3.870991, 3.853464, 
    3.841656, 3.833311, 3.834489, 3.836736, 3.848316, 3.85925, 3.867384, 
    3.872818, 3.878184, 3.8945, 3.903176, 3.922715, 3.919177, 3.925174, 
    3.930914, 3.940584, 3.93899, 3.94326, 3.925014, 3.937126, 3.917163, 
    3.922608, 3.87965, 3.86347, 3.856511, 3.850341, 3.835395, 3.845707, 
    3.841637, 3.85133, 3.857508, 3.85445, 3.872967, 3.865823, 3.903692, 
    3.88731, 3.930244, 3.919902, 3.932729, 3.926175, 3.937416, 3.927297, 
    3.94485, 3.94869, 3.946066, 3.95616, 3.926738, 3.937996, 3.854365, 
    3.854863, 3.857186, 3.846991, 3.846368, 3.837061, 3.84534, 3.848875, 
    3.857866, 3.863108, 3.86803, 3.878884, 3.891063, 3.908193, 3.920572, 
    3.928904, 3.923791, 3.928305, 3.92326, 3.920898, 3.947251, 3.93242, 
    3.954705, 3.953467, 3.943362, 3.953606, 3.855213, 3.852346, 3.842417, 
    3.850184, 3.836049, 3.843952, 3.848508, 3.865973, 3.869744, 3.873247, 
    3.88018, 3.889105, 3.90484, 3.918611, 3.931248, 3.93032, 3.930647, 
    3.933479, 3.926471, 3.934631, 3.936004, 3.932417, 3.953301, 3.947316, 
    3.95344, 3.949542, 3.853277, 3.858105, 3.855495, 3.860402, 3.856946, 
    3.871989, 3.876485, 3.89763, 3.888929, 3.90279, 3.890333, 3.892536, 
    3.903246, 3.891005, 3.917851, 3.89962, 3.933589, 3.915271, 3.934741, 
    3.931194, 3.93707, 3.942345, 3.948997, 3.961319, 3.95846, 3.968799, 
    3.865161, 3.871258, 3.870719, 3.877113, 3.881852, 3.892154, 3.908768, 
    3.902507, 3.914012, 3.916328, 3.898854, 3.90957, 3.875345, 3.880844, 
    3.877568, 3.865642, 3.90395, 3.884218, 3.920777, 3.909995, 3.941593, 
    3.925829, 3.956887, 3.970287, 3.98296, 3.997859, 3.87459, 3.870441, 
    3.877874, 3.888197, 3.897811, 3.910652, 3.911969, 3.914383, 3.920647, 
    3.925926, 3.915148, 3.927251, 3.882123, 3.90567, 3.868875, 3.879899, 
    3.887587, 3.884211, 3.901793, 3.905955, 3.922941, 3.914145, 3.966974, 
    3.943462, 4.00926, 3.990695, 3.868993, 3.874575, 3.894104, 3.884793, 
    3.911511, 3.918132, 3.923527, 3.930441, 3.931188, 3.935295, 3.928569, 
    3.935029, 3.910679, 3.921531, 3.891863, 3.899052, 3.895742, 3.892116, 
    3.903322, 3.915318, 3.915573, 3.919432, 3.930343, 3.911619, 3.970028, 
    3.933797, 3.880677, 3.891494, 3.893041, 3.888843, 3.917467, 3.907058, 
    3.935195, 3.927559, 3.940082, 3.933851, 3.932936, 3.924958, 3.920005, 
    3.907534, 3.897433, 3.889451, 3.891304, 3.900081, 3.916053, 3.931257, 
    3.927918, 3.939128, 3.909564, 3.921919, 3.917137, 3.929625, 3.902342, 
    3.925561, 3.896442, 3.898981, 3.906852, 3.92276, 3.926291, 3.93007, 
    3.927737, 3.916459, 3.914616, 3.90666, 3.904468, 3.898428, 3.893438, 
    3.897997, 3.902793, 3.916463, 3.928848, 3.942421, 3.945753, 3.961732, 
    3.948719, 3.970232, 3.951933, 3.983694, 3.92691, 3.951394, 3.90721, 
    3.911932, 3.920497, 3.940252, 3.929566, 3.942067, 3.914543, 3.900385, 
    3.896732, 3.889936, 3.896888, 3.896322, 3.902991, 3.900846, 3.916919, 
    3.908272, 3.932914, 3.941967, 3.967714, 3.983632, 3.999939, 4.007173, 
    4.009379, 4.010302,
  3.964782, 3.983, 3.979443, 3.994247, 3.986019, 3.995736, 3.968459, 
    3.983728, 3.973965, 3.966413, 4.023343, 3.99491, 4.052797, 4.034863, 
    4.080281, 4.049994, 4.086454, 4.079397, 4.100722, 4.094585, 4.122166, 
    4.103562, 4.136641, 4.117702, 4.120652, 4.102952, 4.000594, 4.019778, 
    3.999464, 4.002185, 4.000963, 3.986189, 3.978792, 3.963395, 3.96618, 
    3.977493, 4.00341, 3.994568, 4.016934, 4.016426, 4.041449, 4.030238, 
    4.072033, 4.060087, 4.094841, 4.086032, 4.094426, 4.091876, 4.09446, 
    4.08156, 4.087075, 4.075768, 4.032372, 4.045061, 4.006854, 3.984089, 
    3.969126, 3.958586, 3.960073, 3.96291, 3.97756, 3.991444, 4.0021, 
    4.009264, 4.016353, 4.037889, 4.049094, 4.07446, 4.069852, 4.077664, 
    4.085159, 4.09782, 4.095729, 4.101332, 4.077456, 4.093287, 4.067233, 
    4.074319, 4.018291, 3.996948, 3.987961, 3.980126, 3.961216, 3.974254, 
    3.969103, 3.981381, 3.989228, 3.985342, 4.009461, 4.000045, 4.04976, 
    4.028439, 4.084283, 4.070796, 4.087531, 4.07897, 4.093666, 4.080434, 
    4.103421, 4.108469, 4.105018, 4.118312, 4.079704, 4.094427, 3.985234, 
    3.985867, 3.988819, 3.97588, 3.975091, 3.96332, 3.973789, 3.978267, 
    3.989684, 3.996473, 4.002951, 4.017279, 4.033422, 4.055589, 4.071668, 
    4.082532, 4.075861, 4.081749, 4.075169, 4.072093, 4.106576, 4.087127, 
    4.116394, 4.11476, 4.101465, 4.114944, 3.986312, 3.98267, 3.970089, 
    3.979927, 3.962042, 3.972032, 3.977802, 4.000243, 4.00521, 4.009831, 
    4.018992, 4.030821, 4.051247, 4.069116, 4.085596, 4.084383, 4.084809, 
    4.088512, 4.079356, 4.09002, 4.091817, 4.087123, 4.114542, 4.106663, 
    4.114726, 4.109591, 3.983853, 3.989988, 3.98667, 3.992915, 3.988514, 
    4.00817, 4.014107, 4.041927, 4.030588, 4.048594, 4.032452, 4.035358, 
    4.049184, 4.033343, 4.068127, 4.044497, 4.088656, 4.064774, 4.090164, 
    4.085524, 4.093213, 4.100131, 4.108873, 4.125128, 4.121349, 4.135034, 
    3.999173, 4.007205, 4.006496, 4.014937, 4.021206, 4.034866, 4.056334, 
    4.048229, 4.063138, 4.066148, 4.043508, 4.057374, 4.012601, 4.019871, 
    4.015538, 3.999806, 4.050095, 4.024339, 4.071935, 4.057925, 4.099143, 
    4.078519, 4.119274, 4.137008, 4.153867, 4.173797, 4.011604, 4.006128, 
    4.015943, 4.029617, 4.042161, 4.058777, 4.060485, 4.06362, 4.071765, 
    4.078645, 4.064614, 4.080374, 4.021564, 4.052321, 4.004064, 4.01862, 
    4.028807, 4.02433, 4.047305, 4.05269, 4.074754, 4.063311, 4.132614, 
    4.101598, 4.189129, 4.1642, 4.00422, 4.011584, 4.037378, 4.025102, 
    4.059891, 4.068492, 4.075517, 4.08454, 4.085516, 4.090889, 4.082094, 
    4.09054, 4.058812, 4.072917, 4.034483, 4.043763, 4.03949, 4.034817, 
    4.049283, 4.064834, 4.065166, 4.070184, 4.084412, 4.060032, 4.136664, 
    4.088928, 4.01965, 4.033994, 4.036008, 4.030473, 4.067628, 4.054118, 
    4.090758, 4.080776, 4.097162, 4.088999, 4.087802, 4.077384, 4.07093, 
    4.054736, 4.041673, 4.031281, 4.033742, 4.045092, 4.06579, 4.085606, 
    4.081245, 4.095911, 4.057366, 4.073422, 4.067199, 4.083474, 4.048015, 
    4.078169, 4.040393, 4.043671, 4.053851, 4.074518, 4.079122, 4.084055, 
    4.081009, 4.066318, 4.063922, 4.053603, 4.050766, 4.042957, 4.03652, 
    4.042401, 4.048599, 4.066323, 4.082459, 4.10023, 4.104607, 4.125674, 
    4.108507, 4.136934, 4.11274, 4.154845, 4.07993, 4.112029, 4.054315, 
    4.060438, 4.071571, 4.097384, 4.083397, 4.099765, 4.063828, 4.045485, 
    4.040769, 4.031924, 4.040969, 4.040239, 4.048854, 4.046081, 4.066915, 
    4.055692, 4.087772, 4.099635, 4.133595, 4.154763, 4.176589, 4.186318, 
    4.189291, 4.190535,
  4.394931, 4.425735, 4.419685, 4.444981, 4.430883, 4.447541, 4.401113, 
    4.426975, 4.410401, 4.397671, 4.495614, 4.446121, 4.549213, 4.516021, 
    4.601168, 4.543991, 4.612795, 4.599476, 4.639682, 4.628071, 4.680817, 
    4.64508, 4.709098, 4.672182, 4.677884, 4.643919, 4.455919, 4.489343, 
    4.453968, 4.458671, 4.456557, 4.431174, 4.41858, 4.392606, 4.39728, 
    4.416376, 4.460792, 4.445531, 4.484354, 4.483463, 4.528148, 4.507799, 
    4.585434, 4.562863, 4.628553, 4.612007, 4.627772, 4.622969, 4.627834, 
    4.60362, 4.613957, 4.592544, 4.511585, 4.53483, 4.466766, 4.427591, 
    4.402236, 4.384558, 4.387042, 4.391791, 4.416488, 4.440167, 4.458524, 
    4.470959, 4.483335, 4.521585, 4.542316, 4.590051, 4.581295, 4.596162, 
    4.610373, 4.634184, 4.630231, 4.64084, 4.595766, 4.625624, 4.576335, 
    4.589783, 4.486733, 4.449629, 4.434201, 4.420846, 4.388955, 4.41089, 
    4.402197, 4.422978, 4.43637, 4.429728, 4.471301, 4.454971, 4.543556, 
    4.504612, 4.608737, 4.583086, 4.614812, 4.59866, 4.626339, 4.601462, 
    4.644811, 4.654441, 4.647852, 4.67336, 4.600064, 4.627773, 4.429543, 
    4.430624, 4.435669, 4.413641, 4.412306, 4.392478, 4.410104, 4.417688, 
    4.43715, 4.44881, 4.459997, 4.484957, 4.51345, 4.554431, 4.58474, 
    4.605471, 4.592722, 4.603983, 4.591402, 4.585548, 4.650825, 4.614055, 
    4.669658, 4.666512, 4.641094, 4.666866, 4.431383, 4.425173, 4.403858, 
    4.420507, 4.390338, 4.407135, 4.4169, 4.455313, 4.463913, 4.471945, 
    4.487963, 4.508832, 4.546323, 4.579899, 4.61119, 4.608923, 4.60972, 
    4.616651, 4.599398, 4.61948, 4.622858, 4.614048, 4.666091, 4.65099, 
    4.666445, 4.656587, 4.427188, 4.437671, 4.431995, 4.44269, 4.435147, 
    4.469054, 4.479405, 4.529032, 4.508419, 4.541387, 4.511727, 4.516931, 
    4.542483, 4.51331, 4.578026, 4.533785, 4.616921, 4.571688, 4.619751, 
    4.611056, 4.625486, 4.638561, 4.655214, 4.68657, 4.679235, 4.705936, 
    4.453466, 4.467378, 4.466145, 4.480857, 4.491853, 4.516028, 4.555826, 
    4.540708, 4.568604, 4.574283, 4.531954, 4.557772, 4.476775, 4.489507, 
    4.481909, 4.454559, 4.544178, 4.49737, 4.585248, 4.558807, 4.636689, 
    4.597797, 4.675217, 4.70982, 4.743316, 4.783701, 4.475035, 4.465506, 
    4.482618, 4.506698, 4.529464, 4.560404, 4.563612, 4.569513, 4.584926, 
    4.598039, 4.571387, 4.601347, 4.492483, 4.548326, 4.461925, 4.487311, 
    4.505264, 4.497354, 4.538991, 4.549014, 4.590611, 4.56893, 4.701188, 
    4.641345, 4.815381, 4.764145, 4.462195, 4.475001, 4.520645, 4.498715, 
    4.562496, 4.578719, 4.592064, 4.609218, 4.611042, 4.621113, 4.604644, 
    4.620458, 4.560471, 4.587114, 4.515338, 4.532426, 4.524535, 4.515938, 
    4.542666, 4.571802, 4.572429, 4.581925, 4.608977, 4.562761, 4.709143, 
    4.617431, 4.489119, 4.514466, 4.518125, 4.508215, 4.577083, 4.551682, 
    4.620866, 4.602116, 4.632938, 4.617565, 4.615319, 4.595627, 4.58334, 
    4.552835, 4.528562, 4.509647, 4.514019, 4.534887, 4.573606, 4.611209, 
    4.603016, 4.630574, 4.557758, 4.588075, 4.57627, 4.607226, 4.540309, 
    4.597127, 4.5262, 4.532257, 4.551182, 4.590162, 4.598949, 4.608312, 
    4.602562, 4.574605, 4.570083, 4.550718, 4.545427, 4.530935, 4.519067, 
    4.529907, 4.541395, 4.574615, 4.605334, 4.638749, 4.647069, 4.687633, 
    4.654514, 4.709675, 4.662626, 4.745278, 4.600495, 4.661262, 4.552049, 
    4.563523, 4.584557, 4.633358, 4.607083, 4.637867, 4.569905, 4.535615, 
    4.526893, 4.51079, 4.527263, 4.525915, 4.541871, 4.53672, 4.575733, 
    4.554623, 4.615264, 4.63762, 4.703111, 4.745113, 4.789431, 4.809533, 
    4.815718, 4.818313,
  6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465,
  6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 6.6465, 
    6.6465, 6.6465, 6.6465, 6.6465, 6.6465,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HC =
  25080.9, 25097.14, 25093.96, 25107.21, 25099.84, 25108.55, 25084.17, 
    25097.79, 25089.07, 25082.35, 25133.42, 25107.81, 25160.67, 25143.88, 
    25186.67, 25158.04, 25192.5, 25185.83, 25205.96, 25200.16, 25226.37, 
    25208.65, 25240.29, 25222.1, 25224.92, 25208.07, 25112.9, 25130.19, 
    25111.89, 25114.33, 25113.23, 25099.99, 25093.38, 25079.67, 25082.14, 
    25092.22, 25115.43, 25107.5, 25127.62, 25127.16, 25150.03, 25139.67, 
    25178.83, 25167.53, 25200.4, 25192.1, 25200.01, 25197.6, 25200.04, 
    25187.89, 25193.08, 25182.38, 25141.61, 25153.41, 25118.53, 25098.11, 
    25084.76, 25075.4, 25076.71, 25079.23, 25092.28, 25104.7, 25114.26, 
    25120.7, 25127.1, 25146.7, 25157.19, 25181.13, 25176.76, 25184.18, 
    25191.28, 25203.21, 25201.24, 25206.54, 25183.98, 25198.93, 25174.28, 
    25181, 25128.85, 25109.63, 25101.58, 25094.57, 25077.73, 25089.33, 
    25084.74, 25095.69, 25102.71, 25099.23, 25120.88, 25112.41, 25157.81, 
    25138.04, 25190.46, 25177.66, 25193.51, 25185.43, 25199.29, 25186.82, 
    25208.51, 25213.31, 25210.03, 25222.69, 25186.12, 25200.01, 25099.14, 
    25099.7, 25102.35, 25090.78, 25090.08, 25079.6, 25088.92, 25092.91, 
    25103.12, 25109.21, 25115.02, 25127.93, 25142.56, 25163.29, 25178.48, 
    25188.81, 25182.47, 25188.07, 25181.81, 25178.89, 25211.51, 25193.13, 
    25220.86, 25219.3, 25206.66, 25219.47, 25100.1, 25096.84, 25085.62, 
    25094.39, 25078.46, 25087.35, 25092.5, 25112.59, 25117.05, 25121.21, 
    25129.48, 25140.2, 25159.21, 25176.07, 25191.69, 25190.55, 25190.95, 
    25194.43, 25185.79, 25195.85, 25197.54, 25193.13, 25219.09, 25211.59, 
    25219.26, 25214.37, 25097.9, 25103.39, 25100.42, 25106.02, 25102.07, 
    25119.71, 25125.07, 25150.47, 25139.99, 25156.72, 25141.68, 25144.34, 
    25157.27, 25142.49, 25175.13, 25152.88, 25194.57, 25171.96, 25195.99, 
    25191.62, 25198.86, 25205.4, 25213.69, 25229.21, 25225.59, 25238.74, 
    25111.63, 25118.85, 25118.21, 25125.82, 25131.48, 25143.88, 25164, 
    25156.38, 25170.41, 25173.26, 25151.95, 25164.97, 25123.71, 25130.28, 
    25126.36, 25112.2, 25158.13, 25134.32, 25178.74, 25165.49, 25204.46, 
    25185, 25223.61, 25240.64, 25256.99, 25276.53, 25122.81, 25117.88, 
    25126.72, 25139.11, 25150.69, 25166.3, 25167.91, 25170.87, 25178.58, 
    25185.12, 25171.81, 25186.76, 25131.81, 25160.22, 25116.02, 25129.14, 
    25138.38, 25134.31, 25155.51, 25160.57, 25181.41, 25170.57, 25236.4, 
    25206.79, 25291.72, 25267.09, 25116.16, 25122.79, 25146.22, 25135.01, 
    25167.35, 25175.48, 25182.14, 25190.7, 25191.62, 25196.67, 25188.4, 
    25196.34, 25166.33, 25179.67, 25143.53, 25152.19, 25148.2, 25143.83, 
    25157.37, 25172.01, 25172.33, 25177.08, 25190.58, 25167.48, 25240.31, 
    25194.82, 25130.08, 25143.08, 25144.95, 25139.89, 25174.66, 25161.91, 
    25196.55, 25187.14, 25202.59, 25194.89, 25193.76, 25183.91, 25177.79, 
    25162.49, 25150.24, 25140.62, 25142.86, 25153.44, 25172.92, 25191.7, 
    25187.59, 25201.41, 25164.97, 25180.15, 25174.25, 25189.7, 25156.18, 
    25184.66, 25149.04, 25152.11, 25161.66, 25181.19, 25185.57, 25190.24, 
    25187.37, 25173.42, 25171.15, 25161.42, 25158.76, 25151.44, 25145.42, 
    25150.92, 25156.72, 25173.42, 25188.75, 25205.49, 25209.64, 25229.73, 
    25213.34, 25240.57, 25217.37, 25257.95, 25186.34, 25216.69, 25162.1, 
    25167.86, 25178.39, 25202.8, 25189.62, 25205.05, 25171.06, 25153.8, 
    25149.39, 25141.2, 25149.58, 25148.9, 25156.96, 25154.36, 25173.98, 
    25163.39, 25193.74, 25204.93, 25237.35, 25257.87, 25279.28, 25288.92, 
    25291.88, 25293.12 ;

 HCSOI =
  25080.9, 25097.14, 25093.96, 25107.21, 25099.84, 25108.55, 25084.17, 
    25097.79, 25089.07, 25082.35, 25133.42, 25107.81, 25160.67, 25143.88, 
    25186.67, 25158.04, 25192.5, 25185.83, 25205.96, 25200.16, 25226.37, 
    25208.65, 25240.29, 25222.1, 25224.92, 25208.07, 25112.9, 25130.19, 
    25111.89, 25114.33, 25113.23, 25099.99, 25093.38, 25079.67, 25082.14, 
    25092.22, 25115.43, 25107.5, 25127.62, 25127.16, 25150.03, 25139.67, 
    25178.83, 25167.53, 25200.4, 25192.1, 25200.01, 25197.6, 25200.04, 
    25187.89, 25193.08, 25182.38, 25141.61, 25153.41, 25118.53, 25098.11, 
    25084.76, 25075.4, 25076.71, 25079.23, 25092.28, 25104.7, 25114.26, 
    25120.7, 25127.1, 25146.7, 25157.19, 25181.13, 25176.76, 25184.18, 
    25191.28, 25203.21, 25201.24, 25206.54, 25183.98, 25198.93, 25174.28, 
    25181, 25128.85, 25109.63, 25101.58, 25094.57, 25077.73, 25089.33, 
    25084.74, 25095.69, 25102.71, 25099.23, 25120.88, 25112.41, 25157.81, 
    25138.04, 25190.46, 25177.66, 25193.51, 25185.43, 25199.29, 25186.82, 
    25208.51, 25213.31, 25210.03, 25222.69, 25186.12, 25200.01, 25099.14, 
    25099.7, 25102.35, 25090.78, 25090.08, 25079.6, 25088.92, 25092.91, 
    25103.12, 25109.21, 25115.02, 25127.93, 25142.56, 25163.29, 25178.48, 
    25188.81, 25182.47, 25188.07, 25181.81, 25178.89, 25211.51, 25193.13, 
    25220.86, 25219.3, 25206.66, 25219.47, 25100.1, 25096.84, 25085.62, 
    25094.39, 25078.46, 25087.35, 25092.5, 25112.59, 25117.05, 25121.21, 
    25129.48, 25140.2, 25159.21, 25176.07, 25191.69, 25190.55, 25190.95, 
    25194.43, 25185.79, 25195.85, 25197.54, 25193.13, 25219.09, 25211.59, 
    25219.26, 25214.37, 25097.9, 25103.39, 25100.42, 25106.02, 25102.07, 
    25119.71, 25125.07, 25150.47, 25139.99, 25156.72, 25141.68, 25144.34, 
    25157.27, 25142.49, 25175.13, 25152.88, 25194.57, 25171.96, 25195.99, 
    25191.62, 25198.86, 25205.4, 25213.69, 25229.21, 25225.59, 25238.74, 
    25111.63, 25118.85, 25118.21, 25125.82, 25131.48, 25143.88, 25164, 
    25156.38, 25170.41, 25173.26, 25151.95, 25164.97, 25123.71, 25130.28, 
    25126.36, 25112.2, 25158.13, 25134.32, 25178.74, 25165.49, 25204.46, 
    25185, 25223.61, 25240.64, 25256.99, 25276.53, 25122.81, 25117.88, 
    25126.72, 25139.11, 25150.69, 25166.3, 25167.91, 25170.87, 25178.58, 
    25185.12, 25171.81, 25186.76, 25131.81, 25160.22, 25116.02, 25129.14, 
    25138.38, 25134.31, 25155.51, 25160.57, 25181.41, 25170.57, 25236.4, 
    25206.79, 25291.72, 25267.09, 25116.16, 25122.79, 25146.22, 25135.01, 
    25167.35, 25175.48, 25182.14, 25190.7, 25191.62, 25196.67, 25188.4, 
    25196.34, 25166.33, 25179.67, 25143.53, 25152.19, 25148.2, 25143.83, 
    25157.37, 25172.01, 25172.33, 25177.08, 25190.58, 25167.48, 25240.31, 
    25194.82, 25130.08, 25143.08, 25144.95, 25139.89, 25174.66, 25161.91, 
    25196.55, 25187.14, 25202.59, 25194.89, 25193.76, 25183.91, 25177.79, 
    25162.49, 25150.24, 25140.62, 25142.86, 25153.44, 25172.92, 25191.7, 
    25187.59, 25201.41, 25164.97, 25180.15, 25174.25, 25189.7, 25156.18, 
    25184.66, 25149.04, 25152.11, 25161.66, 25181.19, 25185.57, 25190.24, 
    25187.37, 25173.42, 25171.15, 25161.42, 25158.76, 25151.44, 25145.42, 
    25150.92, 25156.72, 25173.42, 25188.75, 25205.49, 25209.64, 25229.73, 
    25213.34, 25240.57, 25217.37, 25257.95, 25186.34, 25216.69, 25162.1, 
    25167.86, 25178.39, 25202.8, 25189.62, 25205.05, 25171.06, 25153.8, 
    25149.39, 25141.2, 25149.58, 25148.9, 25156.96, 25154.36, 25173.98, 
    25163.39, 25193.74, 25204.93, 25237.35, 25257.87, 25279.28, 25288.92, 
    25291.88, 25293.12 ;

 HEAT_FROM_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HR =
  7.624269e-08, 7.645139e-08, 7.641083e-08, 7.657911e-08, 7.648578e-08, 
    7.659595e-08, 7.628502e-08, 7.645966e-08, 7.634819e-08, 7.62615e-08, 
    7.690554e-08, 7.658662e-08, 7.723681e-08, 7.70335e-08, 7.754418e-08, 
    7.720516e-08, 7.761253e-08, 7.753444e-08, 7.776953e-08, 7.77022e-08, 
    7.800275e-08, 7.780061e-08, 7.815856e-08, 7.79545e-08, 7.798641e-08, 
    7.779394e-08, 7.665084e-08, 7.686582e-08, 7.663809e-08, 7.666875e-08, 
    7.6655e-08, 7.648769e-08, 7.640334e-08, 7.622676e-08, 7.625883e-08, 
    7.638853e-08, 7.668255e-08, 7.658277e-08, 7.683426e-08, 7.682858e-08, 
    7.710845e-08, 7.698227e-08, 7.745253e-08, 7.731892e-08, 7.7705e-08, 
    7.760792e-08, 7.770044e-08, 7.767239e-08, 7.77008e-08, 7.755842e-08, 
    7.761943e-08, 7.749413e-08, 7.700589e-08, 7.71494e-08, 7.67213e-08, 
    7.646373e-08, 7.629267e-08, 7.617125e-08, 7.618841e-08, 7.622113e-08, 
    7.638929e-08, 7.654739e-08, 7.666784e-08, 7.674839e-08, 7.682777e-08, 
    7.706788e-08, 7.719501e-08, 7.747953e-08, 7.742823e-08, 7.751517e-08, 
    7.759827e-08, 7.773771e-08, 7.771477e-08, 7.777619e-08, 7.75129e-08, 
    7.768788e-08, 7.739899e-08, 7.747801e-08, 7.684923e-08, 7.66097e-08, 
    7.650777e-08, 7.641862e-08, 7.620162e-08, 7.635147e-08, 7.629239e-08, 
    7.643295e-08, 7.652225e-08, 7.647809e-08, 7.67506e-08, 7.664466e-08, 
    7.720254e-08, 7.696229e-08, 7.758857e-08, 7.743876e-08, 7.762448e-08, 
    7.752973e-08, 7.769207e-08, 7.754596e-08, 7.779906e-08, 7.785415e-08, 
    7.78165e-08, 7.796114e-08, 7.753786e-08, 7.770043e-08, 7.647685e-08, 
    7.648405e-08, 7.651761e-08, 7.637008e-08, 7.636106e-08, 7.622587e-08, 
    7.634618e-08, 7.639739e-08, 7.652743e-08, 7.660432e-08, 7.667741e-08, 
    7.683809e-08, 7.701749e-08, 7.72683e-08, 7.744847e-08, 7.75692e-08, 
    7.749518e-08, 7.756054e-08, 7.748747e-08, 7.745323e-08, 7.78335e-08, 
    7.761999e-08, 7.794034e-08, 7.792262e-08, 7.777765e-08, 7.792462e-08, 
    7.648911e-08, 7.644767e-08, 7.630373e-08, 7.641638e-08, 7.621115e-08, 
    7.632602e-08, 7.639206e-08, 7.664685e-08, 7.670285e-08, 7.675474e-08, 
    7.685723e-08, 7.698873e-08, 7.721936e-08, 7.741998e-08, 7.76031e-08, 
    7.758969e-08, 7.759441e-08, 7.76353e-08, 7.7534e-08, 7.765193e-08, 
    7.767171e-08, 7.761997e-08, 7.792025e-08, 7.783448e-08, 7.792224e-08, 
    7.78664e-08, 7.646114e-08, 7.653087e-08, 7.649319e-08, 7.656404e-08, 
    7.651412e-08, 7.673605e-08, 7.680259e-08, 7.711383e-08, 7.698614e-08, 
    7.718939e-08, 7.70068e-08, 7.703915e-08, 7.719597e-08, 7.701667e-08, 
    7.74089e-08, 7.714296e-08, 7.763688e-08, 7.737135e-08, 7.765352e-08, 
    7.760231e-08, 7.768711e-08, 7.776304e-08, 7.785858e-08, 7.803479e-08, 
    7.7994e-08, 7.814135e-08, 7.663483e-08, 7.672524e-08, 7.671731e-08, 
    7.681193e-08, 7.68819e-08, 7.703356e-08, 7.727672e-08, 7.71853e-08, 
    7.735314e-08, 7.738683e-08, 7.713184e-08, 7.728839e-08, 7.678577e-08, 
    7.686698e-08, 7.681864e-08, 7.664195e-08, 7.720634e-08, 7.691673e-08, 
    7.745144e-08, 7.729462e-08, 7.775221e-08, 7.752466e-08, 7.797154e-08, 
    7.816244e-08, 7.834216e-08, 7.855203e-08, 7.677461e-08, 7.671318e-08, 
    7.682319e-08, 7.697533e-08, 7.711654e-08, 7.730418e-08, 7.732339e-08, 
    7.735854e-08, 7.744958e-08, 7.752611e-08, 7.736963e-08, 7.754529e-08, 
    7.688577e-08, 7.723148e-08, 7.668994e-08, 7.685301e-08, 7.696638e-08, 
    7.691667e-08, 7.717485e-08, 7.723568e-08, 7.748282e-08, 7.735509e-08, 
    7.811531e-08, 7.777906e-08, 7.871185e-08, 7.845127e-08, 7.669171e-08, 
    7.677441e-08, 7.706215e-08, 7.692525e-08, 7.731672e-08, 7.741303e-08, 
    7.749135e-08, 7.75914e-08, 7.760222e-08, 7.76615e-08, 7.756436e-08, 
    7.765767e-08, 7.730458e-08, 7.74624e-08, 7.702928e-08, 7.713471e-08, 
    7.708622e-08, 7.703301e-08, 7.719722e-08, 7.737208e-08, 7.737585e-08, 
    7.743191e-08, 7.758979e-08, 7.731831e-08, 7.815863e-08, 7.763973e-08, 
    7.686458e-08, 7.702379e-08, 7.704657e-08, 7.698489e-08, 7.740338e-08, 
    7.725177e-08, 7.766006e-08, 7.754974e-08, 7.77305e-08, 7.764068e-08, 
    7.762746e-08, 7.75121e-08, 7.744025e-08, 7.725872e-08, 7.711099e-08, 
    7.699384e-08, 7.702109e-08, 7.714976e-08, 7.738279e-08, 7.760318e-08, 
    7.755491e-08, 7.771676e-08, 7.728835e-08, 7.7468e-08, 7.739856e-08, 
    7.757962e-08, 7.718286e-08, 7.752063e-08, 7.709649e-08, 7.713369e-08, 
    7.724876e-08, 7.748016e-08, 7.75314e-08, 7.758604e-08, 7.755232e-08, 
    7.738871e-08, 7.736191e-08, 7.724597e-08, 7.721394e-08, 7.71256e-08, 
    7.705243e-08, 7.711927e-08, 7.718945e-08, 7.738879e-08, 7.756837e-08, 
    7.776411e-08, 7.781203e-08, 7.804059e-08, 7.785449e-08, 7.816151e-08, 
    7.790043e-08, 7.835236e-08, 7.754026e-08, 7.789281e-08, 7.725401e-08, 
    7.732286e-08, 7.744735e-08, 7.773286e-08, 7.757877e-08, 7.775899e-08, 
    7.736087e-08, 7.715419e-08, 7.710074e-08, 7.700096e-08, 7.710302e-08, 
    7.709473e-08, 7.719238e-08, 7.7161e-08, 7.739541e-08, 7.72695e-08, 
    7.762712e-08, 7.775758e-08, 7.812591e-08, 7.835159e-08, 7.858132e-08, 
    7.86827e-08, 7.871355e-08, 7.872645e-08 ;

 HR_vr =
  2.780871e-07, 2.787966e-07, 2.786588e-07, 2.792304e-07, 2.789135e-07, 
    2.792876e-07, 2.782311e-07, 2.788246e-07, 2.784459e-07, 2.781512e-07, 
    2.803378e-07, 2.792559e-07, 2.814609e-07, 2.807722e-07, 2.825011e-07, 
    2.813536e-07, 2.827323e-07, 2.824684e-07, 2.832631e-07, 2.830356e-07, 
    2.840504e-07, 2.833681e-07, 2.845762e-07, 2.838877e-07, 2.839953e-07, 
    2.833456e-07, 2.794741e-07, 2.802031e-07, 2.794308e-07, 2.795348e-07, 
    2.794882e-07, 2.789199e-07, 2.786332e-07, 2.780331e-07, 2.781421e-07, 
    2.785829e-07, 2.795816e-07, 2.79243e-07, 2.800966e-07, 2.800774e-07, 
    2.810262e-07, 2.805985e-07, 2.821913e-07, 2.817391e-07, 2.830451e-07, 
    2.827169e-07, 2.830296e-07, 2.829348e-07, 2.830309e-07, 2.825495e-07, 
    2.827557e-07, 2.82332e-07, 2.806786e-07, 2.811649e-07, 2.797132e-07, 
    2.788382e-07, 2.782571e-07, 2.778442e-07, 2.779026e-07, 2.780139e-07, 
    2.785855e-07, 2.791228e-07, 2.795318e-07, 2.798052e-07, 2.800746e-07, 
    2.808884e-07, 2.813193e-07, 2.822825e-07, 2.821091e-07, 2.824031e-07, 
    2.826842e-07, 2.831556e-07, 2.83078e-07, 2.832855e-07, 2.823955e-07, 
    2.829871e-07, 2.820102e-07, 2.822775e-07, 2.801468e-07, 2.793344e-07, 
    2.789879e-07, 2.786852e-07, 2.779475e-07, 2.78457e-07, 2.782562e-07, 
    2.78734e-07, 2.790374e-07, 2.788874e-07, 2.798127e-07, 2.794531e-07, 
    2.813448e-07, 2.805307e-07, 2.826514e-07, 2.821447e-07, 2.827729e-07, 
    2.824524e-07, 2.830013e-07, 2.825074e-07, 2.833629e-07, 2.835488e-07, 
    2.834217e-07, 2.839102e-07, 2.8248e-07, 2.830295e-07, 2.788832e-07, 
    2.789076e-07, 2.790216e-07, 2.785202e-07, 2.784896e-07, 2.7803e-07, 
    2.78439e-07, 2.786131e-07, 2.79055e-07, 2.793161e-07, 2.795643e-07, 
    2.801095e-07, 2.807178e-07, 2.815676e-07, 2.821776e-07, 2.82586e-07, 
    2.823356e-07, 2.825567e-07, 2.823095e-07, 2.821937e-07, 2.834791e-07, 
    2.827576e-07, 2.8384e-07, 2.837802e-07, 2.832905e-07, 2.837869e-07, 
    2.789248e-07, 2.78784e-07, 2.782947e-07, 2.786777e-07, 2.7798e-07, 
    2.783705e-07, 2.785949e-07, 2.794604e-07, 2.796507e-07, 2.798267e-07, 
    2.801745e-07, 2.806204e-07, 2.814019e-07, 2.820811e-07, 2.827006e-07, 
    2.826553e-07, 2.826712e-07, 2.828094e-07, 2.824669e-07, 2.828657e-07, 
    2.829325e-07, 2.827576e-07, 2.837722e-07, 2.834825e-07, 2.837789e-07, 
    2.835904e-07, 2.788298e-07, 2.790667e-07, 2.789387e-07, 2.791793e-07, 
    2.790097e-07, 2.797632e-07, 2.799889e-07, 2.810443e-07, 2.806116e-07, 
    2.813003e-07, 2.806817e-07, 2.807913e-07, 2.813224e-07, 2.807152e-07, 
    2.820435e-07, 2.811429e-07, 2.828148e-07, 2.819162e-07, 2.82871e-07, 
    2.826979e-07, 2.829846e-07, 2.832411e-07, 2.835639e-07, 2.841587e-07, 
    2.84021e-07, 2.845183e-07, 2.794197e-07, 2.797266e-07, 2.796997e-07, 
    2.800208e-07, 2.802581e-07, 2.807724e-07, 2.815962e-07, 2.812866e-07, 
    2.81855e-07, 2.81969e-07, 2.811055e-07, 2.816356e-07, 2.79932e-07, 
    2.802074e-07, 2.800435e-07, 2.794438e-07, 2.813577e-07, 2.803761e-07, 
    2.821876e-07, 2.816568e-07, 2.832046e-07, 2.824352e-07, 2.839452e-07, 
    2.845891e-07, 2.851953e-07, 2.859018e-07, 2.798942e-07, 2.796857e-07, 
    2.800591e-07, 2.805749e-07, 2.810536e-07, 2.816892e-07, 2.817543e-07, 
    2.818732e-07, 2.821813e-07, 2.824402e-07, 2.819106e-07, 2.825051e-07, 
    2.802708e-07, 2.814429e-07, 2.796068e-07, 2.8016e-07, 2.805446e-07, 
    2.803761e-07, 2.812513e-07, 2.814573e-07, 2.822937e-07, 2.818616e-07, 
    2.844301e-07, 2.832951e-07, 2.864398e-07, 2.855626e-07, 2.796128e-07, 
    2.798935e-07, 2.808692e-07, 2.804052e-07, 2.817317e-07, 2.820576e-07, 
    2.823227e-07, 2.82661e-07, 2.826976e-07, 2.82898e-07, 2.825696e-07, 
    2.828851e-07, 2.816905e-07, 2.822247e-07, 2.80758e-07, 2.811152e-07, 
    2.80951e-07, 2.807706e-07, 2.81327e-07, 2.819189e-07, 2.819318e-07, 
    2.821214e-07, 2.826549e-07, 2.81737e-07, 2.845759e-07, 2.828238e-07, 
    2.801995e-07, 2.807391e-07, 2.808165e-07, 2.806075e-07, 2.82025e-07, 
    2.815117e-07, 2.828932e-07, 2.825202e-07, 2.831312e-07, 2.828276e-07, 
    2.827829e-07, 2.823928e-07, 2.821497e-07, 2.815352e-07, 2.810348e-07, 
    2.806378e-07, 2.807302e-07, 2.811662e-07, 2.819552e-07, 2.827008e-07, 
    2.825375e-07, 2.830848e-07, 2.816356e-07, 2.822435e-07, 2.820086e-07, 
    2.826212e-07, 2.812783e-07, 2.824211e-07, 2.809857e-07, 2.811118e-07, 
    2.815015e-07, 2.822846e-07, 2.824581e-07, 2.826428e-07, 2.825289e-07, 
    2.819752e-07, 2.818846e-07, 2.814921e-07, 2.813836e-07, 2.810844e-07, 
    2.808364e-07, 2.810629e-07, 2.813006e-07, 2.819756e-07, 2.82583e-07, 
    2.832448e-07, 2.834067e-07, 2.841779e-07, 2.835498e-07, 2.845855e-07, 
    2.837045e-07, 2.852291e-07, 2.824877e-07, 2.836791e-07, 2.815193e-07, 
    2.817525e-07, 2.821736e-07, 2.831389e-07, 2.826183e-07, 2.832273e-07, 
    2.818811e-07, 2.81181e-07, 2.810002e-07, 2.806619e-07, 2.810079e-07, 
    2.809798e-07, 2.813106e-07, 2.812043e-07, 2.81998e-07, 2.815718e-07, 
    2.827817e-07, 2.832226e-07, 2.844661e-07, 2.852268e-07, 2.860007e-07, 
    2.863418e-07, 2.864456e-07, 2.86489e-07,
  2.756907e-07, 2.764159e-07, 2.762751e-07, 2.768594e-07, 2.765354e-07, 
    2.769179e-07, 2.758379e-07, 2.764446e-07, 2.760574e-07, 2.757562e-07, 
    2.779915e-07, 2.768855e-07, 2.791394e-07, 2.784354e-07, 2.802028e-07, 
    2.790298e-07, 2.804391e-07, 2.801693e-07, 2.809817e-07, 2.807491e-07, 
    2.817864e-07, 2.81089e-07, 2.823239e-07, 2.816201e-07, 2.817302e-07, 
    2.81066e-07, 2.771085e-07, 2.778538e-07, 2.770642e-07, 2.771706e-07, 
    2.771229e-07, 2.76542e-07, 2.762489e-07, 2.756354e-07, 2.757469e-07, 
    2.761976e-07, 2.772184e-07, 2.768722e-07, 2.777448e-07, 2.777252e-07, 
    2.786951e-07, 2.782579e-07, 2.798861e-07, 2.794238e-07, 2.807588e-07, 
    2.804233e-07, 2.80743e-07, 2.806461e-07, 2.807442e-07, 2.802522e-07, 
    2.80463e-07, 2.800299e-07, 2.783398e-07, 2.788369e-07, 2.773529e-07, 
    2.764586e-07, 2.758645e-07, 2.754424e-07, 2.755021e-07, 2.756158e-07, 
    2.762002e-07, 2.767494e-07, 2.771675e-07, 2.77447e-07, 2.777223e-07, 
    2.785543e-07, 2.789947e-07, 2.799793e-07, 2.79802e-07, 2.801026e-07, 
    2.803899e-07, 2.808717e-07, 2.807925e-07, 2.810046e-07, 2.800948e-07, 
    2.806995e-07, 2.797009e-07, 2.799742e-07, 2.777963e-07, 2.769657e-07, 
    2.766116e-07, 2.763021e-07, 2.755479e-07, 2.760688e-07, 2.758635e-07, 
    2.76352e-07, 2.766621e-07, 2.765088e-07, 2.774547e-07, 2.770871e-07, 
    2.790208e-07, 2.781886e-07, 2.803564e-07, 2.798384e-07, 2.804805e-07, 
    2.80153e-07, 2.80714e-07, 2.802092e-07, 2.810836e-07, 2.812738e-07, 
    2.811438e-07, 2.816431e-07, 2.801811e-07, 2.807429e-07, 2.765044e-07, 
    2.765294e-07, 2.76646e-07, 2.761334e-07, 2.761021e-07, 2.756323e-07, 
    2.760505e-07, 2.762283e-07, 2.766801e-07, 2.76947e-07, 2.772007e-07, 
    2.777581e-07, 2.783799e-07, 2.792486e-07, 2.79872e-07, 2.802895e-07, 
    2.800336e-07, 2.802595e-07, 2.800069e-07, 2.798885e-07, 2.812025e-07, 
    2.804649e-07, 2.815713e-07, 2.815102e-07, 2.810096e-07, 2.815171e-07, 
    2.76547e-07, 2.764031e-07, 2.759029e-07, 2.762944e-07, 2.755811e-07, 
    2.759804e-07, 2.762098e-07, 2.770946e-07, 2.77289e-07, 2.77469e-07, 
    2.778245e-07, 2.782803e-07, 2.790791e-07, 2.797734e-07, 2.804067e-07, 
    2.803603e-07, 2.803766e-07, 2.805179e-07, 2.801678e-07, 2.805754e-07, 
    2.806437e-07, 2.80465e-07, 2.81502e-07, 2.812059e-07, 2.815089e-07, 
    2.813162e-07, 2.764499e-07, 2.76692e-07, 2.765612e-07, 2.768072e-07, 
    2.766338e-07, 2.77404e-07, 2.776348e-07, 2.787136e-07, 2.782713e-07, 
    2.789753e-07, 2.783429e-07, 2.78455e-07, 2.789979e-07, 2.783772e-07, 
    2.79735e-07, 2.788144e-07, 2.805234e-07, 2.79605e-07, 2.805809e-07, 
    2.804039e-07, 2.80697e-07, 2.809592e-07, 2.812891e-07, 2.818971e-07, 
    2.817565e-07, 2.822647e-07, 2.770529e-07, 2.773666e-07, 2.773392e-07, 
    2.776674e-07, 2.7791e-07, 2.784357e-07, 2.792777e-07, 2.789613e-07, 
    2.795423e-07, 2.796588e-07, 2.787762e-07, 2.793181e-07, 2.775766e-07, 
    2.778581e-07, 2.776906e-07, 2.770776e-07, 2.79034e-07, 2.780306e-07, 
    2.798823e-07, 2.793397e-07, 2.809218e-07, 2.801354e-07, 2.81679e-07, 
    2.823371e-07, 2.829567e-07, 2.83679e-07, 2.775379e-07, 2.773248e-07, 
    2.777065e-07, 2.782338e-07, 2.787231e-07, 2.793728e-07, 2.794393e-07, 
    2.795609e-07, 2.798759e-07, 2.801405e-07, 2.795992e-07, 2.802068e-07, 
    2.77923e-07, 2.791211e-07, 2.772441e-07, 2.778097e-07, 2.782028e-07, 
    2.780305e-07, 2.789251e-07, 2.791357e-07, 2.799907e-07, 2.79549e-07, 
    2.821746e-07, 2.810144e-07, 2.842289e-07, 2.833323e-07, 2.772503e-07, 
    2.775373e-07, 2.785346e-07, 2.780603e-07, 2.794162e-07, 2.797494e-07, 
    2.800203e-07, 2.803662e-07, 2.804036e-07, 2.806084e-07, 2.802728e-07, 
    2.805953e-07, 2.793742e-07, 2.799202e-07, 2.784209e-07, 2.787861e-07, 
    2.786182e-07, 2.784338e-07, 2.790026e-07, 2.796076e-07, 2.796208e-07, 
    2.798147e-07, 2.803601e-07, 2.794217e-07, 2.823237e-07, 2.805327e-07, 
    2.7785e-07, 2.784017e-07, 2.784807e-07, 2.78267e-07, 2.79716e-07, 
    2.791914e-07, 2.806035e-07, 2.802222e-07, 2.808468e-07, 2.805365e-07, 
    2.804908e-07, 2.800921e-07, 2.798436e-07, 2.792154e-07, 2.787039e-07, 
    2.782981e-07, 2.783925e-07, 2.788382e-07, 2.796447e-07, 2.804069e-07, 
    2.8024e-07, 2.807994e-07, 2.79318e-07, 2.799395e-07, 2.796993e-07, 
    2.803255e-07, 2.789528e-07, 2.801211e-07, 2.786537e-07, 2.787826e-07, 
    2.79181e-07, 2.799814e-07, 2.801588e-07, 2.803476e-07, 2.802311e-07, 
    2.796652e-07, 2.795726e-07, 2.791714e-07, 2.790604e-07, 2.787546e-07, 
    2.785011e-07, 2.787326e-07, 2.789756e-07, 2.796656e-07, 2.802865e-07, 
    2.809629e-07, 2.811285e-07, 2.819169e-07, 2.812748e-07, 2.823336e-07, 
    2.81433e-07, 2.829914e-07, 2.801891e-07, 2.81407e-07, 2.791992e-07, 
    2.794375e-07, 2.79868e-07, 2.808548e-07, 2.803226e-07, 2.809451e-07, 
    2.79569e-07, 2.788534e-07, 2.786685e-07, 2.783227e-07, 2.786764e-07, 
    2.786476e-07, 2.789858e-07, 2.788772e-07, 2.796885e-07, 2.792528e-07, 
    2.804896e-07, 2.809402e-07, 2.822113e-07, 2.82989e-07, 2.8378e-07, 
    2.841288e-07, 2.842349e-07, 2.842792e-07,
  2.758359e-07, 2.765716e-07, 2.764287e-07, 2.770216e-07, 2.766928e-07, 
    2.770809e-07, 2.759852e-07, 2.766007e-07, 2.762079e-07, 2.759023e-07, 
    2.781708e-07, 2.770481e-07, 2.793362e-07, 2.786213e-07, 2.804162e-07, 
    2.792248e-07, 2.806563e-07, 2.803821e-07, 2.812075e-07, 2.809712e-07, 
    2.820255e-07, 2.813166e-07, 2.825719e-07, 2.818564e-07, 2.819683e-07, 
    2.812932e-07, 2.772744e-07, 2.78031e-07, 2.772294e-07, 2.773374e-07, 
    2.77289e-07, 2.766996e-07, 2.764022e-07, 2.757798e-07, 2.758929e-07, 
    2.763501e-07, 2.77386e-07, 2.770346e-07, 2.779202e-07, 2.779002e-07, 
    2.788849e-07, 2.784411e-07, 2.800944e-07, 2.796249e-07, 2.80981e-07, 
    2.806402e-07, 2.80965e-07, 2.808665e-07, 2.809663e-07, 2.804663e-07, 
    2.806806e-07, 2.802405e-07, 2.785241e-07, 2.790289e-07, 2.775224e-07, 
    2.76615e-07, 2.760122e-07, 2.75584e-07, 2.756446e-07, 2.757599e-07, 
    2.763528e-07, 2.769099e-07, 2.773342e-07, 2.776179e-07, 2.778974e-07, 
    2.78742e-07, 2.791892e-07, 2.801892e-07, 2.80009e-07, 2.803144e-07, 
    2.806063e-07, 2.810958e-07, 2.810153e-07, 2.812309e-07, 2.803065e-07, 
    2.809209e-07, 2.799063e-07, 2.801839e-07, 2.779726e-07, 2.771295e-07, 
    2.767702e-07, 2.764561e-07, 2.756911e-07, 2.762195e-07, 2.760112e-07, 
    2.765067e-07, 2.768214e-07, 2.766658e-07, 2.776257e-07, 2.772526e-07, 
    2.792157e-07, 2.783707e-07, 2.805722e-07, 2.80046e-07, 2.806983e-07, 
    2.803656e-07, 2.809356e-07, 2.804226e-07, 2.813111e-07, 2.815044e-07, 
    2.813723e-07, 2.818797e-07, 2.803941e-07, 2.809649e-07, 2.766614e-07, 
    2.766868e-07, 2.76805e-07, 2.76285e-07, 2.762533e-07, 2.757767e-07, 
    2.762008e-07, 2.763813e-07, 2.768396e-07, 2.771105e-07, 2.773679e-07, 
    2.779337e-07, 2.785649e-07, 2.794469e-07, 2.800801e-07, 2.805042e-07, 
    2.802443e-07, 2.804738e-07, 2.802172e-07, 2.800969e-07, 2.814319e-07, 
    2.806825e-07, 2.818068e-07, 2.817447e-07, 2.812359e-07, 2.817517e-07, 
    2.767046e-07, 2.765586e-07, 2.760512e-07, 2.764483e-07, 2.757247e-07, 
    2.761298e-07, 2.763625e-07, 2.772602e-07, 2.774575e-07, 2.776402e-07, 
    2.78001e-07, 2.784638e-07, 2.792749e-07, 2.7998e-07, 2.806233e-07, 
    2.805762e-07, 2.805928e-07, 2.807363e-07, 2.803806e-07, 2.807947e-07, 
    2.808641e-07, 2.806825e-07, 2.817363e-07, 2.814354e-07, 2.817433e-07, 
    2.815474e-07, 2.766061e-07, 2.768518e-07, 2.76719e-07, 2.769686e-07, 
    2.767927e-07, 2.775743e-07, 2.778086e-07, 2.789037e-07, 2.784546e-07, 
    2.791695e-07, 2.785273e-07, 2.786411e-07, 2.791925e-07, 2.785621e-07, 
    2.79941e-07, 2.790062e-07, 2.807419e-07, 2.79809e-07, 2.808003e-07, 
    2.806205e-07, 2.809182e-07, 2.811847e-07, 2.8152e-07, 2.82138e-07, 
    2.81995e-07, 2.825116e-07, 2.77218e-07, 2.775363e-07, 2.775084e-07, 
    2.778416e-07, 2.780878e-07, 2.786215e-07, 2.794765e-07, 2.791552e-07, 
    2.797452e-07, 2.798635e-07, 2.789672e-07, 2.795175e-07, 2.777495e-07, 
    2.780352e-07, 2.778652e-07, 2.77243e-07, 2.792291e-07, 2.782103e-07, 
    2.800905e-07, 2.795395e-07, 2.811467e-07, 2.803477e-07, 2.819162e-07, 
    2.825854e-07, 2.832153e-07, 2.8395e-07, 2.777102e-07, 2.774939e-07, 
    2.778812e-07, 2.784166e-07, 2.789133e-07, 2.795731e-07, 2.796406e-07, 
    2.797641e-07, 2.80084e-07, 2.803529e-07, 2.79803e-07, 2.804203e-07, 
    2.781012e-07, 2.793175e-07, 2.77412e-07, 2.779861e-07, 2.783851e-07, 
    2.782102e-07, 2.791185e-07, 2.793323e-07, 2.802007e-07, 2.79752e-07, 
    2.824201e-07, 2.812408e-07, 2.845094e-07, 2.835973e-07, 2.774183e-07, 
    2.777095e-07, 2.78722e-07, 2.782404e-07, 2.796172e-07, 2.799556e-07, 
    2.802308e-07, 2.805822e-07, 2.806202e-07, 2.808283e-07, 2.804872e-07, 
    2.808149e-07, 2.795745e-07, 2.801291e-07, 2.786065e-07, 2.789773e-07, 
    2.788068e-07, 2.786196e-07, 2.791971e-07, 2.798116e-07, 2.79825e-07, 
    2.800219e-07, 2.805762e-07, 2.796228e-07, 2.825718e-07, 2.807515e-07, 
    2.780269e-07, 2.78587e-07, 2.786672e-07, 2.784503e-07, 2.799217e-07, 
    2.793888e-07, 2.808232e-07, 2.804359e-07, 2.810705e-07, 2.807552e-07, 
    2.807088e-07, 2.803037e-07, 2.800512e-07, 2.794133e-07, 2.788938e-07, 
    2.784818e-07, 2.785777e-07, 2.790302e-07, 2.798493e-07, 2.806235e-07, 
    2.804539e-07, 2.810223e-07, 2.795175e-07, 2.801487e-07, 2.799047e-07, 
    2.805408e-07, 2.791466e-07, 2.803333e-07, 2.788429e-07, 2.789737e-07, 
    2.793783e-07, 2.801913e-07, 2.803714e-07, 2.805633e-07, 2.80445e-07, 
    2.798701e-07, 2.79776e-07, 2.793685e-07, 2.792559e-07, 2.789452e-07, 
    2.786879e-07, 2.78923e-07, 2.791697e-07, 2.798704e-07, 2.805012e-07, 
    2.811885e-07, 2.813567e-07, 2.821581e-07, 2.815055e-07, 2.825819e-07, 
    2.816664e-07, 2.832507e-07, 2.804024e-07, 2.816399e-07, 2.793967e-07, 
    2.796388e-07, 2.800761e-07, 2.810787e-07, 2.805378e-07, 2.811704e-07, 
    2.797723e-07, 2.790457e-07, 2.788578e-07, 2.785068e-07, 2.788659e-07, 
    2.788367e-07, 2.791801e-07, 2.790698e-07, 2.798937e-07, 2.794512e-07, 
    2.807076e-07, 2.811655e-07, 2.824574e-07, 2.832482e-07, 2.840526e-07, 
    2.844074e-07, 2.845154e-07, 2.845605e-07,
  2.694351e-07, 2.701692e-07, 2.700265e-07, 2.706184e-07, 2.702901e-07, 
    2.706776e-07, 2.69584e-07, 2.701983e-07, 2.698062e-07, 2.695012e-07, 
    2.717662e-07, 2.706448e-07, 2.729308e-07, 2.722161e-07, 2.74011e-07, 
    2.728196e-07, 2.742512e-07, 2.739768e-07, 2.748028e-07, 2.745662e-07, 
    2.756221e-07, 2.749121e-07, 2.761693e-07, 2.754526e-07, 2.755647e-07, 
    2.748886e-07, 2.708707e-07, 2.716266e-07, 2.708258e-07, 2.709336e-07, 
    2.708853e-07, 2.702969e-07, 2.700002e-07, 2.69379e-07, 2.694918e-07, 
    2.699481e-07, 2.709821e-07, 2.706313e-07, 2.715156e-07, 2.714957e-07, 
    2.724796e-07, 2.72036e-07, 2.73689e-07, 2.732194e-07, 2.745761e-07, 
    2.74235e-07, 2.745601e-07, 2.744615e-07, 2.745614e-07, 2.740611e-07, 
    2.742754e-07, 2.738352e-07, 2.721191e-07, 2.726236e-07, 2.711184e-07, 
    2.702126e-07, 2.696109e-07, 2.691837e-07, 2.692441e-07, 2.693592e-07, 
    2.699508e-07, 2.705068e-07, 2.709304e-07, 2.712137e-07, 2.714928e-07, 
    2.72337e-07, 2.727839e-07, 2.737839e-07, 2.736035e-07, 2.739091e-07, 
    2.742011e-07, 2.74691e-07, 2.746104e-07, 2.748262e-07, 2.739011e-07, 
    2.745159e-07, 2.735008e-07, 2.737785e-07, 2.715682e-07, 2.70726e-07, 
    2.703675e-07, 2.700539e-07, 2.692906e-07, 2.698177e-07, 2.6961e-07, 
    2.701044e-07, 2.704184e-07, 2.702631e-07, 2.712214e-07, 2.708489e-07, 
    2.728103e-07, 2.719658e-07, 2.74167e-07, 2.736406e-07, 2.742932e-07, 
    2.739602e-07, 2.745307e-07, 2.740173e-07, 2.749066e-07, 2.751001e-07, 
    2.749678e-07, 2.754759e-07, 2.739888e-07, 2.7456e-07, 2.702587e-07, 
    2.702841e-07, 2.704021e-07, 2.698832e-07, 2.698515e-07, 2.693759e-07, 
    2.697991e-07, 2.699792e-07, 2.704366e-07, 2.70707e-07, 2.709641e-07, 
    2.715291e-07, 2.721598e-07, 2.730415e-07, 2.736747e-07, 2.74099e-07, 
    2.738389e-07, 2.740685e-07, 2.738118e-07, 2.736914e-07, 2.750275e-07, 
    2.742774e-07, 2.754029e-07, 2.753407e-07, 2.748313e-07, 2.753476e-07, 
    2.703019e-07, 2.701561e-07, 2.696498e-07, 2.70046e-07, 2.693241e-07, 
    2.697282e-07, 2.699605e-07, 2.708566e-07, 2.710536e-07, 2.71236e-07, 
    2.715964e-07, 2.720587e-07, 2.728695e-07, 2.735746e-07, 2.742181e-07, 
    2.741709e-07, 2.741875e-07, 2.743312e-07, 2.739752e-07, 2.743896e-07, 
    2.744592e-07, 2.742774e-07, 2.753323e-07, 2.75031e-07, 2.753393e-07, 
    2.751432e-07, 2.702035e-07, 2.704487e-07, 2.703162e-07, 2.705654e-07, 
    2.703898e-07, 2.711703e-07, 2.714042e-07, 2.724985e-07, 2.720496e-07, 
    2.727641e-07, 2.721222e-07, 2.72236e-07, 2.727872e-07, 2.72157e-07, 
    2.735356e-07, 2.726009e-07, 2.743368e-07, 2.734037e-07, 2.743952e-07, 
    2.742153e-07, 2.745133e-07, 2.7478e-07, 2.751157e-07, 2.757346e-07, 
    2.755914e-07, 2.761089e-07, 2.708144e-07, 2.711323e-07, 2.711044e-07, 
    2.714371e-07, 2.716831e-07, 2.722163e-07, 2.730711e-07, 2.727497e-07, 
    2.733397e-07, 2.734581e-07, 2.725618e-07, 2.731121e-07, 2.713451e-07, 
    2.716307e-07, 2.714607e-07, 2.708394e-07, 2.728237e-07, 2.718056e-07, 
    2.736851e-07, 2.73134e-07, 2.74742e-07, 2.739424e-07, 2.755125e-07, 
    2.76183e-07, 2.768141e-07, 2.775509e-07, 2.713059e-07, 2.710899e-07, 
    2.714767e-07, 2.720116e-07, 2.72508e-07, 2.731676e-07, 2.732351e-07, 
    2.733586e-07, 2.736786e-07, 2.739475e-07, 2.733976e-07, 2.740149e-07, 
    2.716967e-07, 2.72912e-07, 2.710081e-07, 2.715815e-07, 2.719801e-07, 
    2.718054e-07, 2.72713e-07, 2.729268e-07, 2.737954e-07, 2.733465e-07, 
    2.760174e-07, 2.748363e-07, 2.78112e-07, 2.771972e-07, 2.710144e-07, 
    2.713052e-07, 2.723168e-07, 2.718356e-07, 2.732117e-07, 2.735502e-07, 
    2.738254e-07, 2.74177e-07, 2.74215e-07, 2.744233e-07, 2.740819e-07, 
    2.744098e-07, 2.73169e-07, 2.737236e-07, 2.722013e-07, 2.725719e-07, 
    2.724015e-07, 2.722144e-07, 2.727916e-07, 2.734062e-07, 2.734195e-07, 
    2.736165e-07, 2.741713e-07, 2.732173e-07, 2.761696e-07, 2.743467e-07, 
    2.716222e-07, 2.72182e-07, 2.72262e-07, 2.720452e-07, 2.735162e-07, 
    2.729834e-07, 2.744182e-07, 2.740306e-07, 2.746657e-07, 2.743501e-07, 
    2.743037e-07, 2.738983e-07, 2.736458e-07, 2.730078e-07, 2.724885e-07, 
    2.720767e-07, 2.721725e-07, 2.726248e-07, 2.734439e-07, 2.742184e-07, 
    2.740487e-07, 2.746174e-07, 2.731119e-07, 2.737433e-07, 2.734993e-07, 
    2.741355e-07, 2.727412e-07, 2.739283e-07, 2.724375e-07, 2.725683e-07, 
    2.729728e-07, 2.73786e-07, 2.739661e-07, 2.741581e-07, 2.740396e-07, 
    2.734647e-07, 2.733705e-07, 2.72963e-07, 2.728504e-07, 2.725399e-07, 
    2.722826e-07, 2.725176e-07, 2.727643e-07, 2.734649e-07, 2.74096e-07, 
    2.747838e-07, 2.749522e-07, 2.75755e-07, 2.751013e-07, 2.761797e-07, 
    2.752627e-07, 2.768499e-07, 2.739972e-07, 2.752359e-07, 2.729913e-07, 
    2.732332e-07, 2.736708e-07, 2.74674e-07, 2.741326e-07, 2.747658e-07, 
    2.733668e-07, 2.726404e-07, 2.724525e-07, 2.721017e-07, 2.724605e-07, 
    2.724314e-07, 2.727746e-07, 2.726643e-07, 2.734882e-07, 2.730457e-07, 
    2.743025e-07, 2.747608e-07, 2.760547e-07, 2.768472e-07, 2.776538e-07, 
    2.780097e-07, 2.78118e-07, 2.781633e-07,
  2.510366e-07, 2.517468e-07, 2.516088e-07, 2.521818e-07, 2.518639e-07, 
    2.522391e-07, 2.511806e-07, 2.51775e-07, 2.513955e-07, 2.511005e-07, 
    2.532943e-07, 2.522073e-07, 2.544242e-07, 2.537304e-07, 2.554738e-07, 
    2.543162e-07, 2.557073e-07, 2.554404e-07, 2.562439e-07, 2.560137e-07, 
    2.570418e-07, 2.563502e-07, 2.575751e-07, 2.568766e-07, 2.569859e-07, 
    2.563274e-07, 2.52426e-07, 2.531589e-07, 2.523826e-07, 2.524871e-07, 
    2.524402e-07, 2.518705e-07, 2.515834e-07, 2.509823e-07, 2.510914e-07, 
    2.515329e-07, 2.525341e-07, 2.521942e-07, 2.53051e-07, 2.530317e-07, 
    2.539861e-07, 2.535557e-07, 2.551606e-07, 2.547043e-07, 2.560233e-07, 
    2.556915e-07, 2.560077e-07, 2.559118e-07, 2.560089e-07, 2.555223e-07, 
    2.557308e-07, 2.553027e-07, 2.536363e-07, 2.541258e-07, 2.526661e-07, 
    2.51789e-07, 2.512066e-07, 2.507935e-07, 2.508519e-07, 2.509632e-07, 
    2.515355e-07, 2.520737e-07, 2.524839e-07, 2.527584e-07, 2.530289e-07, 
    2.538478e-07, 2.542815e-07, 2.552529e-07, 2.550776e-07, 2.553746e-07, 
    2.556585e-07, 2.561351e-07, 2.560567e-07, 2.562667e-07, 2.553668e-07, 
    2.559648e-07, 2.549777e-07, 2.552476e-07, 2.531024e-07, 2.522859e-07, 
    2.519389e-07, 2.516353e-07, 2.508968e-07, 2.514068e-07, 2.512057e-07, 
    2.51684e-07, 2.519881e-07, 2.518377e-07, 2.527659e-07, 2.52405e-07, 
    2.543072e-07, 2.534876e-07, 2.556253e-07, 2.551135e-07, 2.557481e-07, 
    2.554243e-07, 2.559791e-07, 2.554798e-07, 2.563449e-07, 2.565333e-07, 
    2.564045e-07, 2.568993e-07, 2.554521e-07, 2.560077e-07, 2.518335e-07, 
    2.51858e-07, 2.519722e-07, 2.514701e-07, 2.514394e-07, 2.509794e-07, 
    2.513887e-07, 2.51563e-07, 2.520057e-07, 2.522676e-07, 2.525165e-07, 
    2.530641e-07, 2.536758e-07, 2.545316e-07, 2.551467e-07, 2.555592e-07, 
    2.553063e-07, 2.555295e-07, 2.552799e-07, 2.55163e-07, 2.564627e-07, 
    2.557327e-07, 2.568281e-07, 2.567675e-07, 2.562717e-07, 2.567743e-07, 
    2.518752e-07, 2.517341e-07, 2.512443e-07, 2.516276e-07, 2.509293e-07, 
    2.513201e-07, 2.515449e-07, 2.524125e-07, 2.526032e-07, 2.5278e-07, 
    2.531293e-07, 2.535777e-07, 2.543646e-07, 2.550495e-07, 2.55675e-07, 
    2.556291e-07, 2.556453e-07, 2.55785e-07, 2.554389e-07, 2.558419e-07, 
    2.559095e-07, 2.557327e-07, 2.567594e-07, 2.56466e-07, 2.567662e-07, 
    2.565752e-07, 2.5178e-07, 2.520174e-07, 2.518891e-07, 2.521304e-07, 
    2.519604e-07, 2.527164e-07, 2.529432e-07, 2.540045e-07, 2.535689e-07, 
    2.542623e-07, 2.536393e-07, 2.537497e-07, 2.542849e-07, 2.53673e-07, 
    2.550117e-07, 2.54104e-07, 2.557905e-07, 2.548836e-07, 2.558473e-07, 
    2.556723e-07, 2.559621e-07, 2.562217e-07, 2.565484e-07, 2.571514e-07, 
    2.570117e-07, 2.575161e-07, 2.523715e-07, 2.526796e-07, 2.526525e-07, 
    2.529749e-07, 2.532135e-07, 2.537306e-07, 2.545603e-07, 2.542482e-07, 
    2.548212e-07, 2.549362e-07, 2.540658e-07, 2.546002e-07, 2.528858e-07, 
    2.531627e-07, 2.529978e-07, 2.523958e-07, 2.543201e-07, 2.533323e-07, 
    2.551569e-07, 2.546214e-07, 2.561847e-07, 2.554071e-07, 2.569349e-07, 
    2.575884e-07, 2.582038e-07, 2.589233e-07, 2.528477e-07, 2.526384e-07, 
    2.530133e-07, 2.535321e-07, 2.540137e-07, 2.546541e-07, 2.547196e-07, 
    2.548396e-07, 2.551505e-07, 2.554119e-07, 2.548775e-07, 2.554775e-07, 
    2.532269e-07, 2.544059e-07, 2.525592e-07, 2.531151e-07, 2.535015e-07, 
    2.53332e-07, 2.542126e-07, 2.544202e-07, 2.552641e-07, 2.548278e-07, 
    2.574271e-07, 2.562766e-07, 2.594713e-07, 2.585779e-07, 2.525652e-07, 
    2.52847e-07, 2.538281e-07, 2.533613e-07, 2.546968e-07, 2.550257e-07, 
    2.552932e-07, 2.556351e-07, 2.55672e-07, 2.558746e-07, 2.555426e-07, 
    2.558615e-07, 2.546554e-07, 2.551943e-07, 2.53716e-07, 2.540757e-07, 
    2.539102e-07, 2.537287e-07, 2.542889e-07, 2.548859e-07, 2.548987e-07, 
    2.550902e-07, 2.556299e-07, 2.547023e-07, 2.575756e-07, 2.558005e-07, 
    2.531544e-07, 2.536974e-07, 2.53775e-07, 2.535646e-07, 2.549928e-07, 
    2.544751e-07, 2.558697e-07, 2.554927e-07, 2.561104e-07, 2.558034e-07, 
    2.557583e-07, 2.553641e-07, 2.551186e-07, 2.544989e-07, 2.539947e-07, 
    2.535951e-07, 2.53688e-07, 2.54127e-07, 2.549225e-07, 2.556753e-07, 
    2.555104e-07, 2.560635e-07, 2.546e-07, 2.552135e-07, 2.549763e-07, 
    2.555948e-07, 2.5424e-07, 2.553935e-07, 2.539452e-07, 2.540721e-07, 
    2.544649e-07, 2.552551e-07, 2.5543e-07, 2.556167e-07, 2.555015e-07, 
    2.549427e-07, 2.548512e-07, 2.544553e-07, 2.54346e-07, 2.540445e-07, 
    2.537949e-07, 2.54023e-07, 2.542625e-07, 2.549429e-07, 2.555564e-07, 
    2.562254e-07, 2.563892e-07, 2.571714e-07, 2.565346e-07, 2.575855e-07, 
    2.56692e-07, 2.582391e-07, 2.554604e-07, 2.566657e-07, 2.544827e-07, 
    2.547178e-07, 2.55143e-07, 2.561186e-07, 2.555919e-07, 2.56208e-07, 
    2.548475e-07, 2.541422e-07, 2.539597e-07, 2.536194e-07, 2.539675e-07, 
    2.539392e-07, 2.542724e-07, 2.541653e-07, 2.549655e-07, 2.545356e-07, 
    2.557571e-07, 2.562031e-07, 2.574633e-07, 2.582363e-07, 2.590236e-07, 
    2.593713e-07, 2.594771e-07, 2.595214e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HTOP =
  0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823 ;

 INT_SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAISHA =
  0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503 ;

 LAISUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAKEICEFRAC =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAKEICETHICK =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAND_UPTAKE =
  7.624269e-08, 7.645139e-08, 7.641083e-08, 7.657911e-08, 7.648578e-08, 
    7.659595e-08, 7.628502e-08, 7.645966e-08, 7.634819e-08, 7.62615e-08, 
    7.690554e-08, 7.658662e-08, 7.723681e-08, 7.70335e-08, 7.754418e-08, 
    7.720516e-08, 7.761253e-08, 7.753444e-08, 7.776953e-08, 7.77022e-08, 
    7.800275e-08, 7.780061e-08, 7.815856e-08, 7.79545e-08, 7.798641e-08, 
    7.779394e-08, 7.665084e-08, 7.686582e-08, 7.663809e-08, 7.666875e-08, 
    7.6655e-08, 7.648769e-08, 7.640334e-08, 7.622676e-08, 7.625883e-08, 
    7.638853e-08, 7.668255e-08, 7.658277e-08, 7.683426e-08, 7.682858e-08, 
    7.710845e-08, 7.698227e-08, 7.745253e-08, 7.731892e-08, 7.7705e-08, 
    7.760792e-08, 7.770044e-08, 7.767239e-08, 7.77008e-08, 7.755842e-08, 
    7.761943e-08, 7.749413e-08, 7.700589e-08, 7.71494e-08, 7.67213e-08, 
    7.646373e-08, 7.629267e-08, 7.617125e-08, 7.618841e-08, 7.622113e-08, 
    7.638929e-08, 7.654739e-08, 7.666784e-08, 7.674839e-08, 7.682777e-08, 
    7.706788e-08, 7.719501e-08, 7.747953e-08, 7.742823e-08, 7.751517e-08, 
    7.759827e-08, 7.773771e-08, 7.771477e-08, 7.777619e-08, 7.75129e-08, 
    7.768788e-08, 7.739899e-08, 7.747801e-08, 7.684923e-08, 7.66097e-08, 
    7.650777e-08, 7.641862e-08, 7.620162e-08, 7.635147e-08, 7.629239e-08, 
    7.643295e-08, 7.652225e-08, 7.647809e-08, 7.67506e-08, 7.664466e-08, 
    7.720254e-08, 7.696229e-08, 7.758857e-08, 7.743876e-08, 7.762448e-08, 
    7.752973e-08, 7.769207e-08, 7.754596e-08, 7.779906e-08, 7.785415e-08, 
    7.78165e-08, 7.796114e-08, 7.753786e-08, 7.770043e-08, 7.647685e-08, 
    7.648405e-08, 7.651761e-08, 7.637008e-08, 7.636106e-08, 7.622587e-08, 
    7.634618e-08, 7.639739e-08, 7.652743e-08, 7.660432e-08, 7.667741e-08, 
    7.683809e-08, 7.701749e-08, 7.72683e-08, 7.744847e-08, 7.75692e-08, 
    7.749518e-08, 7.756054e-08, 7.748747e-08, 7.745323e-08, 7.78335e-08, 
    7.761999e-08, 7.794034e-08, 7.792262e-08, 7.777765e-08, 7.792462e-08, 
    7.648911e-08, 7.644767e-08, 7.630373e-08, 7.641638e-08, 7.621115e-08, 
    7.632602e-08, 7.639206e-08, 7.664685e-08, 7.670285e-08, 7.675474e-08, 
    7.685723e-08, 7.698873e-08, 7.721936e-08, 7.741998e-08, 7.76031e-08, 
    7.758969e-08, 7.759441e-08, 7.76353e-08, 7.7534e-08, 7.765193e-08, 
    7.767171e-08, 7.761997e-08, 7.792025e-08, 7.783448e-08, 7.792224e-08, 
    7.78664e-08, 7.646114e-08, 7.653087e-08, 7.649319e-08, 7.656404e-08, 
    7.651412e-08, 7.673605e-08, 7.680259e-08, 7.711383e-08, 7.698614e-08, 
    7.718939e-08, 7.70068e-08, 7.703915e-08, 7.719597e-08, 7.701667e-08, 
    7.74089e-08, 7.714296e-08, 7.763688e-08, 7.737135e-08, 7.765352e-08, 
    7.760231e-08, 7.768711e-08, 7.776304e-08, 7.785858e-08, 7.803479e-08, 
    7.7994e-08, 7.814135e-08, 7.663483e-08, 7.672524e-08, 7.671731e-08, 
    7.681193e-08, 7.68819e-08, 7.703356e-08, 7.727672e-08, 7.71853e-08, 
    7.735314e-08, 7.738683e-08, 7.713184e-08, 7.728839e-08, 7.678577e-08, 
    7.686698e-08, 7.681864e-08, 7.664195e-08, 7.720634e-08, 7.691673e-08, 
    7.745144e-08, 7.729462e-08, 7.775221e-08, 7.752466e-08, 7.797154e-08, 
    7.816244e-08, 7.834216e-08, 7.855203e-08, 7.677461e-08, 7.671318e-08, 
    7.682319e-08, 7.697533e-08, 7.711654e-08, 7.730418e-08, 7.732339e-08, 
    7.735854e-08, 7.744958e-08, 7.752611e-08, 7.736963e-08, 7.754529e-08, 
    7.688577e-08, 7.723148e-08, 7.668994e-08, 7.685301e-08, 7.696638e-08, 
    7.691667e-08, 7.717485e-08, 7.723568e-08, 7.748282e-08, 7.735509e-08, 
    7.811531e-08, 7.777906e-08, 7.871185e-08, 7.845127e-08, 7.669171e-08, 
    7.677441e-08, 7.706215e-08, 7.692525e-08, 7.731672e-08, 7.741303e-08, 
    7.749135e-08, 7.75914e-08, 7.760222e-08, 7.76615e-08, 7.756436e-08, 
    7.765767e-08, 7.730458e-08, 7.74624e-08, 7.702928e-08, 7.713471e-08, 
    7.708622e-08, 7.703301e-08, 7.719722e-08, 7.737208e-08, 7.737585e-08, 
    7.743191e-08, 7.758979e-08, 7.731831e-08, 7.815863e-08, 7.763973e-08, 
    7.686458e-08, 7.702379e-08, 7.704657e-08, 7.698489e-08, 7.740338e-08, 
    7.725177e-08, 7.766006e-08, 7.754974e-08, 7.77305e-08, 7.764068e-08, 
    7.762746e-08, 7.75121e-08, 7.744025e-08, 7.725872e-08, 7.711099e-08, 
    7.699384e-08, 7.702109e-08, 7.714976e-08, 7.738279e-08, 7.760318e-08, 
    7.755491e-08, 7.771676e-08, 7.728835e-08, 7.7468e-08, 7.739856e-08, 
    7.757962e-08, 7.718286e-08, 7.752063e-08, 7.709649e-08, 7.713369e-08, 
    7.724876e-08, 7.748016e-08, 7.75314e-08, 7.758604e-08, 7.755232e-08, 
    7.738871e-08, 7.736191e-08, 7.724597e-08, 7.721394e-08, 7.71256e-08, 
    7.705243e-08, 7.711927e-08, 7.718945e-08, 7.738879e-08, 7.756837e-08, 
    7.776411e-08, 7.781203e-08, 7.804059e-08, 7.785449e-08, 7.816151e-08, 
    7.790043e-08, 7.835236e-08, 7.754026e-08, 7.789281e-08, 7.725401e-08, 
    7.732286e-08, 7.744735e-08, 7.773286e-08, 7.757877e-08, 7.775899e-08, 
    7.736087e-08, 7.715419e-08, 7.710074e-08, 7.700096e-08, 7.710302e-08, 
    7.709473e-08, 7.719238e-08, 7.7161e-08, 7.739541e-08, 7.72695e-08, 
    7.762712e-08, 7.775758e-08, 7.812591e-08, 7.835159e-08, 7.858132e-08, 
    7.86827e-08, 7.871355e-08, 7.872645e-08 ;

 LAND_USE_FLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC =
  0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203 ;

 LEAFC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC_LOSS =
  8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10 ;

 LEAFN =
  0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507 ;

 LEAF_MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LFC2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LF_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITFALL =
  1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09 ;

 LITHR =
  9.949953e-13, 9.975261e-13, 9.970345e-13, 9.990735e-13, 9.97943e-13, 
    9.992776e-13, 9.95509e-13, 9.97626e-13, 9.96275e-13, 9.952239e-13, 
    1.003024e-12, 9.991646e-13, 1.00703e-12, 1.004573e-12, 1.01074e-12, 
    1.006647e-12, 1.011565e-12, 1.010623e-12, 1.013458e-12, 1.012646e-12, 
    1.016266e-12, 1.013833e-12, 1.018142e-12, 1.015686e-12, 1.01607e-12, 
    1.013752e-12, 9.999428e-13, 1.002544e-12, 9.997884e-13, 1.000159e-12, 
    9.999932e-13, 9.97966e-13, 9.969432e-13, 9.948024e-13, 9.951915e-13, 
    9.96764e-13, 1.000326e-12, 9.991183e-13, 1.002163e-12, 1.002095e-12, 
    1.005479e-12, 1.003954e-12, 1.009635e-12, 1.008022e-12, 1.01268e-12, 
    1.01151e-12, 1.012625e-12, 1.012287e-12, 1.01263e-12, 1.010912e-12, 
    1.011648e-12, 1.010137e-12, 1.004239e-12, 1.005974e-12, 1.000796e-12, 
    9.976748e-13, 9.956017e-13, 9.941288e-13, 9.943371e-13, 9.947339e-13, 
    9.967732e-13, 9.986896e-13, 1.000149e-12, 1.001124e-12, 1.002085e-12, 
    1.004988e-12, 1.006525e-12, 1.009961e-12, 1.009342e-12, 1.010391e-12, 
    1.011393e-12, 1.013074e-12, 1.012798e-12, 1.013538e-12, 1.010364e-12, 
    1.012474e-12, 1.008989e-12, 1.009943e-12, 1.002343e-12, 9.994445e-13, 
    9.982088e-13, 9.971288e-13, 9.944972e-13, 9.963147e-13, 9.955984e-13, 
    9.973029e-13, 9.98385e-13, 9.9785e-13, 1.001151e-12, 9.998679e-13, 
    1.006616e-12, 1.003712e-12, 1.011276e-12, 1.009469e-12, 1.011709e-12, 
    1.010567e-12, 1.012524e-12, 1.010762e-12, 1.013814e-12, 1.014477e-12, 
    1.014024e-12, 1.015766e-12, 1.010665e-12, 1.012625e-12, 9.978348e-13, 
    9.979221e-13, 9.983288e-13, 9.965403e-13, 9.96431e-13, 9.947916e-13, 
    9.962507e-13, 9.968715e-13, 9.98448e-13, 9.993793e-13, 1.000265e-12, 
    1.002209e-12, 1.004379e-12, 1.007411e-12, 1.009586e-12, 1.011043e-12, 
    1.01015e-12, 1.010938e-12, 1.010057e-12, 1.009644e-12, 1.014229e-12, 
    1.011655e-12, 1.015516e-12, 1.015302e-12, 1.013556e-12, 1.015326e-12, 
    9.979834e-13, 9.974813e-13, 9.957359e-13, 9.971019e-13, 9.94613e-13, 
    9.960061e-13, 9.968066e-13, 9.998941e-13, 1.000573e-12, 1.001201e-12, 
    1.002441e-12, 1.004032e-12, 1.006819e-12, 1.009242e-12, 1.011452e-12, 
    1.01129e-12, 1.011347e-12, 1.01184e-12, 1.010618e-12, 1.01204e-12, 
    1.012279e-12, 1.011655e-12, 1.015274e-12, 1.014241e-12, 1.015298e-12, 
    1.014625e-12, 9.976446e-13, 9.984896e-13, 9.980329e-13, 9.988913e-13, 
    9.982864e-13, 1.000974e-12, 1.001779e-12, 1.005544e-12, 1.004e-12, 
    1.006457e-12, 1.00425e-12, 1.004641e-12, 1.006536e-12, 1.00437e-12, 
    1.009108e-12, 1.005896e-12, 1.011859e-12, 1.008654e-12, 1.01206e-12, 
    1.011442e-12, 1.012465e-12, 1.01338e-12, 1.014531e-12, 1.016652e-12, 
    1.016162e-12, 1.017935e-12, 9.997489e-13, 1.000844e-12, 1.000748e-12, 
    1.001893e-12, 1.00274e-12, 1.004574e-12, 1.007512e-12, 1.006408e-12, 
    1.008435e-12, 1.008842e-12, 1.005762e-12, 1.007653e-12, 1.001576e-12, 
    1.002559e-12, 1.001974e-12, 9.99835e-13, 1.006662e-12, 1.003161e-12, 
    1.009622e-12, 1.007729e-12, 1.013249e-12, 1.010505e-12, 1.015891e-12, 
    1.018188e-12, 1.020349e-12, 1.02287e-12, 1.001441e-12, 1.000698e-12, 
    1.002029e-12, 1.003869e-12, 1.005577e-12, 1.007844e-12, 1.008076e-12, 
    1.0085e-12, 1.0096e-12, 1.010523e-12, 1.008634e-12, 1.010754e-12, 
    1.002785e-12, 1.006966e-12, 1.000416e-12, 1.00239e-12, 1.003761e-12, 
    1.00316e-12, 1.006282e-12, 1.007017e-12, 1.01e-12, 1.008459e-12, 
    1.017621e-12, 1.013572e-12, 1.024788e-12, 1.02166e-12, 1.000438e-12, 
    1.001439e-12, 1.004919e-12, 1.003264e-12, 1.007996e-12, 1.009158e-12, 
    1.010104e-12, 1.01131e-12, 1.011441e-12, 1.012156e-12, 1.010984e-12, 
    1.01211e-12, 1.007849e-12, 1.009754e-12, 1.004522e-12, 1.005797e-12, 
    1.005211e-12, 1.004568e-12, 1.006552e-12, 1.008664e-12, 1.00871e-12, 
    1.009386e-12, 1.011289e-12, 1.008015e-12, 1.018141e-12, 1.011892e-12, 
    1.00253e-12, 1.004455e-12, 1.004731e-12, 1.003986e-12, 1.009042e-12, 
    1.007211e-12, 1.012139e-12, 1.010808e-12, 1.012988e-12, 1.011905e-12, 
    1.011745e-12, 1.010354e-12, 1.009487e-12, 1.007295e-12, 1.00551e-12, 
    1.004094e-12, 1.004423e-12, 1.005979e-12, 1.008793e-12, 1.011452e-12, 
    1.01087e-12, 1.012822e-12, 1.007653e-12, 1.009821e-12, 1.008983e-12, 
    1.011168e-12, 1.006379e-12, 1.010455e-12, 1.005335e-12, 1.005785e-12, 
    1.007175e-12, 1.009968e-12, 1.010587e-12, 1.011246e-12, 1.010839e-12, 
    1.008864e-12, 1.008541e-12, 1.007141e-12, 1.006754e-12, 1.005687e-12, 
    1.004802e-12, 1.00561e-12, 1.006458e-12, 1.008866e-12, 1.011033e-12, 
    1.013393e-12, 1.01397e-12, 1.016721e-12, 1.014481e-12, 1.018175e-12, 
    1.015033e-12, 1.020471e-12, 1.010693e-12, 1.014942e-12, 1.007238e-12, 
    1.00807e-12, 1.009572e-12, 1.013015e-12, 1.011158e-12, 1.01333e-12, 
    1.008529e-12, 1.006032e-12, 1.005386e-12, 1.00418e-12, 1.005414e-12, 
    1.005314e-12, 1.006494e-12, 1.006115e-12, 1.008946e-12, 1.007425e-12, 
    1.011741e-12, 1.013314e-12, 1.017749e-12, 1.020462e-12, 1.023222e-12, 
    1.024439e-12, 1.024809e-12, 1.024964e-12 ;

 LITR1C =
  3.066706e-05, 3.066694e-05, 3.066697e-05, 3.066687e-05, 3.066692e-05, 
    3.066687e-05, 3.066704e-05, 3.066694e-05, 3.0667e-05, 3.066705e-05, 
    3.06667e-05, 3.066687e-05, 3.066651e-05, 3.066663e-05, 3.066635e-05, 
    3.066653e-05, 3.066631e-05, 3.066635e-05, 3.066622e-05, 3.066626e-05, 
    3.066609e-05, 3.06662e-05, 3.066601e-05, 3.066612e-05, 3.06661e-05, 
    3.066621e-05, 3.066683e-05, 3.066672e-05, 3.066684e-05, 3.066683e-05, 
    3.066683e-05, 3.066692e-05, 3.066697e-05, 3.066707e-05, 3.066705e-05, 
    3.066698e-05, 3.066682e-05, 3.066687e-05, 3.066674e-05, 3.066674e-05, 
    3.066658e-05, 3.066665e-05, 3.06664e-05, 3.066647e-05, 3.066626e-05, 
    3.066631e-05, 3.066626e-05, 3.066628e-05, 3.066626e-05, 3.066634e-05, 
    3.066631e-05, 3.066637e-05, 3.066664e-05, 3.066656e-05, 3.06668e-05, 
    3.066694e-05, 3.066703e-05, 3.06671e-05, 3.066709e-05, 3.066707e-05, 
    3.066698e-05, 3.066689e-05, 3.066683e-05, 3.066678e-05, 3.066674e-05, 
    3.066661e-05, 3.066654e-05, 3.066638e-05, 3.066641e-05, 3.066636e-05, 
    3.066632e-05, 3.066624e-05, 3.066625e-05, 3.066622e-05, 3.066636e-05, 
    3.066627e-05, 3.066643e-05, 3.066638e-05, 3.066672e-05, 3.066686e-05, 
    3.066691e-05, 3.066696e-05, 3.066708e-05, 3.0667e-05, 3.066703e-05, 
    3.066695e-05, 3.066691e-05, 3.066693e-05, 3.066678e-05, 3.066684e-05, 
    3.066653e-05, 3.066666e-05, 3.066632e-05, 3.06664e-05, 3.06663e-05, 
    3.066635e-05, 3.066627e-05, 3.066635e-05, 3.066621e-05, 3.066618e-05, 
    3.06662e-05, 3.066612e-05, 3.066635e-05, 3.066626e-05, 3.066693e-05, 
    3.066693e-05, 3.066691e-05, 3.066699e-05, 3.066699e-05, 3.066707e-05, 
    3.0667e-05, 3.066698e-05, 3.06669e-05, 3.066686e-05, 3.066682e-05, 
    3.066673e-05, 3.066663e-05, 3.06665e-05, 3.06664e-05, 3.066633e-05, 
    3.066637e-05, 3.066634e-05, 3.066638e-05, 3.06664e-05, 3.066619e-05, 
    3.06663e-05, 3.066613e-05, 3.066614e-05, 3.066622e-05, 3.066614e-05, 
    3.066692e-05, 3.066695e-05, 3.066703e-05, 3.066696e-05, 3.066708e-05, 
    3.066701e-05, 3.066698e-05, 3.066684e-05, 3.06668e-05, 3.066678e-05, 
    3.066672e-05, 3.066665e-05, 3.066652e-05, 3.066642e-05, 3.066631e-05, 
    3.066632e-05, 3.066632e-05, 3.06663e-05, 3.066635e-05, 3.066629e-05, 
    3.066628e-05, 3.06663e-05, 3.066614e-05, 3.066619e-05, 3.066614e-05, 
    3.066617e-05, 3.066694e-05, 3.06669e-05, 3.066692e-05, 3.066688e-05, 
    3.066691e-05, 3.066679e-05, 3.066675e-05, 3.066658e-05, 3.066665e-05, 
    3.066654e-05, 3.066664e-05, 3.066662e-05, 3.066654e-05, 3.066663e-05, 
    3.066642e-05, 3.066656e-05, 3.06663e-05, 3.066644e-05, 3.066628e-05, 
    3.066631e-05, 3.066627e-05, 3.066623e-05, 3.066618e-05, 3.066608e-05, 
    3.06661e-05, 3.066602e-05, 3.066684e-05, 3.066679e-05, 3.06668e-05, 
    3.066675e-05, 3.066671e-05, 3.066663e-05, 3.066649e-05, 3.066654e-05, 
    3.066645e-05, 3.066643e-05, 3.066657e-05, 3.066648e-05, 3.066676e-05, 
    3.066672e-05, 3.066674e-05, 3.066684e-05, 3.066653e-05, 3.066669e-05, 
    3.06664e-05, 3.066648e-05, 3.066623e-05, 3.066636e-05, 3.066611e-05, 
    3.066601e-05, 3.066591e-05, 3.06658e-05, 3.066677e-05, 3.06668e-05, 
    3.066674e-05, 3.066666e-05, 3.066658e-05, 3.066648e-05, 3.066647e-05, 
    3.066645e-05, 3.06664e-05, 3.066636e-05, 3.066644e-05, 3.066635e-05, 
    3.066671e-05, 3.066652e-05, 3.066681e-05, 3.066672e-05, 3.066666e-05, 
    3.066669e-05, 3.066655e-05, 3.066651e-05, 3.066638e-05, 3.066645e-05, 
    3.066603e-05, 3.066622e-05, 3.066571e-05, 3.066585e-05, 3.066681e-05, 
    3.066677e-05, 3.066661e-05, 3.066668e-05, 3.066647e-05, 3.066642e-05, 
    3.066638e-05, 3.066632e-05, 3.066631e-05, 3.066628e-05, 3.066634e-05, 
    3.066628e-05, 3.066648e-05, 3.066639e-05, 3.066663e-05, 3.066657e-05, 
    3.06666e-05, 3.066663e-05, 3.066654e-05, 3.066644e-05, 3.066644e-05, 
    3.066641e-05, 3.066632e-05, 3.066647e-05, 3.066601e-05, 3.06663e-05, 
    3.066672e-05, 3.066663e-05, 3.066662e-05, 3.066665e-05, 3.066642e-05, 
    3.066651e-05, 3.066628e-05, 3.066634e-05, 3.066624e-05, 3.066629e-05, 
    3.06663e-05, 3.066636e-05, 3.06664e-05, 3.06665e-05, 3.066658e-05, 
    3.066665e-05, 3.066663e-05, 3.066656e-05, 3.066643e-05, 3.066631e-05, 
    3.066634e-05, 3.066625e-05, 3.066648e-05, 3.066639e-05, 3.066643e-05, 
    3.066633e-05, 3.066654e-05, 3.066636e-05, 3.066659e-05, 3.066657e-05, 
    3.066651e-05, 3.066638e-05, 3.066635e-05, 3.066632e-05, 3.066634e-05, 
    3.066643e-05, 3.066644e-05, 3.066651e-05, 3.066653e-05, 3.066658e-05, 
    3.066662e-05, 3.066658e-05, 3.066654e-05, 3.066643e-05, 3.066633e-05, 
    3.066623e-05, 3.06662e-05, 3.066607e-05, 3.066618e-05, 3.066601e-05, 
    3.066615e-05, 3.066591e-05, 3.066635e-05, 3.066616e-05, 3.06665e-05, 
    3.066647e-05, 3.06664e-05, 3.066624e-05, 3.066633e-05, 3.066623e-05, 
    3.066644e-05, 3.066656e-05, 3.066659e-05, 3.066664e-05, 3.066659e-05, 
    3.066659e-05, 3.066654e-05, 3.066655e-05, 3.066643e-05, 3.06665e-05, 
    3.06663e-05, 3.066623e-05, 3.066603e-05, 3.066591e-05, 3.066578e-05, 
    3.066572e-05, 3.066571e-05, 3.06657e-05 ;

 LITR1C_TO_SOIL1C =
  6.627068e-13, 6.64392e-13, 6.640647e-13, 6.654226e-13, 6.646697e-13, 
    6.655584e-13, 6.630489e-13, 6.644587e-13, 6.63559e-13, 6.62859e-13, 
    6.680533e-13, 6.654832e-13, 6.707207e-13, 6.690847e-13, 6.731915e-13, 
    6.704659e-13, 6.737406e-13, 6.731136e-13, 6.750013e-13, 6.744609e-13, 
    6.768713e-13, 6.752508e-13, 6.7812e-13, 6.764848e-13, 6.767405e-13, 
    6.751971e-13, 6.660013e-13, 6.677333e-13, 6.658985e-13, 6.661457e-13, 
    6.660349e-13, 6.64685e-13, 6.64004e-13, 6.625783e-13, 6.628374e-13, 
    6.638846e-13, 6.662568e-13, 6.654524e-13, 6.674801e-13, 6.674343e-13, 
    6.696881e-13, 6.686724e-13, 6.724555e-13, 6.713815e-13, 6.744834e-13, 
    6.737039e-13, 6.744467e-13, 6.742216e-13, 6.744496e-13, 6.733062e-13, 
    6.737962e-13, 6.727898e-13, 6.688625e-13, 6.700176e-13, 6.665694e-13, 
    6.644911e-13, 6.631106e-13, 6.621298e-13, 6.622685e-13, 6.625328e-13, 
    6.638907e-13, 6.651669e-13, 6.661385e-13, 6.66788e-13, 6.674278e-13, 
    6.693609e-13, 6.703844e-13, 6.726723e-13, 6.722602e-13, 6.729587e-13, 
    6.736264e-13, 6.747458e-13, 6.745618e-13, 6.750546e-13, 6.729406e-13, 
    6.743458e-13, 6.720253e-13, 6.726603e-13, 6.675995e-13, 6.656696e-13, 
    6.648466e-13, 6.641276e-13, 6.623751e-13, 6.635854e-13, 6.631083e-13, 
    6.642435e-13, 6.64964e-13, 6.646078e-13, 6.668057e-13, 6.659516e-13, 
    6.70445e-13, 6.685113e-13, 6.735485e-13, 6.723448e-13, 6.738369e-13, 
    6.730759e-13, 6.743794e-13, 6.732063e-13, 6.752382e-13, 6.7568e-13, 
    6.75378e-13, 6.765383e-13, 6.731412e-13, 6.744465e-13, 6.645977e-13, 
    6.646558e-13, 6.649267e-13, 6.637356e-13, 6.636629e-13, 6.625712e-13, 
    6.635428e-13, 6.639562e-13, 6.650059e-13, 6.656261e-13, 6.662156e-13, 
    6.675108e-13, 6.689557e-13, 6.709742e-13, 6.724229e-13, 6.73393e-13, 
    6.727984e-13, 6.733234e-13, 6.727364e-13, 6.724613e-13, 6.755143e-13, 
    6.738006e-13, 6.763714e-13, 6.762294e-13, 6.750663e-13, 6.762454e-13, 
    6.646966e-13, 6.643622e-13, 6.632e-13, 6.641096e-13, 6.624522e-13, 
    6.633799e-13, 6.639129e-13, 6.65969e-13, 6.664208e-13, 6.66839e-13, 
    6.676651e-13, 6.687244e-13, 6.705805e-13, 6.721938e-13, 6.736653e-13, 
    6.735575e-13, 6.735955e-13, 6.739238e-13, 6.731101e-13, 6.740573e-13, 
    6.74216e-13, 6.738007e-13, 6.762103e-13, 6.755224e-13, 6.762264e-13, 
    6.757786e-13, 6.64471e-13, 6.650337e-13, 6.647296e-13, 6.653012e-13, 
    6.648984e-13, 6.666881e-13, 6.672243e-13, 6.697311e-13, 6.687034e-13, 
    6.703393e-13, 6.688698e-13, 6.691302e-13, 6.703918e-13, 6.689494e-13, 
    6.721045e-13, 6.699654e-13, 6.739365e-13, 6.718024e-13, 6.740701e-13, 
    6.736589e-13, 6.743398e-13, 6.749491e-13, 6.757157e-13, 6.771284e-13, 
    6.768016e-13, 6.779825e-13, 6.658723e-13, 6.666012e-13, 6.665374e-13, 
    6.673001e-13, 6.678638e-13, 6.690854e-13, 6.71042e-13, 6.703066e-13, 
    6.716567e-13, 6.719275e-13, 6.698765e-13, 6.711357e-13, 6.670891e-13, 
    6.677433e-13, 6.673541e-13, 6.659296e-13, 6.704756e-13, 6.681441e-13, 
    6.724467e-13, 6.71186e-13, 6.748622e-13, 6.730348e-13, 6.766215e-13, 
    6.781508e-13, 6.795903e-13, 6.812685e-13, 6.669992e-13, 6.665041e-13, 
    6.673909e-13, 6.686162e-13, 6.697533e-13, 6.712628e-13, 6.714175e-13, 
    6.716999e-13, 6.724319e-13, 6.730468e-13, 6.717889e-13, 6.732009e-13, 
    6.678941e-13, 6.70678e-13, 6.663165e-13, 6.676307e-13, 6.685442e-13, 
    6.681439e-13, 6.702227e-13, 6.707121e-13, 6.726987e-13, 6.716723e-13, 
    6.777732e-13, 6.750773e-13, 6.825462e-13, 6.80463e-13, 6.66331e-13, 
    6.669977e-13, 6.693152e-13, 6.682131e-13, 6.713638e-13, 6.721381e-13, 
    6.727676e-13, 6.735711e-13, 6.736582e-13, 6.741341e-13, 6.733541e-13, 
    6.741034e-13, 6.712661e-13, 6.725348e-13, 6.69051e-13, 6.698995e-13, 
    6.695094e-13, 6.69081e-13, 6.704026e-13, 6.718086e-13, 6.718393e-13, 
    6.722896e-13, 6.73557e-13, 6.713766e-13, 6.781195e-13, 6.739581e-13, 
    6.677244e-13, 6.690063e-13, 6.6919e-13, 6.686935e-13, 6.720604e-13, 
    6.708414e-13, 6.741225e-13, 6.732367e-13, 6.746881e-13, 6.73967e-13, 
    6.738608e-13, 6.729342e-13, 6.723568e-13, 6.708971e-13, 6.697085e-13, 
    6.687656e-13, 6.68985e-13, 6.700206e-13, 6.718947e-13, 6.736658e-13, 
    6.732779e-13, 6.745778e-13, 6.711356e-13, 6.725797e-13, 6.720215e-13, 
    6.734766e-13, 6.70287e-13, 6.730017e-13, 6.69592e-13, 6.698914e-13, 
    6.708171e-13, 6.726771e-13, 6.730892e-13, 6.73528e-13, 6.732574e-13, 
    6.719424e-13, 6.717271e-13, 6.707948e-13, 6.70537e-13, 6.698263e-13, 
    6.692373e-13, 6.697753e-13, 6.703399e-13, 6.719432e-13, 6.733861e-13, 
    6.749578e-13, 6.753423e-13, 6.771742e-13, 6.756823e-13, 6.781425e-13, 
    6.760499e-13, 6.79671e-13, 6.731598e-13, 6.759895e-13, 6.708595e-13, 
    6.714132e-13, 6.724136e-13, 6.747065e-13, 6.734697e-13, 6.749163e-13, 
    6.717186e-13, 6.70056e-13, 6.696262e-13, 6.688229e-13, 6.696446e-13, 
    6.695778e-13, 6.703637e-13, 6.701113e-13, 6.719964e-13, 6.709841e-13, 
    6.73858e-13, 6.749051e-13, 6.778585e-13, 6.796654e-13, 6.815032e-13, 
    6.823134e-13, 6.8256e-13, 6.82663e-13 ;

 LITR1C_vr =
  0.001751121, 0.001751114, 0.001751115, 0.00175111, 0.001751113, 0.00175111, 
    0.001751119, 0.001751114, 0.001751117, 0.00175112, 0.0017511, 0.00175111, 
    0.00175109, 0.001751096, 0.00175108, 0.001751091, 0.001751078, 
    0.00175108, 0.001751073, 0.001751075, 0.001751066, 0.001751072, 
    0.001751061, 0.001751067, 0.001751066, 0.001751072, 0.001751108, 
    0.001751101, 0.001751108, 0.001751107, 0.001751108, 0.001751113, 
    0.001751116, 0.001751121, 0.00175112, 0.001751116, 0.001751107, 
    0.00175111, 0.001751102, 0.001751102, 0.001751094, 0.001751098, 
    0.001751083, 0.001751087, 0.001751075, 0.001751078, 0.001751075, 
    0.001751076, 0.001751075, 0.00175108, 0.001751078, 0.001751082, 
    0.001751097, 0.001751092, 0.001751106, 0.001751114, 0.001751119, 
    0.001751123, 0.001751122, 0.001751121, 0.001751116, 0.001751111, 
    0.001751107, 0.001751105, 0.001751102, 0.001751095, 0.001751091, 
    0.001751082, 0.001751084, 0.001751081, 0.001751078, 0.001751074, 
    0.001751075, 0.001751073, 0.001751081, 0.001751075, 0.001751085, 
    0.001751082, 0.001751102, 0.001751109, 0.001751112, 0.001751115, 
    0.001751122, 0.001751117, 0.001751119, 0.001751115, 0.001751112, 
    0.001751113, 0.001751105, 0.001751108, 0.001751091, 0.001751098, 
    0.001751079, 0.001751083, 0.001751077, 0.001751081, 0.001751075, 
    0.00175108, 0.001751072, 0.00175107, 0.001751072, 0.001751067, 
    0.00175108, 0.001751075, 0.001751113, 0.001751113, 0.001751112, 
    0.001751117, 0.001751117, 0.001751121, 0.001751118, 0.001751116, 
    0.001751112, 0.001751109, 0.001751107, 0.001751102, 0.001751096, 
    0.001751089, 0.001751083, 0.001751079, 0.001751082, 0.001751079, 
    0.001751082, 0.001751083, 0.001751071, 0.001751078, 0.001751068, 
    0.001751068, 0.001751073, 0.001751068, 0.001751113, 0.001751114, 
    0.001751119, 0.001751115, 0.001751122, 0.001751118, 0.001751116, 
    0.001751108, 0.001751106, 0.001751105, 0.001751101, 0.001751097, 
    0.00175109, 0.001751084, 0.001751078, 0.001751079, 0.001751078, 
    0.001751077, 0.00175108, 0.001751077, 0.001751076, 0.001751078, 
    0.001751068, 0.001751071, 0.001751068, 0.00175107, 0.001751114, 
    0.001751112, 0.001751113, 0.001751111, 0.001751112, 0.001751105, 
    0.001751103, 0.001751093, 0.001751098, 0.001751091, 0.001751097, 
    0.001751096, 0.001751091, 0.001751096, 0.001751084, 0.001751092, 
    0.001751077, 0.001751085, 0.001751077, 0.001751078, 0.001751075, 
    0.001751073, 0.00175107, 0.001751065, 0.001751066, 0.001751061, 
    0.001751108, 0.001751106, 0.001751106, 0.001751103, 0.001751101, 
    0.001751096, 0.001751088, 0.001751091, 0.001751086, 0.001751085, 
    0.001751093, 0.001751088, 0.001751104, 0.001751101, 0.001751103, 
    0.001751108, 0.001751091, 0.0017511, 0.001751083, 0.001751088, 
    0.001751074, 0.001751081, 0.001751067, 0.001751061, 0.001751055, 
    0.001751049, 0.001751104, 0.001751106, 0.001751103, 0.001751098, 
    0.001751093, 0.001751087, 0.001751087, 0.001751086, 0.001751083, 
    0.001751081, 0.001751086, 0.00175108, 0.001751101, 0.00175109, 
    0.001751107, 0.001751102, 0.001751098, 0.0017511, 0.001751092, 
    0.00175109, 0.001751082, 0.001751086, 0.001751062, 0.001751073, 
    0.001751044, 0.001751052, 0.001751107, 0.001751104, 0.001751095, 
    0.001751099, 0.001751087, 0.001751084, 0.001751082, 0.001751079, 
    0.001751078, 0.001751076, 0.001751079, 0.001751076, 0.001751087, 
    0.001751083, 0.001751096, 0.001751093, 0.001751094, 0.001751096, 
    0.001751091, 0.001751085, 0.001751085, 0.001751084, 0.001751079, 
    0.001751087, 0.001751061, 0.001751077, 0.001751101, 0.001751096, 
    0.001751096, 0.001751098, 0.001751084, 0.001751089, 0.001751076, 
    0.00175108, 0.001751074, 0.001751077, 0.001751077, 0.001751081, 
    0.001751083, 0.001751089, 0.001751094, 0.001751097, 0.001751096, 
    0.001751092, 0.001751085, 0.001751078, 0.00175108, 0.001751075, 
    0.001751088, 0.001751082, 0.001751085, 0.001751079, 0.001751091, 
    0.001751081, 0.001751094, 0.001751093, 0.001751089, 0.001751082, 
    0.00175108, 0.001751079, 0.00175108, 0.001751085, 0.001751086, 
    0.001751089, 0.00175109, 0.001751093, 0.001751095, 0.001751093, 
    0.001751091, 0.001751085, 0.001751079, 0.001751073, 0.001751072, 
    0.001751065, 0.00175107, 0.001751061, 0.001751069, 0.001751055, 
    0.00175108, 0.001751069, 0.001751089, 0.001751087, 0.001751083, 
    0.001751074, 0.001751079, 0.001751073, 0.001751086, 0.001751092, 
    0.001751094, 0.001751097, 0.001751094, 0.001751094, 0.001751091, 
    0.001751092, 0.001751085, 0.001751089, 0.001751077, 0.001751073, 
    0.001751062, 0.001751055, 0.001751048, 0.001751045, 0.001751044, 
    0.001751043,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N =
  9.732586e-07, 9.732549e-07, 9.732556e-07, 9.732527e-07, 9.732543e-07, 
    9.732523e-07, 9.732578e-07, 9.732547e-07, 9.732566e-07, 9.732582e-07, 
    9.73247e-07, 9.732526e-07, 9.732412e-07, 9.732447e-07, 9.732358e-07, 
    9.732418e-07, 9.732347e-07, 9.732361e-07, 9.73232e-07, 9.732331e-07, 
    9.73228e-07, 9.732314e-07, 9.732253e-07, 9.732288e-07, 9.732282e-07, 
    9.732315e-07, 9.732514e-07, 9.732477e-07, 9.732516e-07, 9.732511e-07, 
    9.732513e-07, 9.732543e-07, 9.732557e-07, 9.732588e-07, 9.732582e-07, 
    9.73256e-07, 9.732508e-07, 9.732526e-07, 9.732482e-07, 9.732483e-07, 
    9.732435e-07, 9.732456e-07, 9.732374e-07, 9.732398e-07, 9.732331e-07, 
    9.732348e-07, 9.732332e-07, 9.732337e-07, 9.732332e-07, 9.732356e-07, 
    9.732346e-07, 9.732368e-07, 9.732453e-07, 9.732428e-07, 9.732502e-07, 
    9.732547e-07, 9.732577e-07, 9.732598e-07, 9.732595e-07, 9.732589e-07, 
    9.73256e-07, 9.732532e-07, 9.732511e-07, 9.732497e-07, 9.732483e-07, 
    9.732441e-07, 9.73242e-07, 9.73237e-07, 9.732379e-07, 9.732364e-07, 
    9.732349e-07, 9.732325e-07, 9.732329e-07, 9.732319e-07, 9.732364e-07, 
    9.732335e-07, 9.732385e-07, 9.732371e-07, 9.73248e-07, 9.732521e-07, 
    9.732539e-07, 9.732555e-07, 9.732593e-07, 9.732566e-07, 9.732577e-07, 
    9.732552e-07, 9.732537e-07, 9.732544e-07, 9.732497e-07, 9.732515e-07, 
    9.732419e-07, 9.73246e-07, 9.732352e-07, 9.732378e-07, 9.732345e-07, 
    9.732362e-07, 9.732333e-07, 9.732358e-07, 9.732315e-07, 9.732305e-07, 
    9.732312e-07, 9.732287e-07, 9.73236e-07, 9.732332e-07, 9.732545e-07, 
    9.732544e-07, 9.732537e-07, 9.732563e-07, 9.732564e-07, 9.732588e-07, 
    9.732568e-07, 9.732559e-07, 9.732536e-07, 9.732522e-07, 9.73251e-07, 
    9.732481e-07, 9.732451e-07, 9.732407e-07, 9.732375e-07, 9.732355e-07, 
    9.732368e-07, 9.732356e-07, 9.732369e-07, 9.732374e-07, 9.732308e-07, 
    9.732346e-07, 9.73229e-07, 9.732294e-07, 9.732319e-07, 9.732292e-07, 
    9.732543e-07, 9.732549e-07, 9.732574e-07, 9.732555e-07, 9.73259e-07, 
    9.732571e-07, 9.73256e-07, 9.732515e-07, 9.732505e-07, 9.732496e-07, 
    9.732478e-07, 9.732455e-07, 9.732415e-07, 9.73238e-07, 9.732348e-07, 
    9.73235e-07, 9.73235e-07, 9.732344e-07, 9.732361e-07, 9.73234e-07, 
    9.732337e-07, 9.732346e-07, 9.732294e-07, 9.732308e-07, 9.732294e-07, 
    9.732303e-07, 9.732547e-07, 9.732535e-07, 9.732541e-07, 9.732529e-07, 
    9.732538e-07, 9.732499e-07, 9.732488e-07, 9.732433e-07, 9.732456e-07, 
    9.732421e-07, 9.732453e-07, 9.732447e-07, 9.73242e-07, 9.732451e-07, 
    9.732382e-07, 9.732429e-07, 9.732343e-07, 9.732389e-07, 9.73234e-07, 
    9.732349e-07, 9.732335e-07, 9.732321e-07, 9.732304e-07, 9.732274e-07, 
    9.732281e-07, 9.732255e-07, 9.732516e-07, 9.732502e-07, 9.732503e-07, 
    9.732486e-07, 9.732474e-07, 9.732447e-07, 9.732405e-07, 9.732421e-07, 
    9.732393e-07, 9.732386e-07, 9.73243e-07, 9.732403e-07, 9.73249e-07, 
    9.732477e-07, 9.732485e-07, 9.732515e-07, 9.732418e-07, 9.732468e-07, 
    9.732375e-07, 9.732403e-07, 9.732323e-07, 9.732362e-07, 9.732285e-07, 
    9.732252e-07, 9.732221e-07, 9.732184e-07, 9.732493e-07, 9.732503e-07, 
    9.732485e-07, 9.732457e-07, 9.732433e-07, 9.7324e-07, 9.732397e-07, 
    9.732391e-07, 9.732375e-07, 9.732362e-07, 9.732389e-07, 9.732358e-07, 
    9.732473e-07, 9.732413e-07, 9.732507e-07, 9.732479e-07, 9.73246e-07, 
    9.732468e-07, 9.732423e-07, 9.732413e-07, 9.73237e-07, 9.732391e-07, 
    9.73226e-07, 9.732319e-07, 9.732157e-07, 9.732202e-07, 9.732507e-07, 
    9.732493e-07, 9.732443e-07, 9.732466e-07, 9.732398e-07, 9.732381e-07, 
    9.732368e-07, 9.73235e-07, 9.732349e-07, 9.732339e-07, 9.732355e-07, 
    9.732339e-07, 9.7324e-07, 9.732373e-07, 9.732448e-07, 9.73243e-07, 
    9.732438e-07, 9.732448e-07, 9.732419e-07, 9.732389e-07, 9.732388e-07, 
    9.732379e-07, 9.732352e-07, 9.732398e-07, 9.732253e-07, 9.732343e-07, 
    9.732477e-07, 9.732449e-07, 9.732445e-07, 9.732456e-07, 9.732383e-07, 
    9.73241e-07, 9.732339e-07, 9.732358e-07, 9.732327e-07, 9.732343e-07, 
    9.732345e-07, 9.732364e-07, 9.732377e-07, 9.732408e-07, 9.732435e-07, 
    9.732454e-07, 9.732449e-07, 9.732428e-07, 9.732387e-07, 9.732348e-07, 
    9.732357e-07, 9.732329e-07, 9.732403e-07, 9.732372e-07, 9.732385e-07, 
    9.732353e-07, 9.732422e-07, 9.732363e-07, 9.732437e-07, 9.73243e-07, 
    9.732411e-07, 9.73237e-07, 9.732361e-07, 9.732352e-07, 9.732357e-07, 
    9.732386e-07, 9.73239e-07, 9.732411e-07, 9.732416e-07, 9.732431e-07, 
    9.732445e-07, 9.732432e-07, 9.732421e-07, 9.732386e-07, 9.732355e-07, 
    9.732321e-07, 9.732313e-07, 9.732273e-07, 9.732305e-07, 9.732252e-07, 
    9.732297e-07, 9.732219e-07, 9.73236e-07, 9.732298e-07, 9.73241e-07, 
    9.732397e-07, 9.732375e-07, 9.732327e-07, 9.732353e-07, 9.732322e-07, 
    9.73239e-07, 9.732427e-07, 9.732436e-07, 9.732453e-07, 9.732436e-07, 
    9.732437e-07, 9.73242e-07, 9.732425e-07, 9.732385e-07, 9.732406e-07, 
    9.732345e-07, 9.732322e-07, 9.732258e-07, 9.732219e-07, 9.73218e-07, 
    9.732162e-07, 9.732156e-07, 9.732155e-07 ;

 LITR1N_TNDNCY_VERT_TRANS =
  5.097883e-25, 4.166539e-25, -3.235195e-25, 9.803622e-27, 1.073497e-24, 
    2.156797e-25, -2.941087e-26, 6.47039e-25, -3.431268e-25, 1.176435e-25, 
    4.901811e-25, -5.882173e-26, -6.862535e-26, -1.02938e-25, 1.56858e-25, 
    3.921449e-25, 2.156797e-25, 2.646978e-25, 7.107626e-25, -3.235195e-25, 
    -4.509666e-25, 4.705739e-25, 3.62734e-25, 1.450936e-24, -1.612696e-24, 
    3.137159e-25, -4.950829e-25, 2.745014e-25, -5.490028e-25, 2.254833e-25, 
    -6.617445e-25, -1.519561e-25, 4.117521e-25, 2.450906e-25, -5.19592e-25, 
    3.823413e-25, -1.666616e-25, 3.333231e-25, -3.039123e-25, 1.960724e-26, 
    1.960724e-26, -1.068595e-24, -4.901811e-26, -2.548942e-25, 2.548942e-25, 
    -3.725376e-25, -3.529304e-25, -8.235043e-25, -5.391992e-25, 9.803622e-26, 
    1.960724e-26, 2.254833e-25, 1.225453e-25, -6.862535e-26, 4.509666e-25, 
    2.843051e-25, 2.156797e-25, 2.548942e-25, 1.862688e-25, 9.803622e-26, 
    -6.372354e-26, 7.450753e-25, -9.803622e-26, 5.637083e-25, 2.205815e-25, 
    5.882173e-26, -1.323489e-25, -7.842898e-26, -2.156797e-25, -1.058791e-24, 
    8.82326e-26, -4.901811e-26, -2.352869e-25, 3.431268e-25, 2.058761e-25, 
    6.372354e-26, 4.509666e-25, -3.061136e-41, 5.539047e-25, 1.764652e-25, 
    -1.470543e-25, -5.097883e-25, -2.058761e-25, 5.539047e-25, -1.960724e-26, 
    -3.431268e-25, 4.509666e-25, 5.490028e-25, -1.470543e-25, -1.372507e-25, 
    4.509666e-25, -2.990105e-25, -3.039123e-25, 3.235195e-25, 1.519561e-25, 
    -3.235195e-25, 3.578322e-25, -1.960724e-26, 9.803622e-26, -1.666616e-25, 
    -2.450906e-25, 4.705739e-25, -2.450906e-25, -9.803622e-27, -6.372354e-26, 
    -3.088141e-25, -1.274471e-25, 4.901811e-26, 4.41163e-25, -7.058608e-25, 
    4.901811e-26, -6.421373e-25, -3.62734e-25, 1.068595e-24, 6.813517e-25, 
    -9.803622e-27, 7.744861e-25, 5.588064e-25, -5.882173e-26, -9.803622e-26, 
    5.44101e-25, 3.823413e-25, 5.931191e-25, -6.47039e-25, -2.058761e-25, 
    1.078398e-24, -3.38225e-25, 4.65672e-25, 3.039123e-25, 5.735119e-25, 
    -1.960724e-26, -1.274471e-25, 7.842898e-25, -1.666616e-25, 1.960724e-26, 
    9.803622e-27, 0, -2.352869e-25, 2.058761e-25, 2.745014e-25, 5.588064e-25, 
    6.078246e-25, -3.823413e-25, -4.803775e-25, -1.372507e-25, -3.823413e-25, 
    5.784137e-25, -3.235195e-25, 4.705739e-25, -6.47039e-25, -1.024478e-24, 
    -1.470543e-25, 6.176282e-25, -2.450906e-25, -2.254833e-25, -1.176435e-25, 
    7.058608e-25, 6.078246e-25, -1.862688e-25, 1.666616e-25, -3.431268e-25, 
    5.882173e-26, -1.862688e-25, 1.56858e-25, -1.470543e-25, -4.362612e-25, 
    4.117521e-25, 5.342974e-25, -5.19592e-25, 7.00959e-25, -1.960724e-25, 
    -1.078398e-24, -2.009742e-25, -5.391992e-26, 1.274471e-25, 4.215557e-25, 
    -1.862688e-25, 9.803622e-26, 2.254833e-25, -6.862535e-26, -4.705739e-25, 
    -6.862535e-26, 1.274471e-25, 8.431115e-25, 2.646978e-25, -5.490028e-25, 
    1.274471e-25, 9.313441e-25, 8.676206e-25, -2.450905e-26, -3.774394e-25, 
    -3.235195e-25, 7.156644e-25, 2.990105e-25, -8.82326e-26, -1.666616e-25, 
    -6.078246e-25, -3.38225e-25, 5.882173e-26, 1.372507e-25, 6.176282e-25, 
    -1.960724e-25, -1.666616e-25, 9.803622e-27, 4.509666e-25, -1.862688e-25, 
    6.960572e-25, 6.813517e-25, 3.529304e-25, 5.882173e-26, 7.352717e-25, 
    7.940934e-25, 2.646978e-25, 3.431268e-25, 7.646825e-25, 2.450906e-25, 
    1.960724e-25, -1.56858e-25, -7.107626e-25, -1.470543e-26, 8.82326e-26, 
    2.843051e-25, 1.323489e-25, 9.803622e-27, -2.107779e-25, -1.764652e-25, 
    1.176435e-25, -4.901811e-26, -1.470543e-25, 2.205815e-25, 9.803622e-26, 
    4.558684e-25, -5.882173e-26, -2.254833e-25, -1.274471e-25, 5.097883e-25, 
    1.274471e-25, 7.842898e-26, 5.735119e-25, 3.039123e-25, 6.960572e-25, 
    -1.764652e-25, 6.862535e-26, -7.205662e-25, -2.695996e-25, -1.519561e-25, 
    6.960572e-25, 7.352717e-25, 4.215557e-25, -2.058761e-25, 1.470543e-26, 
    -3.921449e-25, -3.921449e-25, 3.039123e-25, 3.431268e-26, -5.98021e-25, 
    2.352869e-25, -3.823413e-25, -9.803622e-27, 3.235195e-25, -2.205815e-25, 
    2.450906e-25, 4.607703e-25, 2.107779e-25, -5.048866e-25, 7.352717e-26, 
    1.56858e-25, -1.176435e-25, -1.666616e-25, -4.803775e-25, -1.078398e-25, 
    -6.47039e-25, -1.519561e-25, 1.372507e-25, -4.509666e-25, 5.882173e-26, 
    4.509666e-25, 5.19592e-25, -6.862535e-26, 4.41163e-25, 2.303851e-25, 
    9.803622e-27, -5.19592e-25, 4.41163e-26, -5.097883e-25, 3.970467e-25, 
    1.323489e-25, 1.02938e-25, 1.56858e-25, 3.921449e-25, -5.882173e-26, 
    3.529304e-25, -1.078398e-25, 5.98021e-25, 9.509513e-25, -1.470543e-25, 
    3.529304e-25, 1.372507e-25, 1.666616e-25, 3.480286e-25, 1.274471e-25, 
    -1.862688e-25, 6.862535e-26, 1.347998e-24, -6.2253e-25, 3.921449e-26, 
    -1.323489e-25, 4.901811e-25, -8.82326e-25, -5.146902e-25, -2.646978e-25, 
    7.842898e-25, -5.490028e-25, -1.960724e-25, -1.274471e-25, 2.450906e-25, 
    -7.352717e-26, -3.921449e-26, -3.284213e-25, -6.960572e-25, 1.960724e-25, 
    -9.509513e-25, -9.803622e-27, 5.588064e-25, 9.803622e-26, 1.372507e-25, 
    -1.274471e-25, 5.19592e-25, 8.03897e-25, 5.882173e-26, 5.490028e-25, 
    -3.970467e-25, -6.176282e-25, 6.862535e-25, 4.705739e-25, -2.107779e-25, 
    -2.058761e-25, -1.078398e-25,
  9.436424e-32, 9.436387e-32, 9.436394e-32, 9.436365e-32, 9.436381e-32, 
    9.436362e-32, 9.436416e-32, 9.436386e-32, 9.436406e-32, 9.43642e-32, 
    9.436308e-32, 9.436364e-32, 9.43625e-32, 9.436286e-32, 9.436196e-32, 
    9.436256e-32, 9.436185e-32, 9.436198e-32, 9.436157e-32, 9.436169e-32, 
    9.436116e-32, 9.436152e-32, 9.436089e-32, 9.436125e-32, 9.436119e-32, 
    9.436153e-32, 9.436352e-32, 9.436314e-32, 9.436354e-32, 9.436349e-32, 
    9.436351e-32, 9.436381e-32, 9.436396e-32, 9.436427e-32, 9.436421e-32, 
    9.436398e-32, 9.436347e-32, 9.436364e-32, 9.43632e-32, 9.436321e-32, 
    9.436272e-32, 9.436294e-32, 9.436212e-32, 9.436236e-32, 9.436168e-32, 
    9.436185e-32, 9.436169e-32, 9.436174e-32, 9.436169e-32, 9.436194e-32, 
    9.436183e-32, 9.436205e-32, 9.43629e-32, 9.436265e-32, 9.43634e-32, 
    9.436385e-32, 9.436415e-32, 9.436436e-32, 9.436433e-32, 9.436427e-32, 
    9.436398e-32, 9.43637e-32, 9.436349e-32, 9.436335e-32, 9.436321e-32, 
    9.436279e-32, 9.436257e-32, 9.436207e-32, 9.436216e-32, 9.436202e-32, 
    9.436187e-32, 9.436163e-32, 9.436166e-32, 9.436156e-32, 9.436202e-32, 
    9.436171e-32, 9.436222e-32, 9.436208e-32, 9.436317e-32, 9.43636e-32, 
    9.436377e-32, 9.436393e-32, 9.436431e-32, 9.436405e-32, 9.436415e-32, 
    9.43639e-32, 9.436375e-32, 9.436383e-32, 9.436335e-32, 9.436353e-32, 
    9.436256e-32, 9.436298e-32, 9.436189e-32, 9.436214e-32, 9.436182e-32, 
    9.436199e-32, 9.43617e-32, 9.436196e-32, 9.436152e-32, 9.436142e-32, 
    9.436149e-32, 9.436123e-32, 9.436197e-32, 9.436169e-32, 9.436383e-32, 
    9.436381e-32, 9.436376e-32, 9.436401e-32, 9.436403e-32, 9.436427e-32, 
    9.436406e-32, 9.436397e-32, 9.436374e-32, 9.43636e-32, 9.436347e-32, 
    9.43632e-32, 9.436288e-32, 9.436244e-32, 9.436213e-32, 9.436192e-32, 
    9.436205e-32, 9.436193e-32, 9.436206e-32, 9.436212e-32, 9.436146e-32, 
    9.436183e-32, 9.436127e-32, 9.43613e-32, 9.436156e-32, 9.43613e-32, 
    9.436381e-32, 9.436388e-32, 9.436413e-32, 9.436393e-32, 9.436429e-32, 
    9.436409e-32, 9.436397e-32, 9.436353e-32, 9.436343e-32, 9.436334e-32, 
    9.436316e-32, 9.436293e-32, 9.436253e-32, 9.436218e-32, 9.436186e-32, 
    9.436188e-32, 9.436187e-32, 9.43618e-32, 9.436198e-32, 9.436177e-32, 
    9.436174e-32, 9.436183e-32, 9.436131e-32, 9.436146e-32, 9.43613e-32, 
    9.43614e-32, 9.436386e-32, 9.436373e-32, 9.43638e-32, 9.436367e-32, 
    9.436376e-32, 9.436337e-32, 9.436326e-32, 9.436271e-32, 9.436294e-32, 
    9.436258e-32, 9.43629e-32, 9.436284e-32, 9.436257e-32, 9.436289e-32, 
    9.43622e-32, 9.436266e-32, 9.43618e-32, 9.436226e-32, 9.436177e-32, 
    9.436186e-32, 9.436172e-32, 9.436158e-32, 9.436142e-32, 9.436111e-32, 
    9.436118e-32, 9.436092e-32, 9.436355e-32, 9.436339e-32, 9.436341e-32, 
    9.436324e-32, 9.436312e-32, 9.436286e-32, 9.436243e-32, 9.436259e-32, 
    9.43623e-32, 9.436224e-32, 9.436268e-32, 9.436241e-32, 9.436329e-32, 
    9.436314e-32, 9.436323e-32, 9.436354e-32, 9.436255e-32, 9.436306e-32, 
    9.436213e-32, 9.43624e-32, 9.43616e-32, 9.4362e-32, 9.436122e-32, 
    9.436089e-32, 9.436058e-32, 9.436021e-32, 9.436331e-32, 9.436341e-32, 
    9.436322e-32, 9.436296e-32, 9.436271e-32, 9.436238e-32, 9.436234e-32, 
    9.436229e-32, 9.436213e-32, 9.436199e-32, 9.436227e-32, 9.436196e-32, 
    9.436311e-32, 9.436251e-32, 9.436346e-32, 9.436317e-32, 9.436297e-32, 
    9.436306e-32, 9.436261e-32, 9.43625e-32, 9.436207e-32, 9.436229e-32, 
    9.436097e-32, 9.436155e-32, 9.435993e-32, 9.436039e-32, 9.436345e-32, 
    9.436331e-32, 9.43628e-32, 9.436304e-32, 9.436236e-32, 9.436219e-32, 
    9.436206e-32, 9.436188e-32, 9.436186e-32, 9.436176e-32, 9.436193e-32, 
    9.436176e-32, 9.436238e-32, 9.43621e-32, 9.436286e-32, 9.436268e-32, 
    9.436276e-32, 9.436286e-32, 9.436257e-32, 9.436226e-32, 9.436226e-32, 
    9.436216e-32, 9.436189e-32, 9.436236e-32, 9.436089e-32, 9.43618e-32, 
    9.436315e-32, 9.436287e-32, 9.436283e-32, 9.436294e-32, 9.436221e-32, 
    9.436247e-32, 9.436176e-32, 9.436195e-32, 9.436164e-32, 9.436179e-32, 
    9.436182e-32, 9.436202e-32, 9.436214e-32, 9.436246e-32, 9.436272e-32, 
    9.436292e-32, 9.436287e-32, 9.436265e-32, 9.436224e-32, 9.436186e-32, 
    9.436195e-32, 9.436166e-32, 9.436241e-32, 9.43621e-32, 9.436222e-32, 
    9.43619e-32, 9.436259e-32, 9.4362e-32, 9.436274e-32, 9.436268e-32, 
    9.436248e-32, 9.436207e-32, 9.436199e-32, 9.436189e-32, 9.436195e-32, 
    9.436223e-32, 9.436228e-32, 9.436248e-32, 9.436254e-32, 9.436269e-32, 
    9.436282e-32, 9.43627e-32, 9.436258e-32, 9.436223e-32, 9.436192e-32, 
    9.436158e-32, 9.43615e-32, 9.43611e-32, 9.436142e-32, 9.436089e-32, 
    9.436135e-32, 9.436056e-32, 9.436197e-32, 9.436136e-32, 9.436247e-32, 
    9.436235e-32, 9.436213e-32, 9.436163e-32, 9.43619e-32, 9.436159e-32, 
    9.436228e-32, 9.436264e-32, 9.436274e-32, 9.436291e-32, 9.436273e-32, 
    9.436274e-32, 9.436257e-32, 9.436263e-32, 9.436222e-32, 9.436244e-32, 
    9.436182e-32, 9.436159e-32, 9.436095e-32, 9.436056e-32, 9.436016e-32, 
    9.435998e-32, 9.435993e-32, 9.435991e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N_TO_SOIL1N =
  4.67374e-14, 4.685625e-14, 4.683317e-14, 4.692893e-14, 4.687584e-14, 
    4.693851e-14, 4.676153e-14, 4.686095e-14, 4.67975e-14, 4.674813e-14, 
    4.711446e-14, 4.69332e-14, 4.730258e-14, 4.71872e-14, 4.747684e-14, 
    4.728461e-14, 4.751556e-14, 4.747134e-14, 4.760447e-14, 4.756636e-14, 
    4.773635e-14, 4.762207e-14, 4.782442e-14, 4.770909e-14, 4.772713e-14, 
    4.761828e-14, 4.696975e-14, 4.70919e-14, 4.69625e-14, 4.697993e-14, 
    4.697212e-14, 4.687692e-14, 4.682888e-14, 4.672834e-14, 4.674661e-14, 
    4.682047e-14, 4.698777e-14, 4.693103e-14, 4.707404e-14, 4.707081e-14, 
    4.722976e-14, 4.715812e-14, 4.742493e-14, 4.734918e-14, 4.756795e-14, 
    4.751297e-14, 4.756536e-14, 4.754948e-14, 4.756557e-14, 4.748492e-14, 
    4.751948e-14, 4.744851e-14, 4.717153e-14, 4.7253e-14, 4.700981e-14, 
    4.686324e-14, 4.676588e-14, 4.669671e-14, 4.670649e-14, 4.672513e-14, 
    4.68209e-14, 4.69109e-14, 4.697942e-14, 4.702523e-14, 4.707035e-14, 
    4.720668e-14, 4.727887e-14, 4.744022e-14, 4.741115e-14, 4.746041e-14, 
    4.75075e-14, 4.758646e-14, 4.757347e-14, 4.760823e-14, 4.745914e-14, 
    4.755824e-14, 4.739459e-14, 4.743937e-14, 4.708247e-14, 4.694635e-14, 
    4.688832e-14, 4.68376e-14, 4.671401e-14, 4.679937e-14, 4.676572e-14, 
    4.684578e-14, 4.689659e-14, 4.687147e-14, 4.702648e-14, 4.696624e-14, 
    4.728314e-14, 4.714676e-14, 4.750201e-14, 4.741712e-14, 4.752235e-14, 
    4.746868e-14, 4.756062e-14, 4.747788e-14, 4.762118e-14, 4.765234e-14, 
    4.763104e-14, 4.771286e-14, 4.747328e-14, 4.756535e-14, 4.687076e-14, 
    4.687485e-14, 4.689396e-14, 4.680996e-14, 4.680483e-14, 4.672784e-14, 
    4.679636e-14, 4.682551e-14, 4.689955e-14, 4.694329e-14, 4.698486e-14, 
    4.70762e-14, 4.71781e-14, 4.732046e-14, 4.742263e-14, 4.749105e-14, 
    4.744911e-14, 4.748613e-14, 4.744474e-14, 4.742533e-14, 4.764065e-14, 
    4.75198e-14, 4.77011e-14, 4.769108e-14, 4.760905e-14, 4.769221e-14, 
    4.687773e-14, 4.685415e-14, 4.677218e-14, 4.683633e-14, 4.671945e-14, 
    4.678487e-14, 4.682246e-14, 4.696747e-14, 4.699933e-14, 4.702882e-14, 
    4.708709e-14, 4.716179e-14, 4.729269e-14, 4.740647e-14, 4.751025e-14, 
    4.750265e-14, 4.750532e-14, 4.752848e-14, 4.747109e-14, 4.753789e-14, 
    4.754909e-14, 4.75198e-14, 4.768974e-14, 4.764122e-14, 4.769087e-14, 
    4.765928e-14, 4.686182e-14, 4.69015e-14, 4.688006e-14, 4.692037e-14, 
    4.689196e-14, 4.701819e-14, 4.7056e-14, 4.72328e-14, 4.716031e-14, 
    4.727568e-14, 4.717205e-14, 4.719041e-14, 4.727938e-14, 4.717766e-14, 
    4.740017e-14, 4.724932e-14, 4.752938e-14, 4.737887e-14, 4.75388e-14, 
    4.75098e-14, 4.755782e-14, 4.76008e-14, 4.765486e-14, 4.775449e-14, 
    4.773143e-14, 4.781472e-14, 4.696065e-14, 4.701205e-14, 4.700755e-14, 
    4.706134e-14, 4.71011e-14, 4.718725e-14, 4.732524e-14, 4.727338e-14, 
    4.736859e-14, 4.738769e-14, 4.724305e-14, 4.733185e-14, 4.704646e-14, 
    4.70926e-14, 4.706515e-14, 4.696469e-14, 4.72853e-14, 4.712087e-14, 
    4.742431e-14, 4.73354e-14, 4.759466e-14, 4.746578e-14, 4.771873e-14, 
    4.782659e-14, 4.792811e-14, 4.804647e-14, 4.704013e-14, 4.700521e-14, 
    4.706775e-14, 4.715416e-14, 4.723435e-14, 4.734082e-14, 4.735172e-14, 
    4.737164e-14, 4.742326e-14, 4.746663e-14, 4.737791e-14, 4.74775e-14, 
    4.710324e-14, 4.729957e-14, 4.699198e-14, 4.708466e-14, 4.714908e-14, 
    4.712085e-14, 4.726746e-14, 4.730197e-14, 4.744208e-14, 4.736969e-14, 
    4.779996e-14, 4.760983e-14, 4.813657e-14, 4.798965e-14, 4.699299e-14, 
    4.704002e-14, 4.720346e-14, 4.712573e-14, 4.734794e-14, 4.740254e-14, 
    4.744694e-14, 4.750361e-14, 4.750975e-14, 4.754331e-14, 4.74883e-14, 
    4.754115e-14, 4.734104e-14, 4.743052e-14, 4.718483e-14, 4.724467e-14, 
    4.721715e-14, 4.718694e-14, 4.728015e-14, 4.737931e-14, 4.738147e-14, 
    4.741323e-14, 4.750261e-14, 4.734884e-14, 4.782438e-14, 4.75309e-14, 
    4.709126e-14, 4.718167e-14, 4.719463e-14, 4.715962e-14, 4.739707e-14, 
    4.731109e-14, 4.75425e-14, 4.748002e-14, 4.758238e-14, 4.753152e-14, 
    4.752404e-14, 4.745869e-14, 4.741797e-14, 4.731503e-14, 4.72312e-14, 
    4.71647e-14, 4.718017e-14, 4.725321e-14, 4.738538e-14, 4.751028e-14, 
    4.748293e-14, 4.75746e-14, 4.733184e-14, 4.743369e-14, 4.739432e-14, 
    4.749694e-14, 4.727199e-14, 4.746345e-14, 4.722298e-14, 4.72441e-14, 
    4.730939e-14, 4.744056e-14, 4.746962e-14, 4.750057e-14, 4.748149e-14, 
    4.738874e-14, 4.737356e-14, 4.730781e-14, 4.728963e-14, 4.723951e-14, 
    4.719797e-14, 4.723591e-14, 4.727573e-14, 4.73888e-14, 4.749056e-14, 
    4.76014e-14, 4.762852e-14, 4.775772e-14, 4.76525e-14, 4.782601e-14, 
    4.767842e-14, 4.79338e-14, 4.74746e-14, 4.767417e-14, 4.731237e-14, 
    4.735142e-14, 4.742197e-14, 4.758368e-14, 4.749646e-14, 4.759848e-14, 
    4.737296e-14, 4.72557e-14, 4.72254e-14, 4.716874e-14, 4.722669e-14, 
    4.722198e-14, 4.72774e-14, 4.72596e-14, 4.739255e-14, 4.732116e-14, 
    4.752384e-14, 4.759768e-14, 4.780598e-14, 4.793341e-14, 4.806302e-14, 
    4.812016e-14, 4.813755e-14, 4.814481e-14 ;

 LITR1N_vr =
  5.557407e-05, 5.557386e-05, 5.55739e-05, 5.557373e-05, 5.557383e-05, 
    5.557372e-05, 5.557403e-05, 5.557385e-05, 5.557396e-05, 5.557405e-05, 
    5.557341e-05, 5.557372e-05, 5.557308e-05, 5.557328e-05, 5.557277e-05, 
    5.557311e-05, 5.557271e-05, 5.557279e-05, 5.557255e-05, 5.557262e-05, 
    5.557232e-05, 5.557252e-05, 5.557217e-05, 5.557237e-05, 5.557234e-05, 
    5.557253e-05, 5.557366e-05, 5.557345e-05, 5.557367e-05, 5.557364e-05, 
    5.557366e-05, 5.557382e-05, 5.557391e-05, 5.557408e-05, 5.557405e-05, 
    5.557392e-05, 5.557363e-05, 5.557373e-05, 5.557348e-05, 5.557348e-05, 
    5.557321e-05, 5.557333e-05, 5.557287e-05, 5.5573e-05, 5.557261e-05, 
    5.557271e-05, 5.557262e-05, 5.557265e-05, 5.557262e-05, 5.557276e-05, 
    5.55727e-05, 5.557283e-05, 5.557331e-05, 5.557317e-05, 5.557359e-05, 
    5.557385e-05, 5.557402e-05, 5.557414e-05, 5.557412e-05, 5.557409e-05, 
    5.557392e-05, 5.557376e-05, 5.557364e-05, 5.557356e-05, 5.557348e-05, 
    5.557325e-05, 5.557312e-05, 5.557284e-05, 5.557289e-05, 5.55728e-05, 
    5.557272e-05, 5.557258e-05, 5.557261e-05, 5.557255e-05, 5.557281e-05, 
    5.557263e-05, 5.557292e-05, 5.557284e-05, 5.557347e-05, 5.55737e-05, 
    5.55738e-05, 5.557389e-05, 5.557411e-05, 5.557396e-05, 5.557402e-05, 
    5.557388e-05, 5.557379e-05, 5.557383e-05, 5.557356e-05, 5.557367e-05, 
    5.557311e-05, 5.557335e-05, 5.557273e-05, 5.557288e-05, 5.557269e-05, 
    5.557279e-05, 5.557263e-05, 5.557277e-05, 5.557252e-05, 5.557247e-05, 
    5.557251e-05, 5.557236e-05, 5.557278e-05, 5.557262e-05, 5.557383e-05, 
    5.557383e-05, 5.557379e-05, 5.557394e-05, 5.557395e-05, 5.557408e-05, 
    5.557396e-05, 5.557391e-05, 5.557379e-05, 5.557371e-05, 5.557364e-05, 
    5.557348e-05, 5.55733e-05, 5.557305e-05, 5.557287e-05, 5.557275e-05, 
    5.557282e-05, 5.557276e-05, 5.557283e-05, 5.557287e-05, 5.557249e-05, 
    5.55727e-05, 5.557238e-05, 5.55724e-05, 5.557255e-05, 5.55724e-05, 
    5.557382e-05, 5.557386e-05, 5.557401e-05, 5.55739e-05, 5.55741e-05, 
    5.557399e-05, 5.557392e-05, 5.557367e-05, 5.557361e-05, 5.557356e-05, 
    5.557346e-05, 5.557333e-05, 5.55731e-05, 5.55729e-05, 5.557272e-05, 
    5.557273e-05, 5.557272e-05, 5.557268e-05, 5.557279e-05, 5.557267e-05, 
    5.557265e-05, 5.55727e-05, 5.55724e-05, 5.557249e-05, 5.55724e-05, 
    5.557245e-05, 5.557385e-05, 5.557378e-05, 5.557382e-05, 5.557375e-05, 
    5.55738e-05, 5.557358e-05, 5.557351e-05, 5.55732e-05, 5.557333e-05, 
    5.557313e-05, 5.557331e-05, 5.557328e-05, 5.557312e-05, 5.55733e-05, 
    5.557291e-05, 5.557317e-05, 5.557268e-05, 5.557295e-05, 5.557267e-05, 
    5.557272e-05, 5.557263e-05, 5.557256e-05, 5.557247e-05, 5.557229e-05, 
    5.557233e-05, 5.557219e-05, 5.557368e-05, 5.557359e-05, 5.55736e-05, 
    5.55735e-05, 5.557343e-05, 5.557328e-05, 5.557304e-05, 5.557313e-05, 
    5.557296e-05, 5.557293e-05, 5.557318e-05, 5.557303e-05, 5.557353e-05, 
    5.557345e-05, 5.55735e-05, 5.557367e-05, 5.557311e-05, 5.55734e-05, 
    5.557287e-05, 5.557302e-05, 5.557257e-05, 5.557279e-05, 5.557235e-05, 
    5.557216e-05, 5.557199e-05, 5.557178e-05, 5.557354e-05, 5.55736e-05, 
    5.557349e-05, 5.557334e-05, 5.55732e-05, 5.557301e-05, 5.557299e-05, 
    5.557296e-05, 5.557287e-05, 5.557279e-05, 5.557295e-05, 5.557277e-05, 
    5.557343e-05, 5.557308e-05, 5.557362e-05, 5.557346e-05, 5.557335e-05, 
    5.55734e-05, 5.557314e-05, 5.557308e-05, 5.557284e-05, 5.557296e-05, 
    5.557221e-05, 5.557254e-05, 5.557162e-05, 5.557188e-05, 5.557362e-05, 
    5.557354e-05, 5.557325e-05, 5.557339e-05, 5.5573e-05, 5.557291e-05, 
    5.557283e-05, 5.557273e-05, 5.557272e-05, 5.557266e-05, 5.557276e-05, 
    5.557266e-05, 5.557301e-05, 5.557285e-05, 5.557328e-05, 5.557318e-05, 
    5.557323e-05, 5.557328e-05, 5.557312e-05, 5.557295e-05, 5.557294e-05, 
    5.557289e-05, 5.557273e-05, 5.5573e-05, 5.557217e-05, 5.557268e-05, 
    5.557345e-05, 5.557329e-05, 5.557327e-05, 5.557333e-05, 5.557291e-05, 
    5.557307e-05, 5.557266e-05, 5.557277e-05, 5.557259e-05, 5.557268e-05, 
    5.557269e-05, 5.557281e-05, 5.557288e-05, 5.557306e-05, 5.55732e-05, 
    5.557332e-05, 5.557329e-05, 5.557317e-05, 5.557293e-05, 5.557272e-05, 
    5.557276e-05, 5.55726e-05, 5.557303e-05, 5.557285e-05, 5.557292e-05, 
    5.557274e-05, 5.557313e-05, 5.55728e-05, 5.557322e-05, 5.557318e-05, 
    5.557307e-05, 5.557284e-05, 5.557279e-05, 5.557273e-05, 5.557277e-05, 
    5.557293e-05, 5.557296e-05, 5.557307e-05, 5.55731e-05, 5.557319e-05, 
    5.557326e-05, 5.55732e-05, 5.557313e-05, 5.557293e-05, 5.557275e-05, 
    5.557256e-05, 5.557251e-05, 5.557228e-05, 5.557247e-05, 5.557216e-05, 
    5.557242e-05, 5.557198e-05, 5.557278e-05, 5.557243e-05, 5.557306e-05, 
    5.557299e-05, 5.557287e-05, 5.557259e-05, 5.557274e-05, 5.557256e-05, 
    5.557296e-05, 5.557316e-05, 5.557321e-05, 5.557331e-05, 5.557321e-05, 
    5.557322e-05, 5.557312e-05, 5.557316e-05, 5.557292e-05, 5.557305e-05, 
    5.557269e-05, 5.557256e-05, 5.55722e-05, 5.557198e-05, 5.557175e-05, 
    5.557165e-05, 5.557162e-05, 5.557161e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1_HR =
  8.09975e-13, 8.120347e-13, 8.116347e-13, 8.132943e-13, 8.123741e-13, 
    8.134603e-13, 8.10393e-13, 8.121162e-13, 8.110166e-13, 8.10161e-13, 
    8.165096e-13, 8.133683e-13, 8.197697e-13, 8.177702e-13, 8.227896e-13, 
    8.194583e-13, 8.234607e-13, 8.226944e-13, 8.250017e-13, 8.24341e-13, 
    8.272871e-13, 8.253065e-13, 8.288134e-13, 8.268147e-13, 8.271273e-13, 
    8.25241e-13, 8.140016e-13, 8.161185e-13, 8.13876e-13, 8.14178e-13, 
    8.140427e-13, 8.123929e-13, 8.115604e-13, 8.09818e-13, 8.101346e-13, 
    8.114145e-13, 8.143139e-13, 8.133307e-13, 8.15809e-13, 8.157531e-13, 
    8.185077e-13, 8.172662e-13, 8.218901e-13, 8.205773e-13, 8.243686e-13, 
    8.234159e-13, 8.243238e-13, 8.240486e-13, 8.243274e-13, 8.229298e-13, 
    8.235287e-13, 8.222987e-13, 8.174986e-13, 8.189105e-13, 8.146959e-13, 
    8.121558e-13, 8.104686e-13, 8.092698e-13, 8.094393e-13, 8.097623e-13, 
    8.11422e-13, 8.129817e-13, 8.141693e-13, 8.149631e-13, 8.15745e-13, 
    8.181078e-13, 8.193587e-13, 8.22155e-13, 8.216513e-13, 8.22505e-13, 
    8.233211e-13, 8.246894e-13, 8.244644e-13, 8.250667e-13, 8.22483e-13, 
    8.242004e-13, 8.213642e-13, 8.221404e-13, 8.159551e-13, 8.135961e-13, 
    8.125904e-13, 8.117115e-13, 8.095696e-13, 8.110488e-13, 8.104657e-13, 
    8.118531e-13, 8.127338e-13, 8.122984e-13, 8.149848e-13, 8.139408e-13, 
    8.194328e-13, 8.170693e-13, 8.232259e-13, 8.217548e-13, 8.235784e-13, 
    8.226483e-13, 8.242416e-13, 8.228076e-13, 8.252911e-13, 8.258311e-13, 
    8.25462e-13, 8.268801e-13, 8.227281e-13, 8.243235e-13, 8.122861e-13, 
    8.123571e-13, 8.126881e-13, 8.112324e-13, 8.111435e-13, 8.098092e-13, 
    8.109967e-13, 8.11502e-13, 8.127851e-13, 8.135431e-13, 8.142635e-13, 
    8.158466e-13, 8.176125e-13, 8.200796e-13, 8.218502e-13, 8.230359e-13, 
    8.223091e-13, 8.229508e-13, 8.222333e-13, 8.218971e-13, 8.256286e-13, 
    8.235341e-13, 8.266762e-13, 8.265026e-13, 8.25081e-13, 8.265222e-13, 
    8.12407e-13, 8.119983e-13, 8.105778e-13, 8.116895e-13, 8.096639e-13, 
    8.107977e-13, 8.114492e-13, 8.139621e-13, 8.145143e-13, 8.150255e-13, 
    8.160351e-13, 8.173298e-13, 8.195983e-13, 8.215702e-13, 8.233687e-13, 
    8.23237e-13, 8.232833e-13, 8.236845e-13, 8.226901e-13, 8.238478e-13, 
    8.240418e-13, 8.235342e-13, 8.264793e-13, 8.256385e-13, 8.264989e-13, 
    8.259516e-13, 8.121312e-13, 8.128189e-13, 8.124473e-13, 8.131459e-13, 
    8.126535e-13, 8.14841e-13, 8.154964e-13, 8.185603e-13, 8.173041e-13, 
    8.193036e-13, 8.175075e-13, 8.178258e-13, 8.193677e-13, 8.176048e-13, 
    8.214611e-13, 8.188467e-13, 8.237002e-13, 8.210918e-13, 8.238634e-13, 
    8.233609e-13, 8.241931e-13, 8.249379e-13, 8.258748e-13, 8.276014e-13, 
    8.272019e-13, 8.286452e-13, 8.138439e-13, 8.147348e-13, 8.146568e-13, 
    8.15589e-13, 8.16278e-13, 8.17771e-13, 8.201624e-13, 8.192637e-13, 
    8.209138e-13, 8.212447e-13, 8.187379e-13, 8.20277e-13, 8.153311e-13, 
    8.161306e-13, 8.15655e-13, 8.139139e-13, 8.194702e-13, 8.166206e-13, 
    8.218793e-13, 8.203385e-13, 8.248316e-13, 8.225981e-13, 8.269818e-13, 
    8.288509e-13, 8.306104e-13, 8.326615e-13, 8.152213e-13, 8.146161e-13, 
    8.157e-13, 8.171975e-13, 8.185873e-13, 8.204324e-13, 8.206213e-13, 
    8.209666e-13, 8.218612e-13, 8.226128e-13, 8.210753e-13, 8.228011e-13, 
    8.163151e-13, 8.197175e-13, 8.143869e-13, 8.159931e-13, 8.171095e-13, 
    8.166203e-13, 8.191611e-13, 8.197592e-13, 8.221874e-13, 8.209328e-13, 
    8.283894e-13, 8.250944e-13, 8.342231e-13, 8.31677e-13, 8.144045e-13, 
    8.152194e-13, 8.18052e-13, 8.167049e-13, 8.205558e-13, 8.215021e-13, 
    8.222715e-13, 8.232536e-13, 8.2336e-13, 8.239417e-13, 8.229883e-13, 
    8.239042e-13, 8.204363e-13, 8.21987e-13, 8.17729e-13, 8.187661e-13, 
    8.182892e-13, 8.177657e-13, 8.19381e-13, 8.210994e-13, 8.211368e-13, 
    8.216873e-13, 8.232363e-13, 8.205714e-13, 8.288128e-13, 8.237266e-13, 
    8.161075e-13, 8.176743e-13, 8.178989e-13, 8.172921e-13, 8.214072e-13, 
    8.199172e-13, 8.239276e-13, 8.228448e-13, 8.246187e-13, 8.237374e-13, 
    8.236077e-13, 8.224752e-13, 8.217695e-13, 8.199854e-13, 8.185327e-13, 
    8.173802e-13, 8.176483e-13, 8.189141e-13, 8.212046e-13, 8.233693e-13, 
    8.228952e-13, 8.24484e-13, 8.202768e-13, 8.220418e-13, 8.213596e-13, 
    8.231381e-13, 8.192396e-13, 8.225576e-13, 8.183902e-13, 8.187562e-13, 
    8.198876e-13, 8.22161e-13, 8.226646e-13, 8.232009e-13, 8.228702e-13, 
    8.212629e-13, 8.209997e-13, 8.198603e-13, 8.195452e-13, 8.186766e-13, 
    8.179568e-13, 8.186143e-13, 8.193043e-13, 8.212638e-13, 8.230274e-13, 
    8.249483e-13, 8.254184e-13, 8.276574e-13, 8.258339e-13, 8.288409e-13, 
    8.262832e-13, 8.30709e-13, 8.227508e-13, 8.262094e-13, 8.199393e-13, 
    8.206161e-13, 8.218388e-13, 8.246413e-13, 8.231297e-13, 8.248977e-13, 
    8.209895e-13, 8.189573e-13, 8.184321e-13, 8.174502e-13, 8.184546e-13, 
    8.183729e-13, 8.193334e-13, 8.190249e-13, 8.213289e-13, 8.200917e-13, 
    8.236042e-13, 8.24884e-13, 8.284937e-13, 8.307022e-13, 8.329484e-13, 
    8.339386e-13, 8.3424e-13, 8.343659e-13 ;

 LITR2C =
  1.939584e-05, 1.939582e-05, 1.939582e-05, 1.939581e-05, 1.939581e-05, 
    1.93958e-05, 1.939583e-05, 1.939582e-05, 1.939583e-05, 1.939583e-05, 
    1.939578e-05, 1.939581e-05, 1.939575e-05, 1.939576e-05, 1.939572e-05, 
    1.939575e-05, 1.939571e-05, 1.939572e-05, 1.93957e-05, 1.93957e-05, 
    1.939567e-05, 1.939569e-05, 1.939566e-05, 1.939568e-05, 1.939568e-05, 
    1.939569e-05, 1.93958e-05, 1.939578e-05, 1.93958e-05, 1.93958e-05, 
    1.93958e-05, 1.939581e-05, 1.939582e-05, 1.939584e-05, 1.939583e-05, 
    1.939582e-05, 1.93958e-05, 1.939581e-05, 1.939578e-05, 1.939578e-05, 
    1.939576e-05, 1.939577e-05, 1.939573e-05, 1.939574e-05, 1.93957e-05, 
    1.939571e-05, 1.93957e-05, 1.939571e-05, 1.93957e-05, 1.939572e-05, 
    1.939571e-05, 1.939572e-05, 1.939577e-05, 1.939575e-05, 1.939579e-05, 
    1.939582e-05, 1.939583e-05, 1.939584e-05, 1.939584e-05, 1.939584e-05, 
    1.939582e-05, 1.939581e-05, 1.93958e-05, 1.939579e-05, 1.939578e-05, 
    1.939576e-05, 1.939575e-05, 1.939572e-05, 1.939573e-05, 1.939572e-05, 
    1.939571e-05, 1.93957e-05, 1.93957e-05, 1.93957e-05, 1.939572e-05, 
    1.93957e-05, 1.939573e-05, 1.939572e-05, 1.939578e-05, 1.93958e-05, 
    1.939581e-05, 1.939582e-05, 1.939584e-05, 1.939583e-05, 1.939583e-05, 
    1.939582e-05, 1.939581e-05, 1.939581e-05, 1.939579e-05, 1.93958e-05, 
    1.939575e-05, 1.939577e-05, 1.939571e-05, 1.939573e-05, 1.939571e-05, 
    1.939572e-05, 1.93957e-05, 1.939572e-05, 1.939569e-05, 1.939569e-05, 
    1.939569e-05, 1.939568e-05, 1.939572e-05, 1.93957e-05, 1.939581e-05, 
    1.939581e-05, 1.939581e-05, 1.939583e-05, 1.939583e-05, 1.939584e-05, 
    1.939583e-05, 1.939582e-05, 1.939581e-05, 1.93958e-05, 1.93958e-05, 
    1.939578e-05, 1.939577e-05, 1.939574e-05, 1.939573e-05, 1.939571e-05, 
    1.939572e-05, 1.939572e-05, 1.939572e-05, 1.939573e-05, 1.939569e-05, 
    1.939571e-05, 1.939568e-05, 1.939568e-05, 1.93957e-05, 1.939568e-05, 
    1.939581e-05, 1.939582e-05, 1.939583e-05, 1.939582e-05, 1.939584e-05, 
    1.939583e-05, 1.939582e-05, 1.93958e-05, 1.939579e-05, 1.939579e-05, 
    1.939578e-05, 1.939577e-05, 1.939575e-05, 1.939573e-05, 1.939571e-05, 
    1.939571e-05, 1.939571e-05, 1.939571e-05, 1.939572e-05, 1.939571e-05, 
    1.939571e-05, 1.939571e-05, 1.939568e-05, 1.939569e-05, 1.939568e-05, 
    1.939569e-05, 1.939582e-05, 1.939581e-05, 1.939581e-05, 1.939581e-05, 
    1.939581e-05, 1.939579e-05, 1.939579e-05, 1.939576e-05, 1.939577e-05, 
    1.939575e-05, 1.939577e-05, 1.939576e-05, 1.939575e-05, 1.939577e-05, 
    1.939573e-05, 1.939575e-05, 1.939571e-05, 1.939573e-05, 1.939571e-05, 
    1.939571e-05, 1.93957e-05, 1.93957e-05, 1.939569e-05, 1.939567e-05, 
    1.939568e-05, 1.939566e-05, 1.93958e-05, 1.939579e-05, 1.939579e-05, 
    1.939578e-05, 1.939578e-05, 1.939576e-05, 1.939574e-05, 1.939575e-05, 
    1.939573e-05, 1.939573e-05, 1.939575e-05, 1.939574e-05, 1.939579e-05, 
    1.939578e-05, 1.939578e-05, 1.93958e-05, 1.939575e-05, 1.939577e-05, 
    1.939573e-05, 1.939574e-05, 1.93957e-05, 1.939572e-05, 1.939568e-05, 
    1.939566e-05, 1.939564e-05, 1.939563e-05, 1.939579e-05, 1.939579e-05, 
    1.939578e-05, 1.939577e-05, 1.939576e-05, 1.939574e-05, 1.939574e-05, 
    1.939573e-05, 1.939573e-05, 1.939572e-05, 1.939573e-05, 1.939572e-05, 
    1.939578e-05, 1.939575e-05, 1.939579e-05, 1.939578e-05, 1.939577e-05, 
    1.939577e-05, 1.939575e-05, 1.939575e-05, 1.939572e-05, 1.939573e-05, 
    1.939567e-05, 1.93957e-05, 1.939561e-05, 1.939563e-05, 1.939579e-05, 
    1.939579e-05, 1.939576e-05, 1.939577e-05, 1.939574e-05, 1.939573e-05, 
    1.939572e-05, 1.939571e-05, 1.939571e-05, 1.939571e-05, 1.939571e-05, 
    1.939571e-05, 1.939574e-05, 1.939573e-05, 1.939576e-05, 1.939575e-05, 
    1.939576e-05, 1.939576e-05, 1.939575e-05, 1.939573e-05, 1.939573e-05, 
    1.939573e-05, 1.939571e-05, 1.939574e-05, 1.939566e-05, 1.939571e-05, 
    1.939578e-05, 1.939577e-05, 1.939576e-05, 1.939577e-05, 1.939573e-05, 
    1.939574e-05, 1.939571e-05, 1.939572e-05, 1.93957e-05, 1.939571e-05, 
    1.939571e-05, 1.939572e-05, 1.939573e-05, 1.939574e-05, 1.939576e-05, 
    1.939577e-05, 1.939577e-05, 1.939575e-05, 1.939573e-05, 1.939571e-05, 
    1.939572e-05, 1.93957e-05, 1.939574e-05, 1.939572e-05, 1.939573e-05, 
    1.939571e-05, 1.939575e-05, 1.939572e-05, 1.939576e-05, 1.939575e-05, 
    1.939574e-05, 1.939572e-05, 1.939572e-05, 1.939571e-05, 1.939572e-05, 
    1.939573e-05, 1.939573e-05, 1.939574e-05, 1.939575e-05, 1.939575e-05, 
    1.939576e-05, 1.939576e-05, 1.939575e-05, 1.939573e-05, 1.939571e-05, 
    1.93957e-05, 1.939569e-05, 1.939567e-05, 1.939569e-05, 1.939566e-05, 
    1.939569e-05, 1.939564e-05, 1.939572e-05, 1.939569e-05, 1.939574e-05, 
    1.939574e-05, 1.939573e-05, 1.93957e-05, 1.939571e-05, 1.93957e-05, 
    1.939573e-05, 1.939575e-05, 1.939576e-05, 1.939577e-05, 1.939576e-05, 
    1.939576e-05, 1.939575e-05, 1.939575e-05, 1.939573e-05, 1.939574e-05, 
    1.939571e-05, 1.93957e-05, 1.939566e-05, 1.939564e-05, 1.939562e-05, 
    1.939561e-05, 1.939561e-05, 1.939561e-05 ;

 LITR2C_TO_SOIL1C =
  1.233469e-13, 1.236609e-13, 1.235999e-13, 1.238529e-13, 1.237126e-13, 
    1.238782e-13, 1.234106e-13, 1.236733e-13, 1.235057e-13, 1.233753e-13, 
    1.243431e-13, 1.238642e-13, 1.248401e-13, 1.245353e-13, 1.253005e-13, 
    1.247926e-13, 1.254028e-13, 1.252859e-13, 1.256377e-13, 1.25537e-13, 
    1.259861e-13, 1.256841e-13, 1.262188e-13, 1.259141e-13, 1.259617e-13, 
    1.256742e-13, 1.239607e-13, 1.242835e-13, 1.239416e-13, 1.239876e-13, 
    1.23967e-13, 1.237155e-13, 1.235886e-13, 1.23323e-13, 1.233712e-13, 
    1.235663e-13, 1.240083e-13, 1.238585e-13, 1.242363e-13, 1.242277e-13, 
    1.246477e-13, 1.244584e-13, 1.251633e-13, 1.249632e-13, 1.255412e-13, 
    1.253959e-13, 1.255343e-13, 1.254924e-13, 1.255349e-13, 1.253218e-13, 
    1.254131e-13, 1.252256e-13, 1.244939e-13, 1.247091e-13, 1.240666e-13, 
    1.236794e-13, 1.234221e-13, 1.232394e-13, 1.232652e-13, 1.233145e-13, 
    1.235675e-13, 1.238053e-13, 1.239863e-13, 1.241073e-13, 1.242265e-13, 
    1.245867e-13, 1.247774e-13, 1.252037e-13, 1.251269e-13, 1.252571e-13, 
    1.253815e-13, 1.255901e-13, 1.255558e-13, 1.256476e-13, 1.252537e-13, 
    1.255155e-13, 1.250832e-13, 1.252015e-13, 1.242585e-13, 1.238989e-13, 
    1.237456e-13, 1.236116e-13, 1.232851e-13, 1.235106e-13, 1.234217e-13, 
    1.236332e-13, 1.237675e-13, 1.237011e-13, 1.241106e-13, 1.239515e-13, 
    1.247887e-13, 1.244284e-13, 1.25367e-13, 1.251427e-13, 1.254207e-13, 
    1.252789e-13, 1.255218e-13, 1.253032e-13, 1.256818e-13, 1.257641e-13, 
    1.257079e-13, 1.259241e-13, 1.252911e-13, 1.255343e-13, 1.236992e-13, 
    1.2371e-13, 1.237605e-13, 1.235386e-13, 1.23525e-13, 1.233216e-13, 
    1.235026e-13, 1.235797e-13, 1.237753e-13, 1.238908e-13, 1.240007e-13, 
    1.24242e-13, 1.245112e-13, 1.248873e-13, 1.251572e-13, 1.25338e-13, 
    1.252272e-13, 1.25325e-13, 1.252156e-13, 1.251644e-13, 1.257333e-13, 
    1.254139e-13, 1.25893e-13, 1.258665e-13, 1.256498e-13, 1.258695e-13, 
    1.237176e-13, 1.236553e-13, 1.234388e-13, 1.236083e-13, 1.232995e-13, 
    1.234723e-13, 1.235716e-13, 1.239547e-13, 1.240389e-13, 1.241168e-13, 
    1.242707e-13, 1.244681e-13, 1.24814e-13, 1.251145e-13, 1.253887e-13, 
    1.253687e-13, 1.253757e-13, 1.254369e-13, 1.252853e-13, 1.254618e-13, 
    1.254913e-13, 1.25414e-13, 1.258629e-13, 1.257348e-13, 1.258659e-13, 
    1.257825e-13, 1.236756e-13, 1.237804e-13, 1.237238e-13, 1.238303e-13, 
    1.237552e-13, 1.240887e-13, 1.241886e-13, 1.246557e-13, 1.244642e-13, 
    1.24769e-13, 1.244952e-13, 1.245437e-13, 1.247788e-13, 1.2451e-13, 
    1.250979e-13, 1.246994e-13, 1.254393e-13, 1.250416e-13, 1.254641e-13, 
    1.253875e-13, 1.255144e-13, 1.25628e-13, 1.257708e-13, 1.26034e-13, 
    1.259731e-13, 1.261931e-13, 1.239367e-13, 1.240725e-13, 1.240606e-13, 
    1.242027e-13, 1.243078e-13, 1.245354e-13, 1.248999e-13, 1.247629e-13, 
    1.250145e-13, 1.250649e-13, 1.246828e-13, 1.249174e-13, 1.241634e-13, 
    1.242853e-13, 1.242128e-13, 1.239474e-13, 1.247944e-13, 1.2436e-13, 
    1.251617e-13, 1.249268e-13, 1.256118e-13, 1.252713e-13, 1.259395e-13, 
    1.262245e-13, 1.264927e-13, 1.268054e-13, 1.241467e-13, 1.240544e-13, 
    1.242196e-13, 1.24448e-13, 1.246598e-13, 1.249411e-13, 1.249699e-13, 
    1.250225e-13, 1.251589e-13, 1.252735e-13, 1.250391e-13, 1.253022e-13, 
    1.243134e-13, 1.248321e-13, 1.240195e-13, 1.242643e-13, 1.244345e-13, 
    1.2436e-13, 1.247473e-13, 1.248385e-13, 1.252086e-13, 1.250174e-13, 
    1.261541e-13, 1.256518e-13, 1.270435e-13, 1.266553e-13, 1.240222e-13, 
    1.241464e-13, 1.245782e-13, 1.243728e-13, 1.249599e-13, 1.251042e-13, 
    1.252215e-13, 1.253712e-13, 1.253874e-13, 1.254761e-13, 1.253307e-13, 
    1.254704e-13, 1.249417e-13, 1.251781e-13, 1.24529e-13, 1.246871e-13, 
    1.246144e-13, 1.245346e-13, 1.247808e-13, 1.250428e-13, 1.250485e-13, 
    1.251324e-13, 1.253685e-13, 1.249623e-13, 1.262187e-13, 1.254433e-13, 
    1.242818e-13, 1.245206e-13, 1.245549e-13, 1.244624e-13, 1.250897e-13, 
    1.248625e-13, 1.254739e-13, 1.253089e-13, 1.255793e-13, 1.254449e-13, 
    1.254252e-13, 1.252525e-13, 1.251449e-13, 1.24873e-13, 1.246515e-13, 
    1.244758e-13, 1.245167e-13, 1.247096e-13, 1.250588e-13, 1.253888e-13, 
    1.253165e-13, 1.255588e-13, 1.249174e-13, 1.251865e-13, 1.250825e-13, 
    1.253536e-13, 1.247593e-13, 1.252651e-13, 1.246298e-13, 1.246856e-13, 
    1.248581e-13, 1.252046e-13, 1.252814e-13, 1.253632e-13, 1.253127e-13, 
    1.250677e-13, 1.250276e-13, 1.248539e-13, 1.248058e-13, 1.246734e-13, 
    1.245637e-13, 1.246639e-13, 1.247691e-13, 1.250679e-13, 1.253367e-13, 
    1.256296e-13, 1.257012e-13, 1.260426e-13, 1.257646e-13, 1.26223e-13, 
    1.25833e-13, 1.265078e-13, 1.252945e-13, 1.258218e-13, 1.248659e-13, 
    1.249691e-13, 1.251555e-13, 1.255827e-13, 1.253523e-13, 1.256218e-13, 
    1.25026e-13, 1.247162e-13, 1.246362e-13, 1.244865e-13, 1.246396e-13, 
    1.246271e-13, 1.247736e-13, 1.247265e-13, 1.250778e-13, 1.248892e-13, 
    1.254246e-13, 1.256197e-13, 1.2617e-13, 1.265067e-13, 1.268492e-13, 
    1.270001e-13, 1.270461e-13, 1.270653e-13 ;

 LITR2C_vr =
  0.001107522, 0.001107521, 0.001107521, 0.001107521, 0.001107521, 
    0.00110752, 0.001107522, 0.001107521, 0.001107522, 0.001107522, 
    0.001107519, 0.001107521, 0.001107517, 0.001107518, 0.001107516, 
    0.001107517, 0.001107515, 0.001107516, 0.001107514, 0.001107515, 
    0.001107513, 0.001107514, 0.001107512, 0.001107513, 0.001107513, 
    0.001107514, 0.00110752, 0.001107519, 0.00110752, 0.00110752, 0.00110752, 
    0.001107521, 0.001107521, 0.001107522, 0.001107522, 0.001107522, 
    0.00110752, 0.001107521, 0.001107519, 0.001107519, 0.001107518, 
    0.001107518, 0.001107516, 0.001107517, 0.001107515, 0.001107515, 
    0.001107515, 0.001107515, 0.001107515, 0.001107515, 0.001107515, 
    0.001107516, 0.001107518, 0.001107518, 0.00110752, 0.001107521, 
    0.001107522, 0.001107523, 0.001107523, 0.001107522, 0.001107522, 
    0.001107521, 0.00110752, 0.00110752, 0.001107519, 0.001107518, 
    0.001107517, 0.001107516, 0.001107516, 0.001107516, 0.001107515, 
    0.001107514, 0.001107515, 0.001107514, 0.001107516, 0.001107515, 
    0.001107516, 0.001107516, 0.001107519, 0.00110752, 0.001107521, 
    0.001107521, 0.001107523, 0.001107522, 0.001107522, 0.001107521, 
    0.001107521, 0.001107521, 0.00110752, 0.00110752, 0.001107517, 
    0.001107519, 0.001107515, 0.001107516, 0.001107515, 0.001107516, 
    0.001107515, 0.001107516, 0.001107514, 0.001107514, 0.001107514, 
    0.001107513, 0.001107516, 0.001107515, 0.001107521, 0.001107521, 
    0.001107521, 0.001107522, 0.001107522, 0.001107522, 0.001107522, 
    0.001107521, 0.001107521, 0.00110752, 0.00110752, 0.001107519, 
    0.001107518, 0.001107517, 0.001107516, 0.001107515, 0.001107516, 
    0.001107515, 0.001107516, 0.001107516, 0.001107514, 0.001107515, 
    0.001107513, 0.001107514, 0.001107514, 0.001107514, 0.001107521, 
    0.001107521, 0.001107522, 0.001107521, 0.001107523, 0.001107522, 
    0.001107522, 0.00110752, 0.00110752, 0.00110752, 0.001107519, 
    0.001107518, 0.001107517, 0.001107516, 0.001107515, 0.001107515, 
    0.001107515, 0.001107515, 0.001107516, 0.001107515, 0.001107515, 
    0.001107515, 0.001107514, 0.001107514, 0.001107514, 0.001107514, 
    0.001107521, 0.001107521, 0.001107521, 0.001107521, 0.001107521, 
    0.00110752, 0.001107519, 0.001107518, 0.001107518, 0.001107517, 
    0.001107518, 0.001107518, 0.001107517, 0.001107518, 0.001107516, 
    0.001107518, 0.001107515, 0.001107516, 0.001107515, 0.001107515, 
    0.001107515, 0.001107514, 0.001107514, 0.001107513, 0.001107513, 
    0.001107512, 0.00110752, 0.00110752, 0.00110752, 0.001107519, 
    0.001107519, 0.001107518, 0.001107517, 0.001107517, 0.001107516, 
    0.001107516, 0.001107518, 0.001107517, 0.001107519, 0.001107519, 
    0.001107519, 0.00110752, 0.001107517, 0.001107519, 0.001107516, 
    0.001107517, 0.001107514, 0.001107516, 0.001107513, 0.001107512, 
    0.001107511, 0.00110751, 0.001107519, 0.00110752, 0.001107519, 
    0.001107518, 0.001107518, 0.001107517, 0.001107517, 0.001107516, 
    0.001107516, 0.001107516, 0.001107516, 0.001107516, 0.001107519, 
    0.001107517, 0.00110752, 0.001107519, 0.001107519, 0.001107519, 
    0.001107517, 0.001107517, 0.001107516, 0.001107516, 0.001107513, 
    0.001107514, 0.001107509, 0.001107511, 0.00110752, 0.001107519, 
    0.001107518, 0.001107519, 0.001107517, 0.001107516, 0.001107516, 
    0.001107515, 0.001107515, 0.001107515, 0.001107515, 0.001107515, 
    0.001107517, 0.001107516, 0.001107518, 0.001107518, 0.001107518, 
    0.001107518, 0.001107517, 0.001107516, 0.001107516, 0.001107516, 
    0.001107515, 0.001107517, 0.001107512, 0.001107515, 0.001107519, 
    0.001107518, 0.001107518, 0.001107518, 0.001107516, 0.001107517, 
    0.001107515, 0.001107516, 0.001107514, 0.001107515, 0.001107515, 
    0.001107516, 0.001107516, 0.001107517, 0.001107518, 0.001107518, 
    0.001107518, 0.001107518, 0.001107516, 0.001107515, 0.001107515, 
    0.001107515, 0.001107517, 0.001107516, 0.001107516, 0.001107515, 
    0.001107517, 0.001107516, 0.001107518, 0.001107518, 0.001107517, 
    0.001107516, 0.001107516, 0.001107515, 0.001107515, 0.001107516, 
    0.001107516, 0.001107517, 0.001107517, 0.001107518, 0.001107518, 
    0.001107518, 0.001107517, 0.001107516, 0.001107515, 0.001107514, 
    0.001107514, 0.001107513, 0.001107514, 0.001107512, 0.001107514, 
    0.001107511, 0.001107516, 0.001107514, 0.001107517, 0.001107517, 
    0.001107516, 0.001107514, 0.001107515, 0.001107514, 0.001107516, 
    0.001107518, 0.001107518, 0.001107518, 0.001107518, 0.001107518, 
    0.001107517, 0.001107518, 0.001107516, 0.001107517, 0.001107515, 
    0.001107514, 0.001107513, 0.001107511, 0.00110751, 0.00110751, 
    0.001107509, 0.001107509,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N =
  2.684241e-07, 2.684239e-07, 2.684239e-07, 2.684237e-07, 2.684238e-07, 
    2.684237e-07, 2.684241e-07, 2.684238e-07, 2.68424e-07, 2.684241e-07, 
    2.684233e-07, 2.684237e-07, 2.684228e-07, 2.684231e-07, 2.684225e-07, 
    2.684229e-07, 2.684224e-07, 2.684225e-07, 2.684222e-07, 2.684223e-07, 
    2.684219e-07, 2.684221e-07, 2.684217e-07, 2.684219e-07, 2.684219e-07, 
    2.684222e-07, 2.684236e-07, 2.684233e-07, 2.684236e-07, 2.684236e-07, 
    2.684236e-07, 2.684238e-07, 2.684239e-07, 2.684241e-07, 2.684241e-07, 
    2.684239e-07, 2.684235e-07, 2.684237e-07, 2.684233e-07, 2.684234e-07, 
    2.68423e-07, 2.684232e-07, 2.684226e-07, 2.684228e-07, 2.684223e-07, 
    2.684224e-07, 2.684223e-07, 2.684223e-07, 2.684223e-07, 2.684224e-07, 
    2.684224e-07, 2.684225e-07, 2.684232e-07, 2.68423e-07, 2.684235e-07, 
    2.684238e-07, 2.684241e-07, 2.684242e-07, 2.684242e-07, 2.684241e-07, 
    2.684239e-07, 2.684237e-07, 2.684236e-07, 2.684235e-07, 2.684234e-07, 
    2.684231e-07, 2.684229e-07, 2.684226e-07, 2.684226e-07, 2.684225e-07, 
    2.684224e-07, 2.684222e-07, 2.684222e-07, 2.684222e-07, 2.684225e-07, 
    2.684223e-07, 2.684226e-07, 2.684226e-07, 2.684233e-07, 2.684237e-07, 
    2.684238e-07, 2.684239e-07, 2.684242e-07, 2.68424e-07, 2.684241e-07, 
    2.684239e-07, 2.684237e-07, 2.684238e-07, 2.684235e-07, 2.684236e-07, 
    2.684229e-07, 2.684232e-07, 2.684224e-07, 2.684226e-07, 2.684224e-07, 
    2.684225e-07, 2.684223e-07, 2.684225e-07, 2.684221e-07, 2.684221e-07, 
    2.684221e-07, 2.684219e-07, 2.684225e-07, 2.684223e-07, 2.684238e-07, 
    2.684238e-07, 2.684238e-07, 2.684239e-07, 2.68424e-07, 2.684241e-07, 
    2.68424e-07, 2.684239e-07, 2.684237e-07, 2.684237e-07, 2.684235e-07, 
    2.684233e-07, 2.684231e-07, 2.684228e-07, 2.684226e-07, 2.684224e-07, 
    2.684225e-07, 2.684224e-07, 2.684225e-07, 2.684226e-07, 2.684221e-07, 
    2.684224e-07, 2.68422e-07, 2.68422e-07, 2.684222e-07, 2.68422e-07, 
    2.684238e-07, 2.684239e-07, 2.68424e-07, 2.684239e-07, 2.684241e-07, 
    2.68424e-07, 2.684239e-07, 2.684236e-07, 2.684235e-07, 2.684235e-07, 
    2.684233e-07, 2.684232e-07, 2.684229e-07, 2.684226e-07, 2.684224e-07, 
    2.684224e-07, 2.684224e-07, 2.684224e-07, 2.684225e-07, 2.684223e-07, 
    2.684223e-07, 2.684224e-07, 2.68422e-07, 2.684221e-07, 2.68422e-07, 
    2.68422e-07, 2.684238e-07, 2.684237e-07, 2.684238e-07, 2.684237e-07, 
    2.684238e-07, 2.684235e-07, 2.684234e-07, 2.68423e-07, 2.684232e-07, 
    2.684229e-07, 2.684232e-07, 2.684231e-07, 2.684229e-07, 2.684231e-07, 
    2.684226e-07, 2.68423e-07, 2.684224e-07, 2.684227e-07, 2.684223e-07, 
    2.684224e-07, 2.684223e-07, 2.684222e-07, 2.684221e-07, 2.684218e-07, 
    2.684219e-07, 2.684217e-07, 2.684236e-07, 2.684235e-07, 2.684235e-07, 
    2.684234e-07, 2.684233e-07, 2.684231e-07, 2.684228e-07, 2.684229e-07, 
    2.684227e-07, 2.684227e-07, 2.68423e-07, 2.684228e-07, 2.684234e-07, 
    2.684233e-07, 2.684234e-07, 2.684236e-07, 2.684229e-07, 2.684233e-07, 
    2.684226e-07, 2.684228e-07, 2.684222e-07, 2.684225e-07, 2.684219e-07, 
    2.684217e-07, 2.684214e-07, 2.684212e-07, 2.684234e-07, 2.684235e-07, 
    2.684234e-07, 2.684232e-07, 2.68423e-07, 2.684228e-07, 2.684228e-07, 
    2.684227e-07, 2.684226e-07, 2.684225e-07, 2.684227e-07, 2.684225e-07, 
    2.684233e-07, 2.684229e-07, 2.684235e-07, 2.684233e-07, 2.684232e-07, 
    2.684233e-07, 2.684229e-07, 2.684229e-07, 2.684225e-07, 2.684227e-07, 
    2.684217e-07, 2.684222e-07, 2.68421e-07, 2.684213e-07, 2.684235e-07, 
    2.684234e-07, 2.684231e-07, 2.684232e-07, 2.684228e-07, 2.684226e-07, 
    2.684225e-07, 2.684224e-07, 2.684224e-07, 2.684223e-07, 2.684224e-07, 
    2.684223e-07, 2.684228e-07, 2.684226e-07, 2.684231e-07, 2.68423e-07, 
    2.68423e-07, 2.684231e-07, 2.684229e-07, 2.684227e-07, 2.684227e-07, 
    2.684226e-07, 2.684224e-07, 2.684228e-07, 2.684217e-07, 2.684224e-07, 
    2.684233e-07, 2.684231e-07, 2.684231e-07, 2.684232e-07, 2.684226e-07, 
    2.684228e-07, 2.684223e-07, 2.684225e-07, 2.684222e-07, 2.684223e-07, 
    2.684224e-07, 2.684225e-07, 2.684226e-07, 2.684228e-07, 2.68423e-07, 
    2.684232e-07, 2.684231e-07, 2.68423e-07, 2.684227e-07, 2.684224e-07, 
    2.684224e-07, 2.684222e-07, 2.684228e-07, 2.684226e-07, 2.684226e-07, 
    2.684224e-07, 2.684229e-07, 2.684225e-07, 2.68423e-07, 2.68423e-07, 
    2.684228e-07, 2.684226e-07, 2.684225e-07, 2.684224e-07, 2.684224e-07, 
    2.684227e-07, 2.684227e-07, 2.684228e-07, 2.684229e-07, 2.68423e-07, 
    2.684231e-07, 2.68423e-07, 2.684229e-07, 2.684227e-07, 2.684224e-07, 
    2.684222e-07, 2.684221e-07, 2.684218e-07, 2.684221e-07, 2.684217e-07, 
    2.68422e-07, 2.684214e-07, 2.684225e-07, 2.68422e-07, 2.684228e-07, 
    2.684228e-07, 2.684226e-07, 2.684222e-07, 2.684224e-07, 2.684222e-07, 
    2.684227e-07, 2.68423e-07, 2.68423e-07, 2.684232e-07, 2.68423e-07, 
    2.68423e-07, 2.684229e-07, 2.68423e-07, 2.684226e-07, 2.684228e-07, 
    2.684224e-07, 2.684222e-07, 2.684217e-07, 2.684214e-07, 2.684212e-07, 
    2.68421e-07, 2.68421e-07, 2.68421e-07 ;

 LITR2N_TNDNCY_VERT_TRANS =
  -6.862535e-26, 9.803622e-27, 9.803622e-26, 1.102908e-25, 7.842898e-26, 
    -2.745014e-25, 1.225453e-25, 1.151926e-25, -3.676358e-26, 2.695996e-26, 
    -3.504795e-25, -2.695996e-26, -1.225453e-26, -9.803622e-26, 
    -1.715634e-26, 4.901811e-26, -1.102908e-25, 2.450906e-25, 2.475414e-25, 
    1.887197e-25, -5.146902e-26, 4.901811e-26, 1.078398e-25, -2.450905e-26, 
    -3.676358e-26, -9.068351e-26, 2.205815e-25, 9.803622e-26, 3.186177e-26, 
    -7.842898e-26, 6.862535e-26, 4.901811e-27, 1.127417e-25, 1.053889e-25, 
    -2.695996e-26, -3.063632e-25, -1.54407e-25, -9.803622e-27, -4.901811e-26, 
    -1.519561e-25, 3.921449e-26, 8.578169e-26, 9.803622e-26, 1.81367e-25, 
    4.166539e-26, -9.803622e-26, 1.470543e-26, 1.960724e-25, -1.102908e-25, 
    2.941087e-26, 2.205815e-26, 2.32836e-25, -1.102908e-25, -3.921449e-26, 
    5.637083e-26, -1.56858e-25, -2.769523e-25, -5.882173e-26, 5.637083e-26, 
    -1.519561e-25, -1.176435e-25, 2.695996e-26, 4.901811e-27, -3.431268e-26, 
    -1.151926e-25, 2.450906e-27, 1.225453e-25, 5.882173e-26, -4.41163e-26, 
    -5.882173e-26, -8.578169e-26, 7.597807e-26, 3.676358e-26, 1.127417e-25, 
    2.156797e-25, 2.205815e-26, 1.078398e-25, 9.803622e-26, -2.034252e-25, 
    -5.882173e-26, -1.495052e-25, 1.127417e-25, 1.54407e-25, 1.81367e-25, 
    -2.303851e-25, 8.087988e-26, -1.470543e-26, -5.882173e-26, 1.936215e-25, 
    2.205815e-26, -3.847922e-25, -1.960724e-25, 8.578169e-26, -1.642107e-25, 
    -2.867559e-25, -1.960724e-26, 9.558531e-26, -1.617598e-25, 2.941087e-26, 
    -1.372507e-25, -2.59796e-25, -1.715634e-25, 2.695996e-26, 1.617598e-25, 
    -1.004871e-25, -1.004871e-25, -1.936215e-25, 9.803622e-26, -1.053889e-25, 
    1.838179e-25, -1.495052e-25, 9.068351e-26, 3.921449e-26, 1.740143e-25, 
    2.058761e-25, 2.941087e-26, 1.29898e-25, -5.146902e-26, -2.450906e-27, 
    3.284213e-25, 8.087988e-26, -7.597807e-26, 5.637083e-26, -4.901811e-27, 
    1.887197e-25, -1.078398e-25, 9.803622e-26, 4.65672e-26, -1.81367e-25, 
    5.146902e-26, 6.617445e-26, 9.803622e-27, -1.470543e-25, -2.205815e-26, 
    -2.450906e-27, 1.102908e-25, 9.803622e-26, -1.985233e-25, 2.941087e-26, 
    6.862535e-26, -4.65672e-26, 5.882173e-26, -5.146902e-26, -8.578169e-26, 
    2.59796e-25, -2.205815e-26, 7.842898e-26, -1.102908e-25, -1.151926e-25, 
    7.352717e-27, -1.127417e-25, -2.695996e-26, -3.676358e-26, -6.127264e-26, 
    -4.166539e-26, 1.838179e-25, 1.274471e-25, 3.186177e-26, 5.146902e-26, 
    3.431268e-26, -1.495052e-25, -7.352717e-26, -2.107779e-25, -1.715634e-26, 
    -2.08327e-25, 4.65672e-26, -1.078398e-25, 1.715634e-26, -9.803622e-27, 
    2.377378e-25, 8.333079e-26, -5.882173e-26, 1.691125e-25, 2.59796e-25, 
    -1.151926e-25, 9.558531e-26, 1.495052e-25, -1.715634e-26, -1.102908e-25, 
    -1.127417e-25, 1.960724e-26, -4.901811e-26, 2.377378e-25, -5.391992e-26, 
    4.65672e-26, -2.132288e-25, 7.352717e-27, -1.225453e-26, 1.666616e-25, 
    3.186177e-26, -1.960724e-26, -1.078398e-25, 2.941087e-26, 6.372354e-26, 
    -1.960724e-26, 2.205815e-26, 1.200944e-25, -1.249962e-25, 2.058761e-25, 
    -7.352717e-27, -1.789161e-25, 1.715634e-25, -7.352717e-27, 7.597807e-26, 
    1.225453e-26, -7.352717e-27, 3.039123e-25, -1.715634e-26, -1.862688e-25, 
    1.470543e-26, 1.078398e-25, 1.715634e-25, -1.715634e-25, 5.882173e-26, 
    -2.058761e-25, 1.715634e-26, 8.82326e-26, 2.32836e-25, 3.186177e-26, 
    1.02938e-25, 2.646978e-25, 8.578169e-26, 2.034252e-25, 3.259704e-25, 
    -1.249962e-25, 7.352717e-27, -1.02938e-25, 1.102908e-25, 2.450906e-27, 
    3.921449e-26, 7.352717e-26, -1.470543e-25, 5.882173e-26, 1.004871e-25, 
    -1.02938e-25, -2.59796e-25, 8.333079e-26, -8.333079e-26, -4.901811e-27, 
    5.882173e-26, 1.102908e-25, 1.078398e-25, -4.901811e-27, -8.333079e-26, 
    0, 3.872431e-25, -7.352717e-26, 9.313441e-26, -2.401887e-25, 
    6.862535e-26, -1.078398e-25, -2.450905e-26, 5.637083e-26, 2.769523e-25, 
    1.004871e-25, -2.450906e-27, -1.004871e-25, -1.715634e-26, -1.715634e-26, 
    4.901811e-27, -2.205815e-26, -1.127417e-25, -9.803622e-26, 1.078398e-25, 
    -9.803622e-27, 8.333079e-26, -1.54407e-25, 1.789161e-25, -7.842898e-26, 
    -2.450905e-26, -9.803622e-26, -1.225453e-25, -5.391992e-26, 1.323489e-25, 
    -1.81367e-25, -1.911706e-25, -2.695996e-26, 7.842898e-26, -1.642107e-25, 
    -1.225453e-25, -4.901811e-27, -1.225453e-25, 1.740143e-25, 1.740143e-25, 
    -1.102908e-25, -6.617445e-26, -1.397016e-25, 1.078398e-25, 2.205815e-26, 
    -1.176435e-25, 1.911706e-25, 1.740143e-25, 1.764652e-25, -4.901811e-27, 
    9.313441e-26, -2.230324e-25, -4.166539e-26, 1.225453e-25, 4.65672e-26, 
    2.009742e-25, -7.842898e-26, 8.333079e-26, -2.426396e-25, 9.558531e-26, 
    -4.65672e-26, -1.838179e-25, -2.671487e-25, -1.911706e-25, -7.842898e-26, 
    4.901811e-26, -9.803622e-26, -1.225453e-26, -1.56858e-25, -6.372354e-26, 
    1.102908e-25, 2.034252e-25, 5.637083e-26, -1.02938e-25, -1.02938e-25, 
    1.02938e-25, -4.65672e-26, -5.637083e-26, 1.274471e-25, -1.372507e-25, 
    -3.676358e-26, 2.450905e-26, -2.254833e-25, 3.676358e-26, 2.794032e-25, 
    -4.65672e-26, 2.32836e-25, -2.303851e-25, 1.004871e-25, -9.558531e-26, 
    -1.887197e-25, -9.803622e-27, -1.249962e-25, 8.578169e-26,
  2.676227e-32, 2.676224e-32, 2.676225e-32, 2.676223e-32, 2.676224e-32, 
    2.676223e-32, 2.676227e-32, 2.676224e-32, 2.676226e-32, 2.676227e-32, 
    2.676219e-32, 2.676223e-32, 2.676214e-32, 2.676217e-32, 2.676211e-32, 
    2.676215e-32, 2.67621e-32, 2.676211e-32, 2.676208e-32, 2.676209e-32, 
    2.676205e-32, 2.676207e-32, 2.676203e-32, 2.676205e-32, 2.676205e-32, 
    2.676207e-32, 2.676222e-32, 2.676219e-32, 2.676222e-32, 2.676222e-32, 
    2.676222e-32, 2.676224e-32, 2.676225e-32, 2.676227e-32, 2.676227e-32, 
    2.676225e-32, 2.676222e-32, 2.676223e-32, 2.67622e-32, 2.67622e-32, 
    2.676216e-32, 2.676218e-32, 2.676212e-32, 2.676214e-32, 2.676209e-32, 
    2.67621e-32, 2.676209e-32, 2.676209e-32, 2.676209e-32, 2.67621e-32, 
    2.67621e-32, 2.676211e-32, 2.676217e-32, 2.676216e-32, 2.676221e-32, 
    2.676224e-32, 2.676227e-32, 2.676228e-32, 2.676228e-32, 2.676227e-32, 
    2.676225e-32, 2.676223e-32, 2.676222e-32, 2.676221e-32, 2.67622e-32, 
    2.676217e-32, 2.676215e-32, 2.676212e-32, 2.676212e-32, 2.676211e-32, 
    2.67621e-32, 2.676208e-32, 2.676209e-32, 2.676208e-32, 2.676211e-32, 
    2.676209e-32, 2.676212e-32, 2.676212e-32, 2.676219e-32, 2.676222e-32, 
    2.676224e-32, 2.676225e-32, 2.676228e-32, 2.676226e-32, 2.676227e-32, 
    2.676225e-32, 2.676224e-32, 2.676224e-32, 2.676221e-32, 2.676222e-32, 
    2.676215e-32, 2.676218e-32, 2.67621e-32, 2.676212e-32, 2.676209e-32, 
    2.676211e-32, 2.676209e-32, 2.676211e-32, 2.676207e-32, 2.676207e-32, 
    2.676207e-32, 2.676205e-32, 2.676211e-32, 2.676209e-32, 2.676224e-32, 
    2.676224e-32, 2.676224e-32, 2.676226e-32, 2.676226e-32, 2.676227e-32, 
    2.676226e-32, 2.676225e-32, 2.676224e-32, 2.676223e-32, 2.676222e-32, 
    2.67622e-32, 2.676217e-32, 2.676214e-32, 2.676212e-32, 2.67621e-32, 
    2.676211e-32, 2.67621e-32, 2.676211e-32, 2.676212e-32, 2.676207e-32, 
    2.67621e-32, 2.676206e-32, 2.676206e-32, 2.676208e-32, 2.676206e-32, 
    2.676224e-32, 2.676225e-32, 2.676227e-32, 2.676225e-32, 2.676228e-32, 
    2.676226e-32, 2.676225e-32, 2.676222e-32, 2.676221e-32, 2.676221e-32, 
    2.676219e-32, 2.676218e-32, 2.676215e-32, 2.676212e-32, 2.67621e-32, 
    2.67621e-32, 2.67621e-32, 2.676209e-32, 2.676211e-32, 2.676209e-32, 
    2.676209e-32, 2.67621e-32, 2.676206e-32, 2.676207e-32, 2.676206e-32, 
    2.676207e-32, 2.676224e-32, 2.676224e-32, 2.676224e-32, 2.676223e-32, 
    2.676224e-32, 2.676221e-32, 2.67622e-32, 2.676216e-32, 2.676218e-32, 
    2.676215e-32, 2.676217e-32, 2.676217e-32, 2.676215e-32, 2.676217e-32, 
    2.676212e-32, 2.676216e-32, 2.676209e-32, 2.676213e-32, 2.676209e-32, 
    2.67621e-32, 2.676209e-32, 2.676208e-32, 2.676207e-32, 2.676204e-32, 
    2.676205e-32, 2.676203e-32, 2.676222e-32, 2.676221e-32, 2.676221e-32, 
    2.67622e-32, 2.676219e-32, 2.676217e-32, 2.676214e-32, 2.676215e-32, 
    2.676213e-32, 2.676213e-32, 2.676216e-32, 2.676214e-32, 2.67622e-32, 
    2.676219e-32, 2.67622e-32, 2.676222e-32, 2.676215e-32, 2.676219e-32, 
    2.676212e-32, 2.676214e-32, 2.676208e-32, 2.676211e-32, 2.676205e-32, 
    2.676203e-32, 2.6762e-32, 2.676198e-32, 2.67622e-32, 2.676221e-32, 
    2.67622e-32, 2.676218e-32, 2.676216e-32, 2.676214e-32, 2.676213e-32, 
    2.676213e-32, 2.676212e-32, 2.676211e-32, 2.676213e-32, 2.676211e-32, 
    2.676219e-32, 2.676214e-32, 2.676222e-32, 2.676219e-32, 2.676218e-32, 
    2.676219e-32, 2.676215e-32, 2.676214e-32, 2.676212e-32, 2.676213e-32, 
    2.676203e-32, 2.676208e-32, 2.676196e-32, 2.676199e-32, 2.676222e-32, 
    2.67622e-32, 2.676217e-32, 2.676219e-32, 2.676214e-32, 2.676212e-32, 
    2.676211e-32, 2.67621e-32, 2.67621e-32, 2.676209e-32, 2.67621e-32, 
    2.676209e-32, 2.676214e-32, 2.676212e-32, 2.676217e-32, 2.676216e-32, 
    2.676217e-32, 2.676217e-32, 2.676215e-32, 2.676213e-32, 2.676213e-32, 
    2.676212e-32, 2.67621e-32, 2.676214e-32, 2.676203e-32, 2.676209e-32, 
    2.676219e-32, 2.676217e-32, 2.676217e-32, 2.676218e-32, 2.676212e-32, 
    2.676214e-32, 2.676209e-32, 2.676211e-32, 2.676208e-32, 2.676209e-32, 
    2.676209e-32, 2.676211e-32, 2.676212e-32, 2.676214e-32, 2.676216e-32, 
    2.676218e-32, 2.676217e-32, 2.676216e-32, 2.676213e-32, 2.67621e-32, 
    2.67621e-32, 2.676208e-32, 2.676214e-32, 2.676212e-32, 2.676212e-32, 
    2.67621e-32, 2.676215e-32, 2.676211e-32, 2.676216e-32, 2.676216e-32, 
    2.676214e-32, 2.676212e-32, 2.676211e-32, 2.67621e-32, 2.676211e-32, 
    2.676213e-32, 2.676213e-32, 2.676214e-32, 2.676215e-32, 2.676216e-32, 
    2.676217e-32, 2.676216e-32, 2.676215e-32, 2.676213e-32, 2.67621e-32, 
    2.676208e-32, 2.676207e-32, 2.676204e-32, 2.676207e-32, 2.676203e-32, 
    2.676206e-32, 2.6762e-32, 2.676211e-32, 2.676206e-32, 2.676214e-32, 
    2.676214e-32, 2.676212e-32, 2.676208e-32, 2.67621e-32, 2.676208e-32, 
    2.676213e-32, 2.676216e-32, 2.676216e-32, 2.676217e-32, 2.676216e-32, 
    2.676216e-32, 2.676215e-32, 2.676216e-32, 2.676212e-32, 2.676214e-32, 
    2.676209e-32, 2.676208e-32, 2.676203e-32, 2.6762e-32, 2.676197e-32, 
    2.676196e-32, 2.676196e-32, 2.676196e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N_TO_SOIL1N =
  3.414061e-15, 3.422752e-15, 3.421064e-15, 3.428066e-15, 3.424184e-15, 
    3.428767e-15, 3.415825e-15, 3.423095e-15, 3.418456e-15, 3.414846e-15, 
    3.441633e-15, 3.428379e-15, 3.45539e-15, 3.446953e-15, 3.468132e-15, 
    3.454076e-15, 3.470964e-15, 3.46773e-15, 3.477466e-15, 3.474679e-15, 
    3.48711e-15, 3.478752e-15, 3.49355e-15, 3.485117e-15, 3.486435e-15, 
    3.478476e-15, 3.431051e-15, 3.439983e-15, 3.430521e-15, 3.431795e-15, 
    3.431224e-15, 3.424263e-15, 3.42075e-15, 3.413398e-15, 3.414734e-15, 
    3.420135e-15, 3.432369e-15, 3.42822e-15, 3.438677e-15, 3.438441e-15, 
    3.450064e-15, 3.444826e-15, 3.464337e-15, 3.458797e-15, 3.474795e-15, 
    3.470775e-15, 3.474606e-15, 3.473445e-15, 3.474621e-15, 3.468724e-15, 
    3.471251e-15, 3.466061e-15, 3.445807e-15, 3.451764e-15, 3.433981e-15, 
    3.423263e-15, 3.416143e-15, 3.411085e-15, 3.4118e-15, 3.413163e-15, 
    3.420166e-15, 3.426748e-15, 3.431758e-15, 3.435108e-15, 3.438407e-15, 
    3.448377e-15, 3.453655e-15, 3.465454e-15, 3.463329e-15, 3.466931e-15, 
    3.470375e-15, 3.476148e-15, 3.475199e-15, 3.477741e-15, 3.466838e-15, 
    3.474085e-15, 3.462118e-15, 3.465393e-15, 3.439293e-15, 3.42934e-15, 
    3.425096e-15, 3.421388e-15, 3.41235e-15, 3.418592e-15, 3.416132e-15, 
    3.421986e-15, 3.425702e-15, 3.423864e-15, 3.4352e-15, 3.430794e-15, 
    3.453968e-15, 3.443995e-15, 3.469973e-15, 3.463766e-15, 3.471461e-15, 
    3.467536e-15, 3.474259e-15, 3.468208e-15, 3.478687e-15, 3.480966e-15, 
    3.479409e-15, 3.485392e-15, 3.467873e-15, 3.474605e-15, 3.423812e-15, 
    3.424112e-15, 3.425509e-15, 3.419367e-15, 3.418991e-15, 3.413361e-15, 
    3.418372e-15, 3.420504e-15, 3.425918e-15, 3.429116e-15, 3.432156e-15, 
    3.438836e-15, 3.446287e-15, 3.456697e-15, 3.464168e-15, 3.469171e-15, 
    3.466105e-15, 3.468812e-15, 3.465785e-15, 3.464366e-15, 3.480112e-15, 
    3.471274e-15, 3.484532e-15, 3.4838e-15, 3.477801e-15, 3.483882e-15, 
    3.424322e-15, 3.422598e-15, 3.416604e-15, 3.421295e-15, 3.412748e-15, 
    3.417532e-15, 3.420281e-15, 3.430884e-15, 3.433214e-15, 3.435371e-15, 
    3.439631e-15, 3.445094e-15, 3.454666e-15, 3.462987e-15, 3.470575e-15, 
    3.47002e-15, 3.470215e-15, 3.471908e-15, 3.467712e-15, 3.472597e-15, 
    3.473416e-15, 3.471274e-15, 3.483701e-15, 3.480153e-15, 3.483784e-15, 
    3.481474e-15, 3.423159e-15, 3.426061e-15, 3.424493e-15, 3.42744e-15, 
    3.425363e-15, 3.434593e-15, 3.437358e-15, 3.450286e-15, 3.444986e-15, 
    3.453423e-15, 3.445844e-15, 3.447187e-15, 3.453693e-15, 3.446255e-15, 
    3.462526e-15, 3.451495e-15, 3.471974e-15, 3.460968e-15, 3.472663e-15, 
    3.470543e-15, 3.474054e-15, 3.477197e-15, 3.48115e-15, 3.488436e-15, 
    3.48675e-15, 3.492841e-15, 3.430385e-15, 3.434145e-15, 3.433815e-15, 
    3.437749e-15, 3.440656e-15, 3.446956e-15, 3.457047e-15, 3.453254e-15, 
    3.460217e-15, 3.461613e-15, 3.451036e-15, 3.45753e-15, 3.436661e-15, 
    3.440034e-15, 3.438027e-15, 3.430681e-15, 3.454126e-15, 3.442102e-15, 
    3.464291e-15, 3.457789e-15, 3.476749e-15, 3.467324e-15, 3.485821e-15, 
    3.493709e-15, 3.501133e-15, 3.509788e-15, 3.436197e-15, 3.433644e-15, 
    3.438217e-15, 3.444536e-15, 3.4504e-15, 3.458186e-15, 3.458983e-15, 
    3.46044e-15, 3.464215e-15, 3.467386e-15, 3.460898e-15, 3.468181e-15, 
    3.440813e-15, 3.455169e-15, 3.432676e-15, 3.439454e-15, 3.444165e-15, 
    3.442101e-15, 3.452821e-15, 3.455345e-15, 3.465591e-15, 3.460297e-15, 
    3.491761e-15, 3.477858e-15, 3.516377e-15, 3.505633e-15, 3.432751e-15, 
    3.436189e-15, 3.448142e-15, 3.442458e-15, 3.458706e-15, 3.462699e-15, 
    3.465946e-15, 3.47009e-15, 3.470539e-15, 3.472993e-15, 3.46897e-15, 
    3.472835e-15, 3.458202e-15, 3.464745e-15, 3.446779e-15, 3.451155e-15, 
    3.449143e-15, 3.446933e-15, 3.453749e-15, 3.461e-15, 3.461158e-15, 
    3.463481e-15, 3.470017e-15, 3.458772e-15, 3.493548e-15, 3.472086e-15, 
    3.439937e-15, 3.446548e-15, 3.447496e-15, 3.444935e-15, 3.462299e-15, 
    3.456012e-15, 3.472934e-15, 3.468365e-15, 3.47585e-15, 3.472131e-15, 
    3.471584e-15, 3.466805e-15, 3.463828e-15, 3.4563e-15, 3.45017e-15, 
    3.445307e-15, 3.446438e-15, 3.451779e-15, 3.461444e-15, 3.470578e-15, 
    3.468578e-15, 3.475282e-15, 3.457529e-15, 3.464977e-15, 3.462098e-15, 
    3.469602e-15, 3.453153e-15, 3.467153e-15, 3.449569e-15, 3.451113e-15, 
    3.455887e-15, 3.46548e-15, 3.467605e-15, 3.469868e-15, 3.468472e-15, 
    3.46169e-15, 3.46058e-15, 3.455772e-15, 3.454442e-15, 3.450777e-15, 
    3.44774e-15, 3.450514e-15, 3.453426e-15, 3.461694e-15, 3.469136e-15, 
    3.477241e-15, 3.479225e-15, 3.488672e-15, 3.480978e-15, 3.493666e-15, 
    3.482874e-15, 3.501549e-15, 3.467968e-15, 3.482562e-15, 3.456105e-15, 
    3.458961e-15, 3.46412e-15, 3.475945e-15, 3.469567e-15, 3.477027e-15, 
    3.460536e-15, 3.451962e-15, 3.449745e-15, 3.445602e-15, 3.44984e-15, 
    3.449496e-15, 3.453549e-15, 3.452247e-15, 3.461969e-15, 3.456748e-15, 
    3.471569e-15, 3.476969e-15, 3.492201e-15, 3.50152e-15, 3.510999e-15, 
    3.515177e-15, 3.516449e-15, 3.51698e-15 ;

 LITR2N_vr =
  1.532729e-05, 1.532728e-05, 1.532728e-05, 1.532727e-05, 1.532728e-05, 
    1.532727e-05, 1.532729e-05, 1.532728e-05, 1.532729e-05, 1.532729e-05, 
    1.532725e-05, 1.532727e-05, 1.532722e-05, 1.532724e-05, 1.53272e-05, 
    1.532722e-05, 1.53272e-05, 1.53272e-05, 1.532718e-05, 1.532719e-05, 
    1.532717e-05, 1.532718e-05, 1.532716e-05, 1.532717e-05, 1.532717e-05, 
    1.532718e-05, 1.532726e-05, 1.532725e-05, 1.532726e-05, 1.532726e-05, 
    1.532726e-05, 1.532728e-05, 1.532728e-05, 1.53273e-05, 1.532729e-05, 
    1.532728e-05, 1.532726e-05, 1.532727e-05, 1.532725e-05, 1.532725e-05, 
    1.532723e-05, 1.532724e-05, 1.532721e-05, 1.532722e-05, 1.532719e-05, 
    1.53272e-05, 1.532719e-05, 1.532719e-05, 1.532719e-05, 1.53272e-05, 
    1.532719e-05, 1.53272e-05, 1.532724e-05, 1.532723e-05, 1.532726e-05, 
    1.532728e-05, 1.532729e-05, 1.53273e-05, 1.53273e-05, 1.53273e-05, 
    1.532728e-05, 1.532727e-05, 1.532726e-05, 1.532726e-05, 1.532725e-05, 
    1.532723e-05, 1.532722e-05, 1.53272e-05, 1.532721e-05, 1.53272e-05, 
    1.53272e-05, 1.532719e-05, 1.532719e-05, 1.532718e-05, 1.53272e-05, 
    1.532719e-05, 1.532721e-05, 1.53272e-05, 1.532725e-05, 1.532727e-05, 
    1.532728e-05, 1.532728e-05, 1.53273e-05, 1.532729e-05, 1.532729e-05, 
    1.532728e-05, 1.532727e-05, 1.532728e-05, 1.532726e-05, 1.532726e-05, 
    1.532722e-05, 1.532724e-05, 1.53272e-05, 1.532721e-05, 1.532719e-05, 
    1.53272e-05, 1.532719e-05, 1.53272e-05, 1.532718e-05, 1.532718e-05, 
    1.532718e-05, 1.532717e-05, 1.53272e-05, 1.532719e-05, 1.532728e-05, 
    1.532728e-05, 1.532727e-05, 1.532728e-05, 1.532728e-05, 1.53273e-05, 
    1.532729e-05, 1.532728e-05, 1.532727e-05, 1.532727e-05, 1.532726e-05, 
    1.532725e-05, 1.532724e-05, 1.532722e-05, 1.532721e-05, 1.53272e-05, 
    1.53272e-05, 1.53272e-05, 1.53272e-05, 1.532721e-05, 1.532718e-05, 
    1.532719e-05, 1.532717e-05, 1.532717e-05, 1.532718e-05, 1.532717e-05, 
    1.532728e-05, 1.532728e-05, 1.532729e-05, 1.532728e-05, 1.53273e-05, 
    1.532729e-05, 1.532728e-05, 1.532726e-05, 1.532726e-05, 1.532726e-05, 
    1.532725e-05, 1.532724e-05, 1.532722e-05, 1.532721e-05, 1.53272e-05, 
    1.53272e-05, 1.53272e-05, 1.532719e-05, 1.53272e-05, 1.532719e-05, 
    1.532719e-05, 1.532719e-05, 1.532717e-05, 1.532718e-05, 1.532717e-05, 
    1.532718e-05, 1.532728e-05, 1.532727e-05, 1.532728e-05, 1.532727e-05, 
    1.532727e-05, 1.532726e-05, 1.532725e-05, 1.532723e-05, 1.532724e-05, 
    1.532722e-05, 1.532724e-05, 1.532724e-05, 1.532722e-05, 1.532724e-05, 
    1.532721e-05, 1.532723e-05, 1.532719e-05, 1.532721e-05, 1.532719e-05, 
    1.53272e-05, 1.532719e-05, 1.532718e-05, 1.532718e-05, 1.532716e-05, 
    1.532717e-05, 1.532716e-05, 1.532727e-05, 1.532726e-05, 1.532726e-05, 
    1.532725e-05, 1.532725e-05, 1.532724e-05, 1.532722e-05, 1.532723e-05, 
    1.532721e-05, 1.532721e-05, 1.532723e-05, 1.532722e-05, 1.532725e-05, 
    1.532725e-05, 1.532725e-05, 1.532726e-05, 1.532722e-05, 1.532724e-05, 
    1.532721e-05, 1.532722e-05, 1.532718e-05, 1.53272e-05, 1.532717e-05, 
    1.532716e-05, 1.532714e-05, 1.532713e-05, 1.532726e-05, 1.532726e-05, 
    1.532725e-05, 1.532724e-05, 1.532723e-05, 1.532722e-05, 1.532722e-05, 
    1.532721e-05, 1.532721e-05, 1.53272e-05, 1.532721e-05, 1.53272e-05, 
    1.532725e-05, 1.532722e-05, 1.532726e-05, 1.532725e-05, 1.532724e-05, 
    1.532724e-05, 1.532723e-05, 1.532722e-05, 1.53272e-05, 1.532721e-05, 
    1.532716e-05, 1.532718e-05, 1.532712e-05, 1.532713e-05, 1.532726e-05, 
    1.532726e-05, 1.532723e-05, 1.532724e-05, 1.532722e-05, 1.532721e-05, 
    1.53272e-05, 1.53272e-05, 1.53272e-05, 1.532719e-05, 1.53272e-05, 
    1.532719e-05, 1.532722e-05, 1.532721e-05, 1.532724e-05, 1.532723e-05, 
    1.532723e-05, 1.532724e-05, 1.532722e-05, 1.532721e-05, 1.532721e-05, 
    1.532721e-05, 1.53272e-05, 1.532722e-05, 1.532716e-05, 1.532719e-05, 
    1.532725e-05, 1.532724e-05, 1.532724e-05, 1.532724e-05, 1.532721e-05, 
    1.532722e-05, 1.532719e-05, 1.53272e-05, 1.532719e-05, 1.532719e-05, 
    1.532719e-05, 1.53272e-05, 1.532721e-05, 1.532722e-05, 1.532723e-05, 
    1.532724e-05, 1.532724e-05, 1.532723e-05, 1.532721e-05, 1.53272e-05, 
    1.53272e-05, 1.532719e-05, 1.532722e-05, 1.53272e-05, 1.532721e-05, 
    1.53272e-05, 1.532723e-05, 1.53272e-05, 1.532723e-05, 1.532723e-05, 
    1.532722e-05, 1.53272e-05, 1.53272e-05, 1.53272e-05, 1.53272e-05, 
    1.532721e-05, 1.532721e-05, 1.532722e-05, 1.532722e-05, 1.532723e-05, 
    1.532724e-05, 1.532723e-05, 1.532722e-05, 1.532721e-05, 1.53272e-05, 
    1.532718e-05, 1.532718e-05, 1.532716e-05, 1.532718e-05, 1.532716e-05, 
    1.532717e-05, 1.532714e-05, 1.53272e-05, 1.532717e-05, 1.532722e-05, 
    1.532722e-05, 1.532721e-05, 1.532719e-05, 1.53272e-05, 1.532718e-05, 
    1.532721e-05, 1.532723e-05, 1.532723e-05, 1.532724e-05, 1.532723e-05, 
    1.532723e-05, 1.532722e-05, 1.532723e-05, 1.532721e-05, 1.532722e-05, 
    1.532719e-05, 1.532718e-05, 1.532716e-05, 1.532714e-05, 1.532712e-05, 
    1.532712e-05, 1.532712e-05, 1.532711e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2_HR =
  1.233469e-13, 1.236609e-13, 1.235999e-13, 1.238529e-13, 1.237126e-13, 
    1.238782e-13, 1.234106e-13, 1.236733e-13, 1.235057e-13, 1.233753e-13, 
    1.243431e-13, 1.238642e-13, 1.248401e-13, 1.245353e-13, 1.253005e-13, 
    1.247926e-13, 1.254028e-13, 1.252859e-13, 1.256377e-13, 1.25537e-13, 
    1.259861e-13, 1.256841e-13, 1.262188e-13, 1.259141e-13, 1.259617e-13, 
    1.256742e-13, 1.239607e-13, 1.242835e-13, 1.239416e-13, 1.239876e-13, 
    1.23967e-13, 1.237155e-13, 1.235886e-13, 1.23323e-13, 1.233712e-13, 
    1.235663e-13, 1.240083e-13, 1.238585e-13, 1.242363e-13, 1.242277e-13, 
    1.246477e-13, 1.244584e-13, 1.251633e-13, 1.249632e-13, 1.255412e-13, 
    1.253959e-13, 1.255343e-13, 1.254924e-13, 1.255349e-13, 1.253218e-13, 
    1.254131e-13, 1.252256e-13, 1.244939e-13, 1.247091e-13, 1.240666e-13, 
    1.236794e-13, 1.234221e-13, 1.232394e-13, 1.232652e-13, 1.233145e-13, 
    1.235675e-13, 1.238053e-13, 1.239863e-13, 1.241073e-13, 1.242265e-13, 
    1.245867e-13, 1.247774e-13, 1.252037e-13, 1.251269e-13, 1.252571e-13, 
    1.253815e-13, 1.255901e-13, 1.255558e-13, 1.256476e-13, 1.252537e-13, 
    1.255155e-13, 1.250832e-13, 1.252015e-13, 1.242585e-13, 1.238989e-13, 
    1.237456e-13, 1.236116e-13, 1.232851e-13, 1.235106e-13, 1.234217e-13, 
    1.236332e-13, 1.237675e-13, 1.237011e-13, 1.241106e-13, 1.239515e-13, 
    1.247887e-13, 1.244284e-13, 1.25367e-13, 1.251427e-13, 1.254207e-13, 
    1.252789e-13, 1.255218e-13, 1.253032e-13, 1.256818e-13, 1.257641e-13, 
    1.257079e-13, 1.259241e-13, 1.252911e-13, 1.255343e-13, 1.236992e-13, 
    1.2371e-13, 1.237605e-13, 1.235386e-13, 1.23525e-13, 1.233216e-13, 
    1.235026e-13, 1.235797e-13, 1.237753e-13, 1.238908e-13, 1.240007e-13, 
    1.24242e-13, 1.245112e-13, 1.248873e-13, 1.251572e-13, 1.25338e-13, 
    1.252272e-13, 1.25325e-13, 1.252156e-13, 1.251644e-13, 1.257333e-13, 
    1.254139e-13, 1.25893e-13, 1.258665e-13, 1.256498e-13, 1.258695e-13, 
    1.237176e-13, 1.236553e-13, 1.234388e-13, 1.236083e-13, 1.232995e-13, 
    1.234723e-13, 1.235716e-13, 1.239547e-13, 1.240389e-13, 1.241168e-13, 
    1.242707e-13, 1.244681e-13, 1.24814e-13, 1.251145e-13, 1.253887e-13, 
    1.253687e-13, 1.253757e-13, 1.254369e-13, 1.252853e-13, 1.254618e-13, 
    1.254913e-13, 1.25414e-13, 1.258629e-13, 1.257348e-13, 1.258659e-13, 
    1.257825e-13, 1.236756e-13, 1.237804e-13, 1.237238e-13, 1.238303e-13, 
    1.237552e-13, 1.240887e-13, 1.241886e-13, 1.246557e-13, 1.244642e-13, 
    1.24769e-13, 1.244952e-13, 1.245437e-13, 1.247788e-13, 1.2451e-13, 
    1.250979e-13, 1.246994e-13, 1.254393e-13, 1.250416e-13, 1.254641e-13, 
    1.253875e-13, 1.255144e-13, 1.25628e-13, 1.257708e-13, 1.26034e-13, 
    1.259731e-13, 1.261931e-13, 1.239367e-13, 1.240725e-13, 1.240606e-13, 
    1.242027e-13, 1.243078e-13, 1.245354e-13, 1.248999e-13, 1.247629e-13, 
    1.250145e-13, 1.250649e-13, 1.246828e-13, 1.249174e-13, 1.241634e-13, 
    1.242853e-13, 1.242128e-13, 1.239474e-13, 1.247944e-13, 1.2436e-13, 
    1.251617e-13, 1.249268e-13, 1.256118e-13, 1.252713e-13, 1.259395e-13, 
    1.262245e-13, 1.264927e-13, 1.268054e-13, 1.241467e-13, 1.240544e-13, 
    1.242196e-13, 1.24448e-13, 1.246598e-13, 1.249411e-13, 1.249699e-13, 
    1.250225e-13, 1.251589e-13, 1.252735e-13, 1.250391e-13, 1.253022e-13, 
    1.243134e-13, 1.248321e-13, 1.240195e-13, 1.242643e-13, 1.244345e-13, 
    1.2436e-13, 1.247473e-13, 1.248385e-13, 1.252086e-13, 1.250174e-13, 
    1.261541e-13, 1.256518e-13, 1.270435e-13, 1.266553e-13, 1.240222e-13, 
    1.241464e-13, 1.245782e-13, 1.243728e-13, 1.249599e-13, 1.251042e-13, 
    1.252215e-13, 1.253712e-13, 1.253874e-13, 1.254761e-13, 1.253307e-13, 
    1.254704e-13, 1.249417e-13, 1.251781e-13, 1.24529e-13, 1.246871e-13, 
    1.246144e-13, 1.245346e-13, 1.247808e-13, 1.250428e-13, 1.250485e-13, 
    1.251324e-13, 1.253685e-13, 1.249623e-13, 1.262187e-13, 1.254433e-13, 
    1.242818e-13, 1.245206e-13, 1.245549e-13, 1.244624e-13, 1.250897e-13, 
    1.248625e-13, 1.254739e-13, 1.253089e-13, 1.255793e-13, 1.254449e-13, 
    1.254252e-13, 1.252525e-13, 1.251449e-13, 1.24873e-13, 1.246515e-13, 
    1.244758e-13, 1.245167e-13, 1.247096e-13, 1.250588e-13, 1.253888e-13, 
    1.253165e-13, 1.255588e-13, 1.249174e-13, 1.251865e-13, 1.250825e-13, 
    1.253536e-13, 1.247593e-13, 1.252651e-13, 1.246298e-13, 1.246856e-13, 
    1.248581e-13, 1.252046e-13, 1.252814e-13, 1.253632e-13, 1.253127e-13, 
    1.250677e-13, 1.250276e-13, 1.248539e-13, 1.248058e-13, 1.246734e-13, 
    1.245637e-13, 1.246639e-13, 1.247691e-13, 1.250679e-13, 1.253367e-13, 
    1.256296e-13, 1.257012e-13, 1.260426e-13, 1.257646e-13, 1.26223e-13, 
    1.25833e-13, 1.265078e-13, 1.252945e-13, 1.258218e-13, 1.248659e-13, 
    1.249691e-13, 1.251555e-13, 1.255827e-13, 1.253523e-13, 1.256218e-13, 
    1.25026e-13, 1.247162e-13, 1.246362e-13, 1.244865e-13, 1.246396e-13, 
    1.246271e-13, 1.247736e-13, 1.247265e-13, 1.250778e-13, 1.248892e-13, 
    1.254246e-13, 1.256197e-13, 1.2617e-13, 1.265067e-13, 1.268492e-13, 
    1.270001e-13, 1.270461e-13, 1.270653e-13 ;

 LITR3C =
  9.697916e-06, 9.697906e-06, 9.697907e-06, 9.6979e-06, 9.697904e-06, 
    9.697899e-06, 9.697914e-06, 9.697906e-06, 9.69791e-06, 9.697915e-06, 
    9.697885e-06, 9.697899e-06, 9.69787e-06, 9.697879e-06, 9.697856e-06, 
    9.697871e-06, 9.697853e-06, 9.697857e-06, 9.697846e-06, 9.697848e-06, 
    9.697835e-06, 9.697844e-06, 9.697827e-06, 9.697837e-06, 9.697836e-06, 
    9.697845e-06, 9.697897e-06, 9.697887e-06, 9.697897e-06, 9.697896e-06, 
    9.697897e-06, 9.697904e-06, 9.697908e-06, 9.697917e-06, 9.697915e-06, 
    9.697908e-06, 9.697896e-06, 9.6979e-06, 9.697888e-06, 9.697888e-06, 
    9.697876e-06, 9.697881e-06, 9.69786e-06, 9.697866e-06, 9.697848e-06, 
    9.697853e-06, 9.697848e-06, 9.69785e-06, 9.697848e-06, 9.697855e-06, 
    9.697852e-06, 9.697858e-06, 9.69788e-06, 9.697874e-06, 9.697894e-06, 
    9.697906e-06, 9.697913e-06, 9.697918e-06, 9.697918e-06, 9.697917e-06, 
    9.697908e-06, 9.697901e-06, 9.697896e-06, 9.697892e-06, 9.697888e-06, 
    9.697877e-06, 9.697872e-06, 9.697858e-06, 9.697861e-06, 9.697857e-06, 
    9.697853e-06, 9.697847e-06, 9.697848e-06, 9.697845e-06, 9.697857e-06, 
    9.697849e-06, 9.697862e-06, 9.697858e-06, 9.697887e-06, 9.697898e-06, 
    9.697903e-06, 9.697907e-06, 9.697917e-06, 9.69791e-06, 9.697913e-06, 
    9.697907e-06, 9.697903e-06, 9.697905e-06, 9.697892e-06, 9.697897e-06, 
    9.697871e-06, 9.697882e-06, 9.697854e-06, 9.69786e-06, 9.697852e-06, 
    9.697857e-06, 9.697849e-06, 9.697856e-06, 9.697844e-06, 9.697842e-06, 
    9.697843e-06, 9.697837e-06, 9.697856e-06, 9.697848e-06, 9.697905e-06, 
    9.697905e-06, 9.697903e-06, 9.697909e-06, 9.69791e-06, 9.697917e-06, 
    9.697911e-06, 9.697908e-06, 9.697902e-06, 9.697898e-06, 9.697896e-06, 
    9.697888e-06, 9.69788e-06, 9.697868e-06, 9.69786e-06, 9.697855e-06, 
    9.697858e-06, 9.697855e-06, 9.697858e-06, 9.69786e-06, 9.697843e-06, 
    9.697852e-06, 9.697837e-06, 9.697838e-06, 9.697845e-06, 9.697838e-06, 
    9.697904e-06, 9.697906e-06, 9.697913e-06, 9.697907e-06, 9.697917e-06, 
    9.697912e-06, 9.697908e-06, 9.697897e-06, 9.697895e-06, 9.697892e-06, 
    9.697887e-06, 9.697881e-06, 9.69787e-06, 9.697861e-06, 9.697853e-06, 
    9.697854e-06, 9.697854e-06, 9.697852e-06, 9.697857e-06, 9.697851e-06, 
    9.69785e-06, 9.697852e-06, 9.697838e-06, 9.697843e-06, 9.697838e-06, 
    9.697841e-06, 9.697906e-06, 9.697902e-06, 9.697904e-06, 9.697901e-06, 
    9.697903e-06, 9.697893e-06, 9.697889e-06, 9.697876e-06, 9.697881e-06, 
    9.697872e-06, 9.69788e-06, 9.697879e-06, 9.697872e-06, 9.69788e-06, 
    9.697862e-06, 9.697874e-06, 9.697851e-06, 9.697864e-06, 9.697851e-06, 
    9.697853e-06, 9.697849e-06, 9.697846e-06, 9.697841e-06, 9.697833e-06, 
    9.697836e-06, 9.697828e-06, 9.697897e-06, 9.697893e-06, 9.697894e-06, 
    9.697889e-06, 9.697886e-06, 9.697879e-06, 9.697868e-06, 9.697872e-06, 
    9.697865e-06, 9.697863e-06, 9.697875e-06, 9.697867e-06, 9.69789e-06, 
    9.697887e-06, 9.697889e-06, 9.697897e-06, 9.697871e-06, 9.697885e-06, 
    9.69786e-06, 9.697867e-06, 9.697847e-06, 9.697857e-06, 9.697837e-06, 
    9.697827e-06, 9.697819e-06, 9.69781e-06, 9.697891e-06, 9.697894e-06, 
    9.697888e-06, 9.697882e-06, 9.697876e-06, 9.697867e-06, 9.697866e-06, 
    9.697864e-06, 9.69786e-06, 9.697857e-06, 9.697864e-06, 9.697856e-06, 
    9.697886e-06, 9.69787e-06, 9.697895e-06, 9.697887e-06, 9.697882e-06, 
    9.697885e-06, 9.697873e-06, 9.69787e-06, 9.697858e-06, 9.697865e-06, 
    9.697829e-06, 9.697845e-06, 9.697803e-06, 9.697815e-06, 9.697895e-06, 
    9.697891e-06, 9.697877e-06, 9.697884e-06, 9.697867e-06, 9.697862e-06, 
    9.697858e-06, 9.697854e-06, 9.697853e-06, 9.69785e-06, 9.697855e-06, 
    9.69785e-06, 9.697867e-06, 9.697859e-06, 9.697879e-06, 9.697875e-06, 
    9.697877e-06, 9.697879e-06, 9.697872e-06, 9.697864e-06, 9.697864e-06, 
    9.697861e-06, 9.697854e-06, 9.697866e-06, 9.697827e-06, 9.697851e-06, 
    9.697887e-06, 9.697879e-06, 9.697878e-06, 9.697881e-06, 9.697862e-06, 
    9.697869e-06, 9.69785e-06, 9.697856e-06, 9.697847e-06, 9.697851e-06, 
    9.697852e-06, 9.697857e-06, 9.69786e-06, 9.697868e-06, 9.697876e-06, 
    9.697881e-06, 9.697879e-06, 9.697874e-06, 9.697863e-06, 9.697853e-06, 
    9.697856e-06, 9.697847e-06, 9.697867e-06, 9.697859e-06, 9.697862e-06, 
    9.697854e-06, 9.697872e-06, 9.697857e-06, 9.697877e-06, 9.697875e-06, 
    9.697869e-06, 9.697858e-06, 9.697857e-06, 9.697854e-06, 9.697856e-06, 
    9.697863e-06, 9.697864e-06, 9.697869e-06, 9.697871e-06, 9.697875e-06, 
    9.697878e-06, 9.697876e-06, 9.697872e-06, 9.697863e-06, 9.697855e-06, 
    9.697846e-06, 9.697844e-06, 9.697833e-06, 9.697842e-06, 9.697827e-06, 
    9.697839e-06, 9.697819e-06, 9.697856e-06, 9.69784e-06, 9.697869e-06, 
    9.697866e-06, 9.69786e-06, 9.697847e-06, 9.697854e-06, 9.697846e-06, 
    9.697864e-06, 9.697874e-06, 9.697876e-06, 9.69788e-06, 9.697876e-06, 
    9.697877e-06, 9.697872e-06, 9.697873e-06, 9.697863e-06, 9.697868e-06, 
    9.697852e-06, 9.697846e-06, 9.697829e-06, 9.697819e-06, 9.697808e-06, 
    9.697804e-06, 9.697802e-06, 9.697802e-06 ;

 LITR3C_TO_SOIL2C =
  6.167343e-14, 6.183042e-14, 6.179994e-14, 6.192643e-14, 6.18563e-14, 
    6.193909e-14, 6.17053e-14, 6.183664e-14, 6.175282e-14, 6.168761e-14, 
    6.217151e-14, 6.193208e-14, 6.242002e-14, 6.226761e-14, 6.265021e-14, 
    6.239628e-14, 6.270136e-14, 6.264295e-14, 6.281882e-14, 6.276846e-14, 
    6.299303e-14, 6.284206e-14, 6.310938e-14, 6.295702e-14, 6.298084e-14, 
    6.283706e-14, 6.198036e-14, 6.214171e-14, 6.197077e-14, 6.19938e-14, 
    6.198348e-14, 6.185773e-14, 6.179427e-14, 6.166146e-14, 6.168559e-14, 
    6.178315e-14, 6.200415e-14, 6.192921e-14, 6.211812e-14, 6.211385e-14, 
    6.232382e-14, 6.222919e-14, 6.258164e-14, 6.248158e-14, 6.277057e-14, 
    6.269794e-14, 6.276715e-14, 6.274617e-14, 6.276742e-14, 6.26609e-14, 
    6.270654e-14, 6.261278e-14, 6.224691e-14, 6.235452e-14, 6.203327e-14, 
    6.183966e-14, 6.171105e-14, 6.161968e-14, 6.16326e-14, 6.165722e-14, 
    6.178372e-14, 6.190261e-14, 6.199314e-14, 6.205364e-14, 6.211324e-14, 
    6.229334e-14, 6.238869e-14, 6.260183e-14, 6.256345e-14, 6.262851e-14, 
    6.269072e-14, 6.279502e-14, 6.277786e-14, 6.282378e-14, 6.262683e-14, 
    6.275774e-14, 6.254156e-14, 6.260072e-14, 6.212924e-14, 6.194944e-14, 
    6.187278e-14, 6.180579e-14, 6.164253e-14, 6.175528e-14, 6.171084e-14, 
    6.181659e-14, 6.188371e-14, 6.185053e-14, 6.205529e-14, 6.197571e-14, 
    6.239434e-14, 6.221418e-14, 6.268346e-14, 6.257133e-14, 6.271033e-14, 
    6.263943e-14, 6.276088e-14, 6.265158e-14, 6.284089e-14, 6.288205e-14, 
    6.285392e-14, 6.296201e-14, 6.264551e-14, 6.276713e-14, 6.184959e-14, 
    6.1855e-14, 6.188023e-14, 6.176927e-14, 6.17625e-14, 6.166079e-14, 
    6.175131e-14, 6.178982e-14, 6.188762e-14, 6.19454e-14, 6.200031e-14, 
    6.212098e-14, 6.225558e-14, 6.244363e-14, 6.25786e-14, 6.266898e-14, 
    6.261358e-14, 6.266249e-14, 6.26078e-14, 6.258218e-14, 6.286661e-14, 
    6.270695e-14, 6.294646e-14, 6.293323e-14, 6.282487e-14, 6.293472e-14, 
    6.18588e-14, 6.182765e-14, 6.171937e-14, 6.180412e-14, 6.164971e-14, 
    6.173614e-14, 6.17858e-14, 6.197734e-14, 6.201943e-14, 6.205839e-14, 
    6.213535e-14, 6.223403e-14, 6.240695e-14, 6.255726e-14, 6.269434e-14, 
    6.268431e-14, 6.268784e-14, 6.271843e-14, 6.264262e-14, 6.273087e-14, 
    6.274565e-14, 6.270696e-14, 6.293146e-14, 6.286736e-14, 6.293295e-14, 
    6.289123e-14, 6.183778e-14, 6.18902e-14, 6.186188e-14, 6.191513e-14, 
    6.18776e-14, 6.204434e-14, 6.209428e-14, 6.232783e-14, 6.223208e-14, 
    6.238448e-14, 6.224758e-14, 6.227184e-14, 6.238938e-14, 6.2255e-14, 
    6.254894e-14, 6.234965e-14, 6.271961e-14, 6.25208e-14, 6.273206e-14, 
    6.269375e-14, 6.275719e-14, 6.281396e-14, 6.288537e-14, 6.301699e-14, 
    6.298653e-14, 6.309655e-14, 6.196833e-14, 6.203623e-14, 6.203029e-14, 
    6.210135e-14, 6.215386e-14, 6.226767e-14, 6.244995e-14, 6.238144e-14, 
    6.250722e-14, 6.253244e-14, 6.234137e-14, 6.245868e-14, 6.208169e-14, 
    6.214263e-14, 6.210637e-14, 6.197367e-14, 6.239718e-14, 6.217998e-14, 
    6.258082e-14, 6.246337e-14, 6.280586e-14, 6.263561e-14, 6.296976e-14, 
    6.311224e-14, 6.324635e-14, 6.34027e-14, 6.207332e-14, 6.202719e-14, 
    6.21098e-14, 6.222396e-14, 6.232989e-14, 6.247053e-14, 6.248493e-14, 
    6.251125e-14, 6.257944e-14, 6.263672e-14, 6.251954e-14, 6.265108e-14, 
    6.215669e-14, 6.241604e-14, 6.200972e-14, 6.213215e-14, 6.221725e-14, 
    6.217996e-14, 6.237362e-14, 6.241921e-14, 6.26043e-14, 6.250867e-14, 
    6.307705e-14, 6.282589e-14, 6.352174e-14, 6.332765e-14, 6.201106e-14, 
    6.207318e-14, 6.228908e-14, 6.21864e-14, 6.247993e-14, 6.255207e-14, 
    6.261071e-14, 6.268557e-14, 6.269368e-14, 6.273802e-14, 6.266535e-14, 
    6.273516e-14, 6.247083e-14, 6.258903e-14, 6.226446e-14, 6.234352e-14, 
    6.230717e-14, 6.226726e-14, 6.239038e-14, 6.252137e-14, 6.252422e-14, 
    6.256619e-14, 6.268426e-14, 6.248112e-14, 6.310932e-14, 6.272162e-14, 
    6.214087e-14, 6.22603e-14, 6.227742e-14, 6.223116e-14, 6.254483e-14, 
    6.243126e-14, 6.273695e-14, 6.265442e-14, 6.278963e-14, 6.272245e-14, 
    6.271256e-14, 6.262623e-14, 6.257244e-14, 6.243646e-14, 6.232572e-14, 
    6.223788e-14, 6.225832e-14, 6.235479e-14, 6.252939e-14, 6.269439e-14, 
    6.265825e-14, 6.277936e-14, 6.245867e-14, 6.259321e-14, 6.254121e-14, 
    6.267677e-14, 6.237961e-14, 6.263252e-14, 6.231487e-14, 6.234276e-14, 
    6.2429e-14, 6.260229e-14, 6.264068e-14, 6.268156e-14, 6.265635e-14, 
    6.253383e-14, 6.251378e-14, 6.242692e-14, 6.24029e-14, 6.233669e-14, 
    6.228182e-14, 6.233194e-14, 6.238455e-14, 6.253391e-14, 6.266834e-14, 
    6.281476e-14, 6.285058e-14, 6.302126e-14, 6.288226e-14, 6.311147e-14, 
    6.29165e-14, 6.325387e-14, 6.264725e-14, 6.291089e-14, 6.243295e-14, 
    6.248454e-14, 6.257773e-14, 6.279135e-14, 6.267613e-14, 6.281089e-14, 
    6.251299e-14, 6.235809e-14, 6.231806e-14, 6.224321e-14, 6.231977e-14, 
    6.231354e-14, 6.238676e-14, 6.236324e-14, 6.253886e-14, 6.244456e-14, 
    6.27123e-14, 6.280985e-14, 6.3085e-14, 6.325334e-14, 6.342457e-14, 
    6.350005e-14, 6.352302e-14, 6.353261e-14 ;

 LITR3C_vr =
  0.000553761, 0.0005537604, 0.0005537606, 0.0005537601, 0.0005537603, 
    0.00055376, 0.0005537609, 0.0005537604, 0.0005537607, 0.000553761, 
    0.0005537593, 0.0005537601, 0.0005537584, 0.0005537589, 0.0005537576, 
    0.0005537585, 0.0005537574, 0.0005537576, 0.000553757, 0.0005537572, 
    0.0005537564, 0.0005537569, 0.000553756, 0.0005537565, 0.0005537564, 
    0.000553757, 0.0005537599, 0.0005537593, 0.00055376, 0.0005537599, 
    0.0005537599, 0.0005537603, 0.0005537606, 0.000553761, 0.000553761, 
    0.0005537606, 0.0005537599, 0.0005537601, 0.0005537595, 0.0005537595, 
    0.0005537587, 0.000553759, 0.0005537578, 0.0005537582, 0.0005537572, 
    0.0005537574, 0.0005537572, 0.0005537572, 0.0005537572, 0.0005537575, 
    0.0005537574, 0.0005537577, 0.000553759, 0.0005537586, 0.0005537597, 
    0.0005537604, 0.0005537609, 0.0005537612, 0.0005537611, 0.000553761, 
    0.0005537606, 0.0005537602, 0.0005537599, 0.0005537597, 0.0005537595, 
    0.0005537588, 0.0005537585, 0.0005537578, 0.0005537579, 0.0005537577, 
    0.0005537574, 0.0005537571, 0.0005537571, 0.000553757, 0.0005537577, 
    0.0005537572, 0.0005537579, 0.0005537578, 0.0005537594, 0.00055376, 
    0.0005537603, 0.0005537605, 0.0005537611, 0.0005537607, 0.0005537609, 
    0.0005537605, 0.0005537603, 0.0005537604, 0.0005537597, 0.0005537599, 
    0.0005537585, 0.0005537591, 0.0005537575, 0.0005537579, 0.0005537574, 
    0.0005537576, 0.0005537572, 0.0005537576, 0.0005537569, 0.0005537568, 
    0.0005537569, 0.0005537565, 0.0005537576, 0.0005537572, 0.0005537604, 
    0.0005537604, 0.0005537603, 0.0005537607, 0.0005537607, 0.000553761, 
    0.0005537607, 0.0005537606, 0.0005537603, 0.00055376, 0.0005537599, 
    0.0005537595, 0.0005537589, 0.0005537583, 0.0005537578, 0.0005537575, 
    0.0005537577, 0.0005537575, 0.0005537577, 0.0005537578, 0.0005537568, 
    0.0005537574, 0.0005537565, 0.0005537566, 0.000553757, 0.0005537566, 
    0.0005537603, 0.0005537604, 0.0005537609, 0.0005537606, 0.0005537611, 
    0.0005537608, 0.0005537606, 0.0005537599, 0.0005537598, 0.0005537596, 
    0.0005537594, 0.000553759, 0.0005537584, 0.0005537579, 0.0005537574, 
    0.0005537575, 0.0005537575, 0.0005537574, 0.0005537576, 0.0005537573, 
    0.0005537572, 0.0005537574, 0.0005537566, 0.0005537568, 0.0005537566, 
    0.0005537567, 0.0005537604, 0.0005537602, 0.0005537603, 0.0005537602, 
    0.0005537603, 0.0005537597, 0.0005537595, 0.0005537587, 0.000553759, 
    0.0005537585, 0.000553759, 0.0005537589, 0.0005537585, 0.000553759, 
    0.0005537579, 0.0005537586, 0.0005537574, 0.0005537581, 0.0005537573, 
    0.0005537574, 0.0005537572, 0.000553757, 0.0005537568, 0.0005537563, 
    0.0005537564, 0.000553756, 0.00055376, 0.0005537597, 0.0005537597, 
    0.0005537595, 0.0005537593, 0.0005537589, 0.0005537583, 0.0005537585, 
    0.0005537581, 0.000553758, 0.0005537586, 0.0005537582, 0.0005537596, 
    0.0005537593, 0.0005537595, 0.0005537599, 0.0005537585, 0.0005537592, 
    0.0005537578, 0.0005537582, 0.0005537571, 0.0005537577, 0.0005537565, 
    0.000553756, 0.0005537555, 0.000553755, 0.0005537596, 0.0005537597, 
    0.0005537595, 0.000553759, 0.0005537587, 0.0005537582, 0.0005537582, 
    0.0005537581, 0.0005537578, 0.0005537577, 0.0005537581, 0.0005537576, 
    0.0005537593, 0.0005537584, 0.0005537598, 0.0005537594, 0.0005537591, 
    0.0005537592, 0.0005537585, 0.0005537584, 0.0005537578, 0.0005537581, 
    0.0005537561, 0.000553757, 0.0005537546, 0.0005537552, 0.0005537598, 
    0.0005537596, 0.0005537588, 0.0005537592, 0.0005537582, 0.0005537579, 
    0.0005537577, 0.0005537575, 0.0005537574, 0.0005537573, 0.0005537575, 
    0.0005537573, 0.0005537582, 0.0005537578, 0.0005537589, 0.0005537586, 
    0.0005537588, 0.0005537589, 0.0005537585, 0.0005537581, 0.000553758, 
    0.0005537579, 0.0005537575, 0.0005537582, 0.000553756, 0.0005537574, 
    0.0005537593, 0.0005537589, 0.0005537589, 0.000553759, 0.0005537579, 
    0.0005537583, 0.0005537573, 0.0005537576, 0.0005537571, 0.0005537574, 
    0.0005537574, 0.0005537577, 0.0005537578, 0.0005537583, 0.0005537587, 
    0.000553759, 0.0005537589, 0.0005537586, 0.000553758, 0.0005537574, 
    0.0005537575, 0.0005537571, 0.0005537582, 0.0005537578, 0.0005537579, 
    0.0005537575, 0.0005537585, 0.0005537577, 0.0005537588, 0.0005537586, 
    0.0005537583, 0.0005537578, 0.0005537576, 0.0005537575, 0.0005537575, 
    0.000553758, 0.0005537581, 0.0005537583, 0.0005537585, 0.0005537587, 
    0.0005537589, 0.0005537587, 0.0005537585, 0.000553758, 0.0005537575, 
    0.000553757, 0.0005537569, 0.0005537563, 0.0005537568, 0.000553756, 
    0.0005537567, 0.0005537555, 0.0005537576, 0.0005537567, 0.0005537583, 
    0.0005537582, 0.0005537578, 0.0005537571, 0.0005537575, 0.000553757, 
    0.0005537581, 0.0005537586, 0.0005537588, 0.000553759, 0.0005537588, 
    0.0005537588, 0.0005537585, 0.0005537586, 0.000553758, 0.0005537583, 
    0.0005537574, 0.000553757, 0.0005537561, 0.0005537555, 0.0005537549, 
    0.0005537546, 0.0005537545, 0.0005537545,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N =
  1.342121e-07, 1.342119e-07, 1.342119e-07, 1.342118e-07, 1.342119e-07, 
    1.342118e-07, 1.34212e-07, 1.342119e-07, 1.34212e-07, 1.34212e-07, 
    1.342116e-07, 1.342118e-07, 1.342114e-07, 1.342115e-07, 1.342112e-07, 
    1.342114e-07, 1.342112e-07, 1.342112e-07, 1.342111e-07, 1.342111e-07, 
    1.342109e-07, 1.342111e-07, 1.342108e-07, 1.34211e-07, 1.342109e-07, 
    1.342111e-07, 1.342118e-07, 1.342117e-07, 1.342118e-07, 1.342118e-07, 
    1.342118e-07, 1.342119e-07, 1.342119e-07, 1.342121e-07, 1.34212e-07, 
    1.34212e-07, 1.342118e-07, 1.342118e-07, 1.342117e-07, 1.342117e-07, 
    1.342115e-07, 1.342116e-07, 1.342113e-07, 1.342114e-07, 1.342111e-07, 
    1.342112e-07, 1.342111e-07, 1.342111e-07, 1.342111e-07, 1.342112e-07, 
    1.342112e-07, 1.342113e-07, 1.342116e-07, 1.342115e-07, 1.342117e-07, 
    1.342119e-07, 1.34212e-07, 1.342121e-07, 1.342121e-07, 1.342121e-07, 
    1.34212e-07, 1.342119e-07, 1.342118e-07, 1.342117e-07, 1.342117e-07, 
    1.342115e-07, 1.342114e-07, 1.342113e-07, 1.342113e-07, 1.342112e-07, 
    1.342112e-07, 1.342111e-07, 1.342111e-07, 1.342111e-07, 1.342112e-07, 
    1.342111e-07, 1.342113e-07, 1.342113e-07, 1.342117e-07, 1.342118e-07, 
    1.342119e-07, 1.342119e-07, 1.342121e-07, 1.34212e-07, 1.34212e-07, 
    1.342119e-07, 1.342119e-07, 1.342119e-07, 1.342117e-07, 1.342118e-07, 
    1.342114e-07, 1.342116e-07, 1.342112e-07, 1.342113e-07, 1.342112e-07, 
    1.342112e-07, 1.342111e-07, 1.342112e-07, 1.342111e-07, 1.34211e-07, 
    1.34211e-07, 1.34211e-07, 1.342112e-07, 1.342111e-07, 1.342119e-07, 
    1.342119e-07, 1.342119e-07, 1.34212e-07, 1.34212e-07, 1.342121e-07, 
    1.34212e-07, 1.34212e-07, 1.342119e-07, 1.342118e-07, 1.342118e-07, 
    1.342117e-07, 1.342116e-07, 1.342114e-07, 1.342113e-07, 1.342112e-07, 
    1.342113e-07, 1.342112e-07, 1.342113e-07, 1.342113e-07, 1.34211e-07, 
    1.342112e-07, 1.34211e-07, 1.34211e-07, 1.342111e-07, 1.34211e-07, 
    1.342119e-07, 1.342119e-07, 1.34212e-07, 1.342119e-07, 1.342121e-07, 
    1.34212e-07, 1.34212e-07, 1.342118e-07, 1.342118e-07, 1.342117e-07, 
    1.342117e-07, 1.342116e-07, 1.342114e-07, 1.342113e-07, 1.342112e-07, 
    1.342112e-07, 1.342112e-07, 1.342112e-07, 1.342112e-07, 1.342112e-07, 
    1.342111e-07, 1.342112e-07, 1.34211e-07, 1.34211e-07, 1.34211e-07, 
    1.34211e-07, 1.342119e-07, 1.342119e-07, 1.342119e-07, 1.342118e-07, 
    1.342119e-07, 1.342117e-07, 1.342117e-07, 1.342115e-07, 1.342116e-07, 
    1.342114e-07, 1.342116e-07, 1.342115e-07, 1.342114e-07, 1.342116e-07, 
    1.342113e-07, 1.342115e-07, 1.342112e-07, 1.342113e-07, 1.342111e-07, 
    1.342112e-07, 1.342111e-07, 1.342111e-07, 1.34211e-07, 1.342109e-07, 
    1.342109e-07, 1.342109e-07, 1.342118e-07, 1.342117e-07, 1.342117e-07, 
    1.342117e-07, 1.342116e-07, 1.342115e-07, 1.342114e-07, 1.342114e-07, 
    1.342113e-07, 1.342113e-07, 1.342115e-07, 1.342114e-07, 1.342117e-07, 
    1.342117e-07, 1.342117e-07, 1.342118e-07, 1.342114e-07, 1.342116e-07, 
    1.342113e-07, 1.342114e-07, 1.342111e-07, 1.342112e-07, 1.342109e-07, 
    1.342108e-07, 1.342107e-07, 1.342106e-07, 1.342117e-07, 1.342117e-07, 
    1.342117e-07, 1.342116e-07, 1.342115e-07, 1.342114e-07, 1.342114e-07, 
    1.342113e-07, 1.342113e-07, 1.342112e-07, 1.342113e-07, 1.342112e-07, 
    1.342116e-07, 1.342114e-07, 1.342118e-07, 1.342117e-07, 1.342116e-07, 
    1.342116e-07, 1.342115e-07, 1.342114e-07, 1.342113e-07, 1.342113e-07, 
    1.342109e-07, 1.342111e-07, 1.342105e-07, 1.342107e-07, 1.342118e-07, 
    1.342117e-07, 1.342115e-07, 1.342116e-07, 1.342114e-07, 1.342113e-07, 
    1.342113e-07, 1.342112e-07, 1.342112e-07, 1.342111e-07, 1.342112e-07, 
    1.342111e-07, 1.342114e-07, 1.342113e-07, 1.342115e-07, 1.342115e-07, 
    1.342115e-07, 1.342115e-07, 1.342114e-07, 1.342113e-07, 1.342113e-07, 
    1.342113e-07, 1.342112e-07, 1.342114e-07, 1.342108e-07, 1.342112e-07, 
    1.342117e-07, 1.342116e-07, 1.342115e-07, 1.342116e-07, 1.342113e-07, 
    1.342114e-07, 1.342111e-07, 1.342112e-07, 1.342111e-07, 1.342112e-07, 
    1.342112e-07, 1.342112e-07, 1.342113e-07, 1.342114e-07, 1.342115e-07, 
    1.342116e-07, 1.342116e-07, 1.342115e-07, 1.342113e-07, 1.342112e-07, 
    1.342112e-07, 1.342111e-07, 1.342114e-07, 1.342113e-07, 1.342113e-07, 
    1.342112e-07, 1.342114e-07, 1.342112e-07, 1.342115e-07, 1.342115e-07, 
    1.342114e-07, 1.342113e-07, 1.342112e-07, 1.342112e-07, 1.342112e-07, 
    1.342113e-07, 1.342113e-07, 1.342114e-07, 1.342114e-07, 1.342115e-07, 
    1.342115e-07, 1.342115e-07, 1.342114e-07, 1.342113e-07, 1.342112e-07, 
    1.342111e-07, 1.34211e-07, 1.342109e-07, 1.34211e-07, 1.342108e-07, 
    1.34211e-07, 1.342107e-07, 1.342112e-07, 1.34211e-07, 1.342114e-07, 
    1.342114e-07, 1.342113e-07, 1.342111e-07, 1.342112e-07, 1.342111e-07, 
    1.342113e-07, 1.342115e-07, 1.342115e-07, 1.342116e-07, 1.342115e-07, 
    1.342115e-07, 1.342114e-07, 1.342115e-07, 1.342113e-07, 1.342114e-07, 
    1.342112e-07, 1.342111e-07, 1.342109e-07, 1.342107e-07, 1.342106e-07, 
    1.342105e-07, 1.342105e-07, 1.342105e-07 ;

 LITR3N_TNDNCY_VERT_TRANS =
  7.352717e-27, -1.838179e-26, -4.901811e-26, -2.450905e-26, 9.190896e-26, 
    -1.237707e-25, 3.553813e-26, -5.514538e-26, -8.700715e-26, 6.862535e-26, 
    9.190896e-26, 1.139671e-25, -5.146902e-26, 3.798904e-26, -3.676358e-26, 
    6.862535e-26, -3.921449e-26, 1.936215e-25, 9.803622e-27, 1.017126e-25, 
    1.274471e-25, -5.637083e-26, 5.269447e-26, -2.941087e-26, -5.759628e-26, 
    1.347998e-26, 1.139671e-25, -3.308722e-26, -7.352717e-27, -4.779266e-26, 
    2.450905e-26, -1.225453e-27, 7.230172e-26, -9.926167e-26, 1.960724e-26, 
    8.333079e-26, -2.450906e-27, 1.188689e-25, 1.556325e-25, 6.73999e-26, 
    7.107626e-26, 4.65672e-26, 1.397016e-25, -2.941087e-26, 5.514538e-26, 
    3.676358e-26, 1.017126e-25, -4.901811e-27, 6.249809e-26, 5.514538e-26, 
    -5.146902e-26, -2.941087e-26, 6.127264e-27, -1.470543e-26, 1.02938e-25, 
    9.190896e-26, -4.289085e-26, -3.063632e-26, -9.803622e-27, -1.090653e-25, 
    1.102908e-26, -2.941087e-26, -8.455624e-26, 5.759628e-26, 6.98508e-26, 
    -1.176435e-25, -3.553813e-26, -1.017126e-25, -3.676358e-27, 
    -6.249809e-26, 6.73999e-26, -1.188689e-25, -5.391992e-26, 1.066144e-25, 
    3.798904e-26, -9.681077e-26, 1.139671e-25, -4.41163e-26, 5.759628e-26, 
    3.308722e-26, -3.186177e-26, 5.024356e-26, -1.176435e-25, 1.115162e-25, 
    4.043994e-26, 4.043994e-26, 3.063632e-26, 7.965443e-26, -6.4949e-26, 
    -7.720352e-26, 5.882173e-26, -4.901811e-27, 4.779266e-26, -3.308722e-26, 
    6.004719e-26, 2.08327e-26, 2.32836e-26, -4.779266e-26, 6.98508e-26, 
    1.225453e-26, -1.887197e-25, 2.450906e-27, -1.397016e-25, -4.41163e-26, 
    5.514538e-26, 1.090653e-25, -3.798904e-26, -2.450905e-26, -2.818541e-26, 
    -8.578169e-27, 8.087988e-26, 1.249962e-25, 5.759628e-26, -4.289085e-26, 
    6.127264e-26, 7.597807e-26, 1.02938e-25, 9.068351e-26, 1.078398e-25, 
    2.941087e-26, 9.190896e-26, -1.053889e-25, 1.188689e-25, -3.063632e-26, 
    -9.681077e-26, -1.67887e-25, 3.676358e-26, 4.901811e-27, 1.470543e-26, 
    7.107626e-26, -5.882173e-26, -4.043994e-26, -6.4949e-26, -1.985233e-25, 
    6.98508e-26, -7.475262e-26, -1.102908e-25, 8.945805e-26, -9.803622e-26, 
    -7.107626e-26, -1.593089e-26, 7.352717e-27, -1.225453e-27, -5.637083e-26, 
    6.862535e-26, -5.759628e-26, 3.676358e-27, 4.043994e-26, 4.779266e-26, 
    -1.703379e-25, 5.024356e-26, -1.225453e-27, -4.779266e-26, -1.838179e-26, 
    3.921449e-26, 4.779266e-26, 7.965443e-26, -1.838179e-26, 8.945805e-26, 
    -3.308722e-26, -7.475262e-26, -1.225453e-26, -3.676358e-26, -4.41163e-26, 
    -6.004719e-26, 2.450906e-27, -1.960724e-26, 6.98508e-26, -4.534175e-26, 
    1.225453e-27, -8.210533e-26, -4.41163e-26, 1.225453e-27, -2.573451e-26, 
    -7.352717e-27, 8.578169e-27, 2.32836e-26, -2.450905e-26, 1.715634e-26, 
    -1.188689e-25, -5.146902e-26, -6.127264e-26, -1.347998e-25, 
    -1.188689e-25, -1.115162e-25, 7.842898e-26, -5.269447e-26, -9.803622e-27, 
    9.313441e-26, 2.205815e-26, 1.629852e-25, 2.450906e-27, 1.102908e-26, 
    -6.249809e-26, 4.901811e-26, 4.901811e-26, 1.213198e-25, -2.450906e-27, 
    -1.225453e-27, 2.205815e-26, -3.676358e-26, 2.08327e-26, -9.803622e-27, 
    -1.347998e-26, 9.926167e-26, 2.695996e-26, -3.063632e-26, -1.139671e-25, 
    4.779266e-26, -3.921449e-26, 5.514538e-26, -3.553813e-26, -5.269447e-26, 
    -3.676358e-27, 4.166539e-26, 3.921449e-26, 1.360253e-25, -1.531816e-25, 
    4.901811e-27, 9.803622e-27, -1.715634e-26, 1.838179e-26, 5.637083e-26, 
    3.676358e-27, -1.053889e-25, -1.02938e-25, -5.146902e-26, 4.901811e-27, 
    2.695996e-26, 8.333079e-26, -5.024356e-26, -7.475262e-26, 1.02938e-25, 
    -1.102908e-26, -1.470543e-26, 5.391992e-26, -7.842898e-26, -5.391992e-26, 
    1.960724e-26, 2.450906e-27, 1.225453e-27, -3.798904e-26, -3.186177e-26, 
    2.941087e-26, -4.043994e-26, 8.210533e-26, 1.02938e-25, -5.882173e-26, 
    -6.127264e-27, -1.102908e-26, -9.803622e-27, 2.450905e-26, -3.308722e-26, 
    -2.450905e-26, -8.455624e-26, -6.862535e-26, -9.803622e-26, 7.107626e-26, 
    4.901811e-27, -6.4949e-26, -6.372354e-26, 1.347998e-25, 3.676358e-26, 
    4.534175e-26, -9.803622e-26, -4.901811e-26, 3.798904e-26, 5.146902e-26, 
    1.43378e-25, 1.188689e-25, -5.759628e-26, -1.066144e-25, -2.450905e-26, 
    1.593089e-26, 3.186177e-26, -5.514538e-26, -8.210533e-26, 8.945805e-26, 
    -6.127264e-27, 9.681077e-26, -4.41163e-26, -3.676358e-27, 9.803622e-26, 
    2.32836e-26, 3.308722e-26, -6.249809e-26, 6.4949e-26, 3.921449e-26, 
    4.289085e-26, -7.230172e-26, 1.593089e-25, 2.450906e-27, 6.004719e-26, 
    -4.901811e-27, 8.578169e-26, 3.186177e-26, 1.29898e-25, -2.08327e-26, 
    2.695996e-26, 1.225453e-26, -5.514538e-26, -1.593089e-26, -2.450906e-27, 
    4.901811e-27, -1.29898e-25, -1.225453e-26, -1.004871e-25, -1.384762e-25, 
    5.269447e-26, -2.450906e-27, 1.593089e-26, -8.210533e-26, 9.803622e-27, 
    4.289085e-26, -2.32836e-26, -1.81367e-25, 6.127264e-27, 3.676358e-27, 
    5.882173e-26, -4.901811e-27, 6.98508e-26, -1.102908e-26, 3.186177e-26, 
    -8.578169e-27, 1.347998e-26, -3.676358e-26, -1.213198e-25, 3.553813e-26, 
    -1.02938e-25, 5.146902e-26, 1.262216e-25, -8.578169e-26, -8.945805e-26, 
    1.960724e-26, 3.431268e-26, -9.681077e-26, 2.818541e-26, 1.017126e-25,
  1.338114e-32, 1.338112e-32, 1.338113e-32, 1.338111e-32, 1.338112e-32, 
    1.338111e-32, 1.338113e-32, 1.338112e-32, 1.338113e-32, 1.338113e-32, 
    1.338109e-32, 1.338111e-32, 1.338107e-32, 1.338109e-32, 1.338105e-32, 
    1.338107e-32, 1.338105e-32, 1.338105e-32, 1.338104e-32, 1.338104e-32, 
    1.338102e-32, 1.338104e-32, 1.338101e-32, 1.338103e-32, 1.338102e-32, 
    1.338104e-32, 1.338111e-32, 1.33811e-32, 1.338111e-32, 1.338111e-32, 
    1.338111e-32, 1.338112e-32, 1.338113e-32, 1.338114e-32, 1.338113e-32, 
    1.338113e-32, 1.338111e-32, 1.338111e-32, 1.33811e-32, 1.33811e-32, 
    1.338108e-32, 1.338109e-32, 1.338106e-32, 1.338107e-32, 1.338104e-32, 
    1.338105e-32, 1.338104e-32, 1.338104e-32, 1.338104e-32, 1.338105e-32, 
    1.338105e-32, 1.338106e-32, 1.338109e-32, 1.338108e-32, 1.33811e-32, 
    1.338112e-32, 1.338113e-32, 1.338114e-32, 1.338114e-32, 1.338114e-32, 
    1.338113e-32, 1.338112e-32, 1.338111e-32, 1.33811e-32, 1.33811e-32, 
    1.338108e-32, 1.338108e-32, 1.338106e-32, 1.338106e-32, 1.338105e-32, 
    1.338105e-32, 1.338104e-32, 1.338104e-32, 1.338104e-32, 1.338105e-32, 
    1.338104e-32, 1.338106e-32, 1.338106e-32, 1.33811e-32, 1.338111e-32, 
    1.338112e-32, 1.338112e-32, 1.338114e-32, 1.338113e-32, 1.338113e-32, 
    1.338112e-32, 1.338112e-32, 1.338112e-32, 1.33811e-32, 1.338111e-32, 
    1.338107e-32, 1.338109e-32, 1.338105e-32, 1.338106e-32, 1.338105e-32, 
    1.338105e-32, 1.338104e-32, 1.338105e-32, 1.338104e-32, 1.338103e-32, 
    1.338104e-32, 1.338103e-32, 1.338105e-32, 1.338104e-32, 1.338112e-32, 
    1.338112e-32, 1.338112e-32, 1.338113e-32, 1.338113e-32, 1.338114e-32, 
    1.338113e-32, 1.338113e-32, 1.338112e-32, 1.338111e-32, 1.338111e-32, 
    1.33811e-32, 1.338109e-32, 1.338107e-32, 1.338106e-32, 1.338105e-32, 
    1.338106e-32, 1.338105e-32, 1.338106e-32, 1.338106e-32, 1.338103e-32, 
    1.338105e-32, 1.338103e-32, 1.338103e-32, 1.338104e-32, 1.338103e-32, 
    1.338112e-32, 1.338112e-32, 1.338113e-32, 1.338113e-32, 1.338114e-32, 
    1.338113e-32, 1.338113e-32, 1.338111e-32, 1.338111e-32, 1.33811e-32, 
    1.33811e-32, 1.338109e-32, 1.338107e-32, 1.338106e-32, 1.338105e-32, 
    1.338105e-32, 1.338105e-32, 1.338105e-32, 1.338105e-32, 1.338105e-32, 
    1.338104e-32, 1.338105e-32, 1.338103e-32, 1.338103e-32, 1.338103e-32, 
    1.338103e-32, 1.338112e-32, 1.338112e-32, 1.338112e-32, 1.338112e-32, 
    1.338112e-32, 1.33811e-32, 1.33811e-32, 1.338108e-32, 1.338109e-32, 
    1.338108e-32, 1.338109e-32, 1.338108e-32, 1.338108e-32, 1.338109e-32, 
    1.338106e-32, 1.338108e-32, 1.338105e-32, 1.338106e-32, 1.338105e-32, 
    1.338105e-32, 1.338104e-32, 1.338104e-32, 1.338103e-32, 1.338102e-32, 
    1.338102e-32, 1.338102e-32, 1.338111e-32, 1.33811e-32, 1.33811e-32, 
    1.33811e-32, 1.338109e-32, 1.338109e-32, 1.338107e-32, 1.338108e-32, 
    1.338107e-32, 1.338106e-32, 1.338108e-32, 1.338107e-32, 1.33811e-32, 
    1.33811e-32, 1.33811e-32, 1.338111e-32, 1.338107e-32, 1.338109e-32, 
    1.338106e-32, 1.338107e-32, 1.338104e-32, 1.338105e-32, 1.338103e-32, 
    1.338101e-32, 1.3381e-32, 1.338099e-32, 1.33811e-32, 1.338111e-32, 
    1.33811e-32, 1.338109e-32, 1.338108e-32, 1.338107e-32, 1.338107e-32, 
    1.338107e-32, 1.338106e-32, 1.338105e-32, 1.338106e-32, 1.338105e-32, 
    1.338109e-32, 1.338107e-32, 1.338111e-32, 1.33811e-32, 1.338109e-32, 
    1.338109e-32, 1.338108e-32, 1.338107e-32, 1.338106e-32, 1.338107e-32, 
    1.338102e-32, 1.338104e-32, 1.338098e-32, 1.338099e-32, 1.338111e-32, 
    1.33811e-32, 1.338108e-32, 1.338109e-32, 1.338107e-32, 1.338106e-32, 
    1.338106e-32, 1.338105e-32, 1.338105e-32, 1.338104e-32, 1.338105e-32, 
    1.338105e-32, 1.338107e-32, 1.338106e-32, 1.338109e-32, 1.338108e-32, 
    1.338108e-32, 1.338109e-32, 1.338108e-32, 1.338106e-32, 1.338106e-32, 
    1.338106e-32, 1.338105e-32, 1.338107e-32, 1.338101e-32, 1.338105e-32, 
    1.33811e-32, 1.338109e-32, 1.338108e-32, 1.338109e-32, 1.338106e-32, 
    1.338107e-32, 1.338104e-32, 1.338105e-32, 1.338104e-32, 1.338105e-32, 
    1.338105e-32, 1.338105e-32, 1.338106e-32, 1.338107e-32, 1.338108e-32, 
    1.338109e-32, 1.338109e-32, 1.338108e-32, 1.338106e-32, 1.338105e-32, 
    1.338105e-32, 1.338104e-32, 1.338107e-32, 1.338106e-32, 1.338106e-32, 
    1.338105e-32, 1.338108e-32, 1.338105e-32, 1.338108e-32, 1.338108e-32, 
    1.338107e-32, 1.338106e-32, 1.338105e-32, 1.338105e-32, 1.338105e-32, 
    1.338106e-32, 1.338106e-32, 1.338107e-32, 1.338107e-32, 1.338108e-32, 
    1.338108e-32, 1.338108e-32, 1.338108e-32, 1.338106e-32, 1.338105e-32, 
    1.338104e-32, 1.338104e-32, 1.338102e-32, 1.338103e-32, 1.338101e-32, 
    1.338103e-32, 1.3381e-32, 1.338105e-32, 1.338103e-32, 1.338107e-32, 
    1.338107e-32, 1.338106e-32, 1.338104e-32, 1.338105e-32, 1.338104e-32, 
    1.338106e-32, 1.338108e-32, 1.338108e-32, 1.338109e-32, 1.338108e-32, 
    1.338108e-32, 1.338108e-32, 1.338108e-32, 1.338106e-32, 1.338107e-32, 
    1.338105e-32, 1.338104e-32, 1.338102e-32, 1.3381e-32, 1.338099e-32, 
    1.338098e-32, 1.338098e-32, 1.338098e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N_TO_SOIL2N =
  1.70703e-15, 1.711376e-15, 1.710532e-15, 1.714033e-15, 1.712092e-15, 
    1.714383e-15, 1.707912e-15, 1.711547e-15, 1.709228e-15, 1.707423e-15, 
    1.720817e-15, 1.714189e-15, 1.727695e-15, 1.723476e-15, 1.734066e-15, 
    1.727038e-15, 1.735482e-15, 1.733865e-15, 1.738733e-15, 1.737339e-15, 
    1.743555e-15, 1.739376e-15, 1.746775e-15, 1.742558e-15, 1.743218e-15, 
    1.739238e-15, 1.715525e-15, 1.719992e-15, 1.71526e-15, 1.715898e-15, 
    1.715612e-15, 1.712131e-15, 1.710375e-15, 1.706699e-15, 1.707367e-15, 
    1.710067e-15, 1.716184e-15, 1.71411e-15, 1.719338e-15, 1.719221e-15, 
    1.725032e-15, 1.722413e-15, 1.732168e-15, 1.729399e-15, 1.737397e-15, 
    1.735387e-15, 1.737303e-15, 1.736722e-15, 1.73731e-15, 1.734362e-15, 
    1.735625e-15, 1.73303e-15, 1.722903e-15, 1.725882e-15, 1.71699e-15, 
    1.711631e-15, 1.708072e-15, 1.705542e-15, 1.7059e-15, 1.706582e-15, 
    1.710083e-15, 1.713374e-15, 1.715879e-15, 1.717554e-15, 1.719204e-15, 
    1.724189e-15, 1.726828e-15, 1.732727e-15, 1.731665e-15, 1.733466e-15, 
    1.735187e-15, 1.738074e-15, 1.737599e-15, 1.73887e-15, 1.733419e-15, 
    1.737042e-15, 1.731059e-15, 1.732696e-15, 1.719647e-15, 1.71467e-15, 
    1.712548e-15, 1.710694e-15, 1.706175e-15, 1.709296e-15, 1.708066e-15, 
    1.710993e-15, 1.712851e-15, 1.711932e-15, 1.7176e-15, 1.715397e-15, 
    1.726984e-15, 1.721998e-15, 1.734986e-15, 1.731883e-15, 1.73573e-15, 
    1.733768e-15, 1.737129e-15, 1.734104e-15, 1.739344e-15, 1.740483e-15, 
    1.739704e-15, 1.742696e-15, 1.733936e-15, 1.737302e-15, 1.711906e-15, 
    1.712056e-15, 1.712754e-15, 1.709683e-15, 1.709495e-15, 1.706681e-15, 
    1.709186e-15, 1.710252e-15, 1.712959e-15, 1.714558e-15, 1.716078e-15, 
    1.719418e-15, 1.723143e-15, 1.728348e-15, 1.732084e-15, 1.734586e-15, 
    1.733052e-15, 1.734406e-15, 1.732892e-15, 1.732183e-15, 1.740056e-15, 
    1.735637e-15, 1.742266e-15, 1.7419e-15, 1.7389e-15, 1.741941e-15, 
    1.712161e-15, 1.711299e-15, 1.708302e-15, 1.710648e-15, 1.706374e-15, 
    1.708766e-15, 1.71014e-15, 1.715442e-15, 1.716607e-15, 1.717685e-15, 
    1.719816e-15, 1.722547e-15, 1.727333e-15, 1.731493e-15, 1.735288e-15, 
    1.73501e-15, 1.735108e-15, 1.735954e-15, 1.733856e-15, 1.736299e-15, 
    1.736708e-15, 1.735637e-15, 1.741851e-15, 1.740077e-15, 1.741892e-15, 
    1.740737e-15, 1.711579e-15, 1.71303e-15, 1.712246e-15, 1.71372e-15, 
    1.712681e-15, 1.717296e-15, 1.718679e-15, 1.725143e-15, 1.722493e-15, 
    1.726711e-15, 1.722922e-15, 1.723593e-15, 1.726847e-15, 1.723127e-15, 
    1.731263e-15, 1.725747e-15, 1.735987e-15, 1.730484e-15, 1.736332e-15, 
    1.735271e-15, 1.737027e-15, 1.738598e-15, 1.740575e-15, 1.744218e-15, 
    1.743375e-15, 1.74642e-15, 1.715193e-15, 1.717072e-15, 1.716908e-15, 
    1.718874e-15, 1.720328e-15, 1.723478e-15, 1.728523e-15, 1.726627e-15, 
    1.730108e-15, 1.730806e-15, 1.725518e-15, 1.728765e-15, 1.71833e-15, 
    1.720017e-15, 1.719014e-15, 1.71534e-15, 1.727063e-15, 1.721051e-15, 
    1.732146e-15, 1.728895e-15, 1.738374e-15, 1.733662e-15, 1.742911e-15, 
    1.746854e-15, 1.750566e-15, 1.754894e-15, 1.718099e-15, 1.716822e-15, 
    1.719109e-15, 1.722268e-15, 1.7252e-15, 1.729093e-15, 1.729491e-15, 
    1.73022e-15, 1.732107e-15, 1.733693e-15, 1.730449e-15, 1.73409e-15, 
    1.720406e-15, 1.727585e-15, 1.716338e-15, 1.719727e-15, 1.722082e-15, 
    1.72105e-15, 1.726411e-15, 1.727672e-15, 1.732795e-15, 1.730149e-15, 
    1.74588e-15, 1.738929e-15, 1.758189e-15, 1.752817e-15, 1.716375e-15, 
    1.718095e-15, 1.724071e-15, 1.721229e-15, 1.729353e-15, 1.73135e-15, 
    1.732973e-15, 1.735045e-15, 1.735269e-15, 1.736497e-15, 1.734485e-15, 
    1.736418e-15, 1.729101e-15, 1.732373e-15, 1.723389e-15, 1.725577e-15, 
    1.724571e-15, 1.723467e-15, 1.726875e-15, 1.7305e-15, 1.730579e-15, 
    1.731741e-15, 1.735009e-15, 1.729386e-15, 1.746774e-15, 1.736043e-15, 
    1.719968e-15, 1.723274e-15, 1.723748e-15, 1.722467e-15, 1.73115e-15, 
    1.728006e-15, 1.736467e-15, 1.734183e-15, 1.737925e-15, 1.736066e-15, 
    1.735792e-15, 1.733403e-15, 1.731914e-15, 1.72815e-15, 1.725085e-15, 
    1.722653e-15, 1.723219e-15, 1.725889e-15, 1.730722e-15, 1.735289e-15, 
    1.734289e-15, 1.737641e-15, 1.728765e-15, 1.732488e-15, 1.731049e-15, 
    1.734801e-15, 1.726576e-15, 1.733576e-15, 1.724784e-15, 1.725556e-15, 
    1.727944e-15, 1.73274e-15, 1.733802e-15, 1.734934e-15, 1.734236e-15, 
    1.730845e-15, 1.73029e-15, 1.727886e-15, 1.727221e-15, 1.725388e-15, 
    1.72387e-15, 1.725257e-15, 1.726713e-15, 1.730847e-15, 1.734568e-15, 
    1.73862e-15, 1.739612e-15, 1.744336e-15, 1.740489e-15, 1.746833e-15, 
    1.741437e-15, 1.750774e-15, 1.733984e-15, 1.741281e-15, 1.728053e-15, 
    1.72948e-15, 1.73206e-15, 1.737973e-15, 1.734784e-15, 1.738514e-15, 
    1.730268e-15, 1.725981e-15, 1.724873e-15, 1.722801e-15, 1.72492e-15, 
    1.724748e-15, 1.726774e-15, 1.726123e-15, 1.730984e-15, 1.728374e-15, 
    1.735785e-15, 1.738485e-15, 1.746101e-15, 1.75076e-15, 1.755499e-15, 
    1.757588e-15, 1.758224e-15, 1.75849e-15 ;

 LITR3N_vr =
  7.663647e-06, 7.663639e-06, 7.663641e-06, 7.663634e-06, 7.663638e-06, 
    7.663634e-06, 7.663645e-06, 7.663639e-06, 7.663643e-06, 7.663646e-06, 
    7.663622e-06, 7.663634e-06, 7.663611e-06, 7.663618e-06, 7.6636e-06, 
    7.663612e-06, 7.663597e-06, 7.6636e-06, 7.663592e-06, 7.663594e-06, 
    7.663583e-06, 7.663591e-06, 7.663577e-06, 7.663585e-06, 7.663583e-06, 
    7.663591e-06, 7.663632e-06, 7.663624e-06, 7.663632e-06, 7.663632e-06, 
    7.663632e-06, 7.663638e-06, 7.663641e-06, 7.663647e-06, 7.663646e-06, 
    7.663642e-06, 7.663631e-06, 7.663634e-06, 7.663625e-06, 7.663625e-06, 
    7.663615e-06, 7.66362e-06, 7.663603e-06, 7.663608e-06, 7.663593e-06, 
    7.663597e-06, 7.663594e-06, 7.663595e-06, 7.663594e-06, 7.663599e-06, 
    7.663597e-06, 7.663602e-06, 7.663619e-06, 7.663614e-06, 7.66363e-06, 
    7.663639e-06, 7.663645e-06, 7.66365e-06, 7.663649e-06, 7.663648e-06, 
    7.663642e-06, 7.663636e-06, 7.663632e-06, 7.663629e-06, 7.663625e-06, 
    7.663617e-06, 7.663612e-06, 7.663602e-06, 7.663604e-06, 7.663601e-06, 
    7.663598e-06, 7.663592e-06, 7.663593e-06, 7.663592e-06, 7.663601e-06, 
    7.663594e-06, 7.663605e-06, 7.663602e-06, 7.663625e-06, 7.663633e-06, 
    7.663637e-06, 7.663641e-06, 7.663648e-06, 7.663642e-06, 7.663645e-06, 
    7.66364e-06, 7.663637e-06, 7.663638e-06, 7.663629e-06, 7.663632e-06, 
    7.663612e-06, 7.663621e-06, 7.663598e-06, 7.663603e-06, 7.663597e-06, 
    7.6636e-06, 7.663594e-06, 7.6636e-06, 7.663591e-06, 7.663589e-06, 
    7.66359e-06, 7.663584e-06, 7.6636e-06, 7.663594e-06, 7.663638e-06, 
    7.663638e-06, 7.663637e-06, 7.663642e-06, 7.663642e-06, 7.663647e-06, 
    7.663643e-06, 7.663642e-06, 7.663636e-06, 7.663633e-06, 7.663631e-06, 
    7.663625e-06, 7.663619e-06, 7.66361e-06, 7.663603e-06, 7.663599e-06, 
    7.663602e-06, 7.663599e-06, 7.663602e-06, 7.663603e-06, 7.663589e-06, 
    7.663597e-06, 7.663585e-06, 7.663586e-06, 7.663592e-06, 7.663586e-06, 
    7.663638e-06, 7.66364e-06, 7.663644e-06, 7.663641e-06, 7.663648e-06, 
    7.663643e-06, 7.663642e-06, 7.663632e-06, 7.66363e-06, 7.663628e-06, 
    7.663624e-06, 7.66362e-06, 7.663612e-06, 7.663604e-06, 7.663598e-06, 
    7.663598e-06, 7.663598e-06, 7.663596e-06, 7.6636e-06, 7.663596e-06, 
    7.663595e-06, 7.663597e-06, 7.663586e-06, 7.663589e-06, 7.663586e-06, 
    7.663588e-06, 7.663639e-06, 7.663636e-06, 7.663638e-06, 7.663635e-06, 
    7.663637e-06, 7.663629e-06, 7.663626e-06, 7.663615e-06, 7.66362e-06, 
    7.663612e-06, 7.663619e-06, 7.663618e-06, 7.663612e-06, 7.663619e-06, 
    7.663604e-06, 7.663614e-06, 7.663596e-06, 7.663606e-06, 7.663596e-06, 
    7.663598e-06, 7.663594e-06, 7.663592e-06, 7.663588e-06, 7.663582e-06, 
    7.663583e-06, 7.663578e-06, 7.663632e-06, 7.66363e-06, 7.66363e-06, 
    7.663626e-06, 7.663623e-06, 7.663618e-06, 7.66361e-06, 7.663612e-06, 
    7.663606e-06, 7.663605e-06, 7.663614e-06, 7.663609e-06, 7.663627e-06, 
    7.663624e-06, 7.663626e-06, 7.663632e-06, 7.663612e-06, 7.663622e-06, 
    7.663603e-06, 7.663609e-06, 7.663592e-06, 7.663601e-06, 7.663584e-06, 
    7.663577e-06, 7.663571e-06, 7.663563e-06, 7.663628e-06, 7.66363e-06, 
    7.663626e-06, 7.663621e-06, 7.663615e-06, 7.663608e-06, 7.663608e-06, 
    7.663606e-06, 7.663603e-06, 7.663601e-06, 7.663606e-06, 7.6636e-06, 
    7.663623e-06, 7.663611e-06, 7.663631e-06, 7.663624e-06, 7.663621e-06, 
    7.663622e-06, 7.663613e-06, 7.663611e-06, 7.663602e-06, 7.663606e-06, 
    7.663579e-06, 7.663592e-06, 7.663558e-06, 7.663567e-06, 7.663631e-06, 
    7.663628e-06, 7.663617e-06, 7.663622e-06, 7.663608e-06, 7.663604e-06, 
    7.663602e-06, 7.663598e-06, 7.663598e-06, 7.663595e-06, 7.663599e-06, 
    7.663595e-06, 7.663608e-06, 7.663602e-06, 7.663618e-06, 7.663614e-06, 
    7.663616e-06, 7.663618e-06, 7.663612e-06, 7.663606e-06, 7.663606e-06, 
    7.663603e-06, 7.663598e-06, 7.663608e-06, 7.663577e-06, 7.663596e-06, 
    7.663624e-06, 7.663619e-06, 7.663618e-06, 7.66362e-06, 7.663604e-06, 
    7.663611e-06, 7.663595e-06, 7.6636e-06, 7.663592e-06, 7.663596e-06, 
    7.663597e-06, 7.663601e-06, 7.663603e-06, 7.66361e-06, 7.663615e-06, 
    7.66362e-06, 7.663619e-06, 7.663614e-06, 7.663605e-06, 7.663598e-06, 
    7.663599e-06, 7.663593e-06, 7.663609e-06, 7.663602e-06, 7.663605e-06, 
    7.663598e-06, 7.663612e-06, 7.663601e-06, 7.663616e-06, 7.663614e-06, 
    7.663611e-06, 7.663602e-06, 7.6636e-06, 7.663598e-06, 7.6636e-06, 
    7.663605e-06, 7.663606e-06, 7.663611e-06, 7.663612e-06, 7.663615e-06, 
    7.663617e-06, 7.663615e-06, 7.663612e-06, 7.663605e-06, 7.663599e-06, 
    7.663592e-06, 7.66359e-06, 7.663582e-06, 7.663589e-06, 7.663577e-06, 
    7.663587e-06, 7.663571e-06, 7.6636e-06, 7.663587e-06, 7.66361e-06, 
    7.663608e-06, 7.663603e-06, 7.663592e-06, 7.663599e-06, 7.663592e-06, 
    7.663606e-06, 7.663613e-06, 7.663616e-06, 7.66362e-06, 7.663615e-06, 
    7.663616e-06, 7.663612e-06, 7.663613e-06, 7.663605e-06, 7.66361e-06, 
    7.663597e-06, 7.663592e-06, 7.663579e-06, 7.663571e-06, 7.663562e-06, 
    7.663559e-06, 7.663557e-06, 7.663557e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3_HR =
  6.167343e-14, 6.183042e-14, 6.179994e-14, 6.192643e-14, 6.18563e-14, 
    6.193909e-14, 6.17053e-14, 6.183664e-14, 6.175282e-14, 6.168761e-14, 
    6.217151e-14, 6.193208e-14, 6.242002e-14, 6.226761e-14, 6.265021e-14, 
    6.239628e-14, 6.270136e-14, 6.264295e-14, 6.281882e-14, 6.276846e-14, 
    6.299303e-14, 6.284206e-14, 6.310938e-14, 6.295702e-14, 6.298084e-14, 
    6.283706e-14, 6.198036e-14, 6.214171e-14, 6.197077e-14, 6.19938e-14, 
    6.198348e-14, 6.185773e-14, 6.179427e-14, 6.166146e-14, 6.168559e-14, 
    6.178315e-14, 6.200415e-14, 6.192921e-14, 6.211812e-14, 6.211385e-14, 
    6.232382e-14, 6.222919e-14, 6.258164e-14, 6.248158e-14, 6.277057e-14, 
    6.269794e-14, 6.276715e-14, 6.274617e-14, 6.276742e-14, 6.26609e-14, 
    6.270654e-14, 6.261278e-14, 6.224691e-14, 6.235452e-14, 6.203327e-14, 
    6.183966e-14, 6.171105e-14, 6.161968e-14, 6.16326e-14, 6.165722e-14, 
    6.178372e-14, 6.190261e-14, 6.199314e-14, 6.205364e-14, 6.211324e-14, 
    6.229334e-14, 6.238869e-14, 6.260183e-14, 6.256345e-14, 6.262851e-14, 
    6.269072e-14, 6.279502e-14, 6.277786e-14, 6.282378e-14, 6.262683e-14, 
    6.275774e-14, 6.254156e-14, 6.260072e-14, 6.212924e-14, 6.194944e-14, 
    6.187278e-14, 6.180579e-14, 6.164253e-14, 6.175528e-14, 6.171084e-14, 
    6.181659e-14, 6.188371e-14, 6.185053e-14, 6.205529e-14, 6.197571e-14, 
    6.239434e-14, 6.221418e-14, 6.268346e-14, 6.257133e-14, 6.271033e-14, 
    6.263943e-14, 6.276088e-14, 6.265158e-14, 6.284089e-14, 6.288205e-14, 
    6.285392e-14, 6.296201e-14, 6.264551e-14, 6.276713e-14, 6.184959e-14, 
    6.1855e-14, 6.188023e-14, 6.176927e-14, 6.17625e-14, 6.166079e-14, 
    6.175131e-14, 6.178982e-14, 6.188762e-14, 6.19454e-14, 6.200031e-14, 
    6.212098e-14, 6.225558e-14, 6.244363e-14, 6.25786e-14, 6.266898e-14, 
    6.261358e-14, 6.266249e-14, 6.26078e-14, 6.258218e-14, 6.286661e-14, 
    6.270695e-14, 6.294646e-14, 6.293323e-14, 6.282487e-14, 6.293472e-14, 
    6.18588e-14, 6.182765e-14, 6.171937e-14, 6.180412e-14, 6.164971e-14, 
    6.173614e-14, 6.17858e-14, 6.197734e-14, 6.201943e-14, 6.205839e-14, 
    6.213535e-14, 6.223403e-14, 6.240695e-14, 6.255726e-14, 6.269434e-14, 
    6.268431e-14, 6.268784e-14, 6.271843e-14, 6.264262e-14, 6.273087e-14, 
    6.274565e-14, 6.270696e-14, 6.293146e-14, 6.286736e-14, 6.293295e-14, 
    6.289123e-14, 6.183778e-14, 6.18902e-14, 6.186188e-14, 6.191513e-14, 
    6.18776e-14, 6.204434e-14, 6.209428e-14, 6.232783e-14, 6.223208e-14, 
    6.238448e-14, 6.224758e-14, 6.227184e-14, 6.238938e-14, 6.2255e-14, 
    6.254894e-14, 6.234965e-14, 6.271961e-14, 6.25208e-14, 6.273206e-14, 
    6.269375e-14, 6.275719e-14, 6.281396e-14, 6.288537e-14, 6.301699e-14, 
    6.298653e-14, 6.309655e-14, 6.196833e-14, 6.203623e-14, 6.203029e-14, 
    6.210135e-14, 6.215386e-14, 6.226767e-14, 6.244995e-14, 6.238144e-14, 
    6.250722e-14, 6.253244e-14, 6.234137e-14, 6.245868e-14, 6.208169e-14, 
    6.214263e-14, 6.210637e-14, 6.197367e-14, 6.239718e-14, 6.217998e-14, 
    6.258082e-14, 6.246337e-14, 6.280586e-14, 6.263561e-14, 6.296976e-14, 
    6.311224e-14, 6.324635e-14, 6.34027e-14, 6.207332e-14, 6.202719e-14, 
    6.21098e-14, 6.222396e-14, 6.232989e-14, 6.247053e-14, 6.248493e-14, 
    6.251125e-14, 6.257944e-14, 6.263672e-14, 6.251954e-14, 6.265108e-14, 
    6.215669e-14, 6.241604e-14, 6.200972e-14, 6.213215e-14, 6.221725e-14, 
    6.217996e-14, 6.237362e-14, 6.241921e-14, 6.26043e-14, 6.250867e-14, 
    6.307705e-14, 6.282589e-14, 6.352174e-14, 6.332765e-14, 6.201106e-14, 
    6.207318e-14, 6.228908e-14, 6.21864e-14, 6.247993e-14, 6.255207e-14, 
    6.261071e-14, 6.268557e-14, 6.269368e-14, 6.273802e-14, 6.266535e-14, 
    6.273516e-14, 6.247083e-14, 6.258903e-14, 6.226446e-14, 6.234352e-14, 
    6.230717e-14, 6.226726e-14, 6.239038e-14, 6.252137e-14, 6.252422e-14, 
    6.256619e-14, 6.268426e-14, 6.248112e-14, 6.310932e-14, 6.272162e-14, 
    6.214087e-14, 6.22603e-14, 6.227742e-14, 6.223116e-14, 6.254483e-14, 
    6.243126e-14, 6.273695e-14, 6.265442e-14, 6.278963e-14, 6.272245e-14, 
    6.271256e-14, 6.262623e-14, 6.257244e-14, 6.243646e-14, 6.232572e-14, 
    6.223788e-14, 6.225832e-14, 6.235479e-14, 6.252939e-14, 6.269439e-14, 
    6.265825e-14, 6.277936e-14, 6.245867e-14, 6.259321e-14, 6.254121e-14, 
    6.267677e-14, 6.237961e-14, 6.263252e-14, 6.231487e-14, 6.234276e-14, 
    6.2429e-14, 6.260229e-14, 6.264068e-14, 6.268156e-14, 6.265635e-14, 
    6.253383e-14, 6.251378e-14, 6.242692e-14, 6.24029e-14, 6.233669e-14, 
    6.228182e-14, 6.233194e-14, 6.238455e-14, 6.253391e-14, 6.266834e-14, 
    6.281476e-14, 6.285058e-14, 6.302126e-14, 6.288226e-14, 6.311147e-14, 
    6.29165e-14, 6.325387e-14, 6.264725e-14, 6.291089e-14, 6.243295e-14, 
    6.248454e-14, 6.257773e-14, 6.279135e-14, 6.267613e-14, 6.281089e-14, 
    6.251299e-14, 6.235809e-14, 6.231806e-14, 6.224321e-14, 6.231977e-14, 
    6.231354e-14, 6.238676e-14, 6.236324e-14, 6.253886e-14, 6.244456e-14, 
    6.27123e-14, 6.280985e-14, 6.3085e-14, 6.325334e-14, 6.342457e-14, 
    6.350005e-14, 6.352302e-14, 6.353261e-14 ;

 LITTERC =
  5.976081e-05, 5.976067e-05, 5.97607e-05, 5.976058e-05, 5.976064e-05, 
    5.976057e-05, 5.976078e-05, 5.976066e-05, 5.976074e-05, 5.97608e-05, 
    5.976036e-05, 5.976058e-05, 5.976013e-05, 5.976027e-05, 5.975992e-05, 
    5.976015e-05, 5.975987e-05, 5.975992e-05, 5.975976e-05, 5.975981e-05, 
    5.97596e-05, 5.975974e-05, 5.97595e-05, 5.975964e-05, 5.975962e-05, 
    5.975975e-05, 5.976053e-05, 5.976038e-05, 5.976054e-05, 5.976052e-05, 
    5.976053e-05, 5.976064e-05, 5.97607e-05, 5.976082e-05, 5.97608e-05, 
    5.976071e-05, 5.976051e-05, 5.976058e-05, 5.97604e-05, 5.976041e-05, 
    5.976022e-05, 5.97603e-05, 5.975998e-05, 5.976007e-05, 5.975981e-05, 
    5.975987e-05, 5.975981e-05, 5.975983e-05, 5.975981e-05, 5.975991e-05, 
    5.975987e-05, 5.975995e-05, 5.976029e-05, 5.976019e-05, 5.976048e-05, 
    5.976066e-05, 5.976078e-05, 5.976086e-05, 5.976085e-05, 5.976083e-05, 
    5.976071e-05, 5.97606e-05, 5.976052e-05, 5.976046e-05, 5.976041e-05, 
    5.976024e-05, 5.976016e-05, 5.975996e-05, 5.976e-05, 5.975994e-05, 
    5.975988e-05, 5.975979e-05, 5.97598e-05, 5.975976e-05, 5.975994e-05, 
    5.975982e-05, 5.976002e-05, 5.975996e-05, 5.976039e-05, 5.976056e-05, 
    5.976063e-05, 5.976069e-05, 5.976084e-05, 5.976074e-05, 5.976078e-05, 
    5.976068e-05, 5.976062e-05, 5.976065e-05, 5.976046e-05, 5.976054e-05, 
    5.976015e-05, 5.976032e-05, 5.975989e-05, 5.975999e-05, 5.975986e-05, 
    5.975993e-05, 5.975982e-05, 5.975992e-05, 5.975974e-05, 5.975971e-05, 
    5.975973e-05, 5.975963e-05, 5.975992e-05, 5.975981e-05, 5.976065e-05, 
    5.976064e-05, 5.976062e-05, 5.976072e-05, 5.976073e-05, 5.976082e-05, 
    5.976074e-05, 5.97607e-05, 5.976062e-05, 5.976056e-05, 5.976051e-05, 
    5.97604e-05, 5.976028e-05, 5.976011e-05, 5.975998e-05, 5.97599e-05, 
    5.975995e-05, 5.975991e-05, 5.975996e-05, 5.975998e-05, 5.975972e-05, 
    5.975987e-05, 5.975965e-05, 5.975966e-05, 5.975976e-05, 5.975966e-05, 
    5.976064e-05, 5.976067e-05, 5.976077e-05, 5.976069e-05, 5.976083e-05, 
    5.976075e-05, 5.976071e-05, 5.976053e-05, 5.97605e-05, 5.976046e-05, 
    5.976039e-05, 5.97603e-05, 5.976014e-05, 5.976e-05, 5.975988e-05, 
    5.975989e-05, 5.975988e-05, 5.975986e-05, 5.975992e-05, 5.975984e-05, 
    5.975983e-05, 5.975987e-05, 5.975966e-05, 5.975972e-05, 5.975966e-05, 
    5.97597e-05, 5.976066e-05, 5.976061e-05, 5.976064e-05, 5.976059e-05, 
    5.976062e-05, 5.976047e-05, 5.976043e-05, 5.976021e-05, 5.97603e-05, 
    5.976016e-05, 5.976028e-05, 5.976026e-05, 5.976016e-05, 5.976028e-05, 
    5.976001e-05, 5.976019e-05, 5.975986e-05, 5.976004e-05, 5.975984e-05, 
    5.975988e-05, 5.975982e-05, 5.975977e-05, 5.97597e-05, 5.975958e-05, 
    5.975961e-05, 5.975951e-05, 5.976054e-05, 5.976048e-05, 5.976048e-05, 
    5.976042e-05, 5.976037e-05, 5.976027e-05, 5.97601e-05, 5.976016e-05, 
    5.976005e-05, 5.976003e-05, 5.97602e-05, 5.976009e-05, 5.976044e-05, 
    5.976038e-05, 5.976042e-05, 5.976054e-05, 5.976015e-05, 5.976035e-05, 
    5.975998e-05, 5.976009e-05, 5.975978e-05, 5.975993e-05, 5.975963e-05, 
    5.97595e-05, 5.975938e-05, 5.975923e-05, 5.976044e-05, 5.976049e-05, 
    5.976041e-05, 5.976031e-05, 5.976021e-05, 5.976008e-05, 5.976007e-05, 
    5.976004e-05, 5.975998e-05, 5.975993e-05, 5.976004e-05, 5.975992e-05, 
    5.976037e-05, 5.976013e-05, 5.97605e-05, 5.976039e-05, 5.976031e-05, 
    5.976035e-05, 5.976017e-05, 5.976013e-05, 5.975996e-05, 5.976005e-05, 
    5.975953e-05, 5.975976e-05, 5.975912e-05, 5.97593e-05, 5.97605e-05, 
    5.976044e-05, 5.976025e-05, 5.976034e-05, 5.976007e-05, 5.976001e-05, 
    5.975995e-05, 5.975988e-05, 5.975988e-05, 5.975984e-05, 5.975991e-05, 
    5.975984e-05, 5.976008e-05, 5.975998e-05, 5.976027e-05, 5.97602e-05, 
    5.976023e-05, 5.976027e-05, 5.976016e-05, 5.976004e-05, 5.976003e-05, 
    5.975999e-05, 5.975989e-05, 5.976007e-05, 5.97595e-05, 5.975985e-05, 
    5.976038e-05, 5.976027e-05, 5.976026e-05, 5.97603e-05, 5.976002e-05, 
    5.976012e-05, 5.975984e-05, 5.975991e-05, 5.975979e-05, 5.975985e-05, 
    5.975986e-05, 5.975994e-05, 5.975999e-05, 5.976011e-05, 5.976022e-05, 
    5.97603e-05, 5.976028e-05, 5.976019e-05, 5.976003e-05, 5.975988e-05, 
    5.975991e-05, 5.97598e-05, 5.976009e-05, 5.975997e-05, 5.976002e-05, 
    5.97599e-05, 5.976016e-05, 5.975994e-05, 5.976023e-05, 5.97602e-05, 
    5.976012e-05, 5.975996e-05, 5.975993e-05, 5.975989e-05, 5.975991e-05, 
    5.976003e-05, 5.976004e-05, 5.976012e-05, 5.976014e-05, 5.97602e-05, 
    5.976026e-05, 5.976021e-05, 5.976016e-05, 5.976003e-05, 5.97599e-05, 
    5.975977e-05, 5.975974e-05, 5.975958e-05, 5.975971e-05, 5.97595e-05, 
    5.975968e-05, 5.975937e-05, 5.975992e-05, 5.975968e-05, 5.976012e-05, 
    5.976007e-05, 5.975999e-05, 5.975979e-05, 5.97599e-05, 5.975977e-05, 
    5.976004e-05, 5.976019e-05, 5.976022e-05, 5.976029e-05, 5.976022e-05, 
    5.976023e-05, 5.976016e-05, 5.976018e-05, 5.976002e-05, 5.976011e-05, 
    5.975986e-05, 5.975977e-05, 5.975952e-05, 5.975937e-05, 5.975921e-05, 
    5.975914e-05, 5.975912e-05, 5.975911e-05 ;

 LITTERC_HR =
  9.949953e-13, 9.975261e-13, 9.970345e-13, 9.990735e-13, 9.97943e-13, 
    9.992776e-13, 9.95509e-13, 9.97626e-13, 9.96275e-13, 9.952239e-13, 
    1.003024e-12, 9.991646e-13, 1.00703e-12, 1.004573e-12, 1.01074e-12, 
    1.006647e-12, 1.011565e-12, 1.010623e-12, 1.013458e-12, 1.012646e-12, 
    1.016266e-12, 1.013833e-12, 1.018142e-12, 1.015686e-12, 1.01607e-12, 
    1.013752e-12, 9.999428e-13, 1.002544e-12, 9.997884e-13, 1.000159e-12, 
    9.999932e-13, 9.97966e-13, 9.969432e-13, 9.948024e-13, 9.951915e-13, 
    9.96764e-13, 1.000326e-12, 9.991183e-13, 1.002163e-12, 1.002095e-12, 
    1.005479e-12, 1.003954e-12, 1.009635e-12, 1.008022e-12, 1.01268e-12, 
    1.01151e-12, 1.012625e-12, 1.012287e-12, 1.01263e-12, 1.010912e-12, 
    1.011648e-12, 1.010137e-12, 1.004239e-12, 1.005974e-12, 1.000796e-12, 
    9.976748e-13, 9.956017e-13, 9.941288e-13, 9.943371e-13, 9.947339e-13, 
    9.967732e-13, 9.986896e-13, 1.000149e-12, 1.001124e-12, 1.002085e-12, 
    1.004988e-12, 1.006525e-12, 1.009961e-12, 1.009342e-12, 1.010391e-12, 
    1.011393e-12, 1.013074e-12, 1.012798e-12, 1.013538e-12, 1.010364e-12, 
    1.012474e-12, 1.008989e-12, 1.009943e-12, 1.002343e-12, 9.994445e-13, 
    9.982088e-13, 9.971288e-13, 9.944972e-13, 9.963147e-13, 9.955984e-13, 
    9.973029e-13, 9.98385e-13, 9.9785e-13, 1.001151e-12, 9.998679e-13, 
    1.006616e-12, 1.003712e-12, 1.011276e-12, 1.009469e-12, 1.011709e-12, 
    1.010567e-12, 1.012524e-12, 1.010762e-12, 1.013814e-12, 1.014477e-12, 
    1.014024e-12, 1.015766e-12, 1.010665e-12, 1.012625e-12, 9.978348e-13, 
    9.979221e-13, 9.983288e-13, 9.965403e-13, 9.96431e-13, 9.947916e-13, 
    9.962507e-13, 9.968715e-13, 9.98448e-13, 9.993793e-13, 1.000265e-12, 
    1.002209e-12, 1.004379e-12, 1.007411e-12, 1.009586e-12, 1.011043e-12, 
    1.01015e-12, 1.010938e-12, 1.010057e-12, 1.009644e-12, 1.014229e-12, 
    1.011655e-12, 1.015516e-12, 1.015302e-12, 1.013556e-12, 1.015326e-12, 
    9.979834e-13, 9.974813e-13, 9.957359e-13, 9.971019e-13, 9.94613e-13, 
    9.960061e-13, 9.968066e-13, 9.998941e-13, 1.000573e-12, 1.001201e-12, 
    1.002441e-12, 1.004032e-12, 1.006819e-12, 1.009242e-12, 1.011452e-12, 
    1.01129e-12, 1.011347e-12, 1.01184e-12, 1.010618e-12, 1.01204e-12, 
    1.012279e-12, 1.011655e-12, 1.015274e-12, 1.014241e-12, 1.015298e-12, 
    1.014625e-12, 9.976446e-13, 9.984896e-13, 9.980329e-13, 9.988913e-13, 
    9.982864e-13, 1.000974e-12, 1.001779e-12, 1.005544e-12, 1.004e-12, 
    1.006457e-12, 1.00425e-12, 1.004641e-12, 1.006536e-12, 1.00437e-12, 
    1.009108e-12, 1.005896e-12, 1.011859e-12, 1.008654e-12, 1.01206e-12, 
    1.011442e-12, 1.012465e-12, 1.01338e-12, 1.014531e-12, 1.016652e-12, 
    1.016162e-12, 1.017935e-12, 9.997489e-13, 1.000844e-12, 1.000748e-12, 
    1.001893e-12, 1.00274e-12, 1.004574e-12, 1.007512e-12, 1.006408e-12, 
    1.008435e-12, 1.008842e-12, 1.005762e-12, 1.007653e-12, 1.001576e-12, 
    1.002559e-12, 1.001974e-12, 9.99835e-13, 1.006662e-12, 1.003161e-12, 
    1.009622e-12, 1.007729e-12, 1.013249e-12, 1.010505e-12, 1.015891e-12, 
    1.018188e-12, 1.020349e-12, 1.02287e-12, 1.001441e-12, 1.000698e-12, 
    1.002029e-12, 1.003869e-12, 1.005577e-12, 1.007844e-12, 1.008076e-12, 
    1.0085e-12, 1.0096e-12, 1.010523e-12, 1.008634e-12, 1.010754e-12, 
    1.002785e-12, 1.006966e-12, 1.000416e-12, 1.00239e-12, 1.003761e-12, 
    1.00316e-12, 1.006282e-12, 1.007017e-12, 1.01e-12, 1.008459e-12, 
    1.017621e-12, 1.013572e-12, 1.024788e-12, 1.02166e-12, 1.000438e-12, 
    1.001439e-12, 1.004919e-12, 1.003264e-12, 1.007996e-12, 1.009158e-12, 
    1.010104e-12, 1.01131e-12, 1.011441e-12, 1.012156e-12, 1.010984e-12, 
    1.01211e-12, 1.007849e-12, 1.009754e-12, 1.004522e-12, 1.005797e-12, 
    1.005211e-12, 1.004568e-12, 1.006552e-12, 1.008664e-12, 1.00871e-12, 
    1.009386e-12, 1.011289e-12, 1.008015e-12, 1.018141e-12, 1.011892e-12, 
    1.00253e-12, 1.004455e-12, 1.004731e-12, 1.003986e-12, 1.009042e-12, 
    1.007211e-12, 1.012139e-12, 1.010808e-12, 1.012988e-12, 1.011905e-12, 
    1.011745e-12, 1.010354e-12, 1.009487e-12, 1.007295e-12, 1.00551e-12, 
    1.004094e-12, 1.004423e-12, 1.005979e-12, 1.008793e-12, 1.011452e-12, 
    1.01087e-12, 1.012822e-12, 1.007653e-12, 1.009821e-12, 1.008983e-12, 
    1.011168e-12, 1.006379e-12, 1.010455e-12, 1.005335e-12, 1.005785e-12, 
    1.007175e-12, 1.009968e-12, 1.010587e-12, 1.011246e-12, 1.010839e-12, 
    1.008864e-12, 1.008541e-12, 1.007141e-12, 1.006754e-12, 1.005687e-12, 
    1.004802e-12, 1.00561e-12, 1.006458e-12, 1.008866e-12, 1.011033e-12, 
    1.013393e-12, 1.01397e-12, 1.016721e-12, 1.014481e-12, 1.018175e-12, 
    1.015033e-12, 1.020471e-12, 1.010693e-12, 1.014942e-12, 1.007238e-12, 
    1.00807e-12, 1.009572e-12, 1.013015e-12, 1.011158e-12, 1.01333e-12, 
    1.008529e-12, 1.006032e-12, 1.005386e-12, 1.00418e-12, 1.005414e-12, 
    1.005314e-12, 1.006494e-12, 1.006115e-12, 1.008946e-12, 1.007425e-12, 
    1.011741e-12, 1.013314e-12, 1.017749e-12, 1.020462e-12, 1.023222e-12, 
    1.024439e-12, 1.024809e-12, 1.024964e-12 ;

 LITTERC_LOSS =
  1.842723e-12, 1.847409e-12, 1.846499e-12, 1.850275e-12, 1.848182e-12, 
    1.850653e-12, 1.843674e-12, 1.847595e-12, 1.845092e-12, 1.843146e-12, 
    1.857592e-12, 1.850444e-12, 1.865011e-12, 1.860461e-12, 1.871883e-12, 
    1.864302e-12, 1.87341e-12, 1.871666e-12, 1.876916e-12, 1.875413e-12, 
    1.882117e-12, 1.87761e-12, 1.88559e-12, 1.881042e-12, 1.881753e-12, 
    1.877461e-12, 1.851885e-12, 1.856702e-12, 1.851599e-12, 1.852287e-12, 
    1.851978e-12, 1.848224e-12, 1.84633e-12, 1.842365e-12, 1.843086e-12, 
    1.845998e-12, 1.852596e-12, 1.850358e-12, 1.855998e-12, 1.855871e-12, 
    1.862139e-12, 1.859314e-12, 1.869835e-12, 1.866848e-12, 1.875475e-12, 
    1.873307e-12, 1.875374e-12, 1.874747e-12, 1.875382e-12, 1.872201e-12, 
    1.873564e-12, 1.870765e-12, 1.859843e-12, 1.863055e-12, 1.853465e-12, 
    1.847685e-12, 1.843846e-12, 1.841118e-12, 1.841504e-12, 1.842238e-12, 
    1.846015e-12, 1.849564e-12, 1.852267e-12, 1.854073e-12, 1.855852e-12, 
    1.861229e-12, 1.864075e-12, 1.870438e-12, 1.869292e-12, 1.871235e-12, 
    1.873092e-12, 1.876205e-12, 1.875693e-12, 1.877064e-12, 1.871185e-12, 
    1.875093e-12, 1.868639e-12, 1.870405e-12, 1.85633e-12, 1.850962e-12, 
    1.848674e-12, 1.846674e-12, 1.8418e-12, 1.845166e-12, 1.843839e-12, 
    1.846996e-12, 1.849e-12, 1.848009e-12, 1.854122e-12, 1.851747e-12, 
    1.864244e-12, 1.858866e-12, 1.872875e-12, 1.869528e-12, 1.873677e-12, 
    1.871561e-12, 1.875186e-12, 1.871923e-12, 1.877575e-12, 1.878804e-12, 
    1.877964e-12, 1.881191e-12, 1.871742e-12, 1.875373e-12, 1.847981e-12, 
    1.848143e-12, 1.848896e-12, 1.845584e-12, 1.845381e-12, 1.842345e-12, 
    1.845047e-12, 1.846197e-12, 1.849117e-12, 1.850842e-12, 1.852481e-12, 
    1.856083e-12, 1.860102e-12, 1.865716e-12, 1.869745e-12, 1.872443e-12, 
    1.870789e-12, 1.872249e-12, 1.870617e-12, 1.869851e-12, 1.878343e-12, 
    1.873577e-12, 1.880726e-12, 1.880331e-12, 1.877097e-12, 1.880376e-12, 
    1.848257e-12, 1.847327e-12, 1.844094e-12, 1.846624e-12, 1.842014e-12, 
    1.844595e-12, 1.846077e-12, 1.851795e-12, 1.853052e-12, 1.854215e-12, 
    1.856512e-12, 1.859458e-12, 1.864621e-12, 1.869108e-12, 1.8732e-12, 
    1.8729e-12, 1.873006e-12, 1.873919e-12, 1.871656e-12, 1.87429e-12, 
    1.874732e-12, 1.873577e-12, 1.880278e-12, 1.878365e-12, 1.880323e-12, 
    1.879077e-12, 1.847629e-12, 1.849194e-12, 1.848348e-12, 1.849938e-12, 
    1.848818e-12, 1.853795e-12, 1.855287e-12, 1.862259e-12, 1.8594e-12, 
    1.86395e-12, 1.859863e-12, 1.860587e-12, 1.864096e-12, 1.860084e-12, 
    1.868859e-12, 1.86291e-12, 1.873954e-12, 1.868019e-12, 1.874326e-12, 
    1.873182e-12, 1.875076e-12, 1.876771e-12, 1.878903e-12, 1.882832e-12, 
    1.881923e-12, 1.885207e-12, 1.851526e-12, 1.853553e-12, 1.853376e-12, 
    1.855497e-12, 1.857065e-12, 1.860463e-12, 1.865904e-12, 1.863859e-12, 
    1.867614e-12, 1.868367e-12, 1.862663e-12, 1.866165e-12, 1.85491e-12, 
    1.85673e-12, 1.855647e-12, 1.851685e-12, 1.864329e-12, 1.857845e-12, 
    1.869811e-12, 1.866305e-12, 1.876529e-12, 1.871447e-12, 1.881422e-12, 
    1.885675e-12, 1.889679e-12, 1.894346e-12, 1.854661e-12, 1.853283e-12, 
    1.85575e-12, 1.859158e-12, 1.86232e-12, 1.866518e-12, 1.866948e-12, 
    1.867734e-12, 1.86977e-12, 1.87148e-12, 1.867981e-12, 1.871909e-12, 
    1.857149e-12, 1.864892e-12, 1.852762e-12, 1.856417e-12, 1.858957e-12, 
    1.857844e-12, 1.863626e-12, 1.864987e-12, 1.870512e-12, 1.867657e-12, 
    1.884625e-12, 1.877127e-12, 1.8979e-12, 1.892106e-12, 1.852802e-12, 
    1.854656e-12, 1.861102e-12, 1.858037e-12, 1.866799e-12, 1.868953e-12, 
    1.870703e-12, 1.872938e-12, 1.87318e-12, 1.874504e-12, 1.872335e-12, 
    1.874419e-12, 1.866528e-12, 1.870056e-12, 1.860367e-12, 1.862727e-12, 
    1.861642e-12, 1.86045e-12, 1.864126e-12, 1.868036e-12, 1.868122e-12, 
    1.869374e-12, 1.872899e-12, 1.866835e-12, 1.885588e-12, 1.874014e-12, 
    1.856677e-12, 1.860242e-12, 1.860754e-12, 1.859373e-12, 1.868737e-12, 
    1.865346e-12, 1.874472e-12, 1.872008e-12, 1.876045e-12, 1.874039e-12, 
    1.873744e-12, 1.871167e-12, 1.869561e-12, 1.865501e-12, 1.862196e-12, 
    1.859573e-12, 1.860183e-12, 1.863064e-12, 1.868276e-12, 1.873201e-12, 
    1.872123e-12, 1.875738e-12, 1.866165e-12, 1.870181e-12, 1.868629e-12, 
    1.872675e-12, 1.863804e-12, 1.871354e-12, 1.861872e-12, 1.862704e-12, 
    1.865279e-12, 1.870452e-12, 1.871598e-12, 1.872818e-12, 1.872066e-12, 
    1.868408e-12, 1.86781e-12, 1.865217e-12, 1.8645e-12, 1.862523e-12, 
    1.860885e-12, 1.862381e-12, 1.863951e-12, 1.868411e-12, 1.872424e-12, 
    1.876795e-12, 1.877864e-12, 1.882959e-12, 1.87881e-12, 1.885652e-12, 
    1.879832e-12, 1.889903e-12, 1.871794e-12, 1.879664e-12, 1.865397e-12, 
    1.866937e-12, 1.869719e-12, 1.876096e-12, 1.872656e-12, 1.87668e-12, 
    1.867786e-12, 1.863162e-12, 1.861967e-12, 1.859732e-12, 1.862018e-12, 
    1.861832e-12, 1.864018e-12, 1.863316e-12, 1.868558e-12, 1.865743e-12, 
    1.873736e-12, 1.876648e-12, 1.884862e-12, 1.889888e-12, 1.894999e-12, 
    1.897252e-12, 1.897938e-12, 1.898225e-12 ;

 LIVECROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVECROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 MEG_acetaldehyde =
  1.712902e-18, 1.713157e-18, 1.71311e-18, 1.713305e-18, 1.713199e-18, 
    1.713325e-18, 1.712964e-18, 1.713164e-18, 1.713037e-18, 1.712927e-18, 
    1.713678e-18, 1.713315e-18, 1.714078e-18, 1.713843e-18, 1.714442e-18, 
    1.714039e-18, 1.714525e-18, 1.714436e-18, 1.714717e-18, 1.714637e-18, 
    1.714985e-18, 1.714754e-18, 1.715174e-18, 1.714932e-18, 1.714968e-18, 
    1.714745e-18, 1.713393e-18, 1.713631e-18, 1.713378e-18, 1.713412e-18, 
    1.713398e-18, 1.7132e-18, 1.713096e-18, 1.712887e-18, 1.712924e-18, 
    1.713082e-18, 1.713427e-18, 1.713314e-18, 1.713611e-18, 1.713604e-18, 
    1.713932e-18, 1.713784e-18, 1.714339e-18, 1.714182e-18, 1.71464e-18, 
    1.714524e-18, 1.714634e-18, 1.714601e-18, 1.714634e-18, 1.714464e-18, 
    1.714537e-18, 1.714389e-18, 1.71381e-18, 1.713979e-18, 1.713474e-18, 
    1.713164e-18, 1.712971e-18, 1.712821e-18, 1.712841e-18, 1.712878e-18, 
    1.713083e-18, 1.713272e-18, 1.713414e-18, 1.713509e-18, 1.713603e-18, 
    1.713874e-18, 1.714029e-18, 1.714368e-18, 1.714311e-18, 1.714411e-18, 
    1.714513e-18, 1.714677e-18, 1.714651e-18, 1.714722e-18, 1.714412e-18, 
    1.714616e-18, 1.714278e-18, 1.71437e-18, 1.71361e-18, 1.713345e-18, 
    1.713217e-18, 1.713119e-18, 1.712856e-18, 1.713039e-18, 1.71297e-18, 
    1.713138e-18, 1.713242e-18, 1.713192e-18, 1.713512e-18, 1.713386e-18, 
    1.714038e-18, 1.713757e-18, 1.714501e-18, 1.714323e-18, 1.714544e-18, 
    1.714432e-18, 1.714622e-18, 1.714451e-18, 1.71475e-18, 1.714814e-18, 
    1.71477e-18, 1.714944e-18, 1.714441e-18, 1.714632e-18, 1.713189e-18, 
    1.713197e-18, 1.713238e-18, 1.713061e-18, 1.713051e-18, 1.712885e-18, 
    1.713035e-18, 1.713094e-18, 1.71325e-18, 1.713339e-18, 1.713424e-18, 
    1.713613e-18, 1.713821e-18, 1.714119e-18, 1.714335e-18, 1.714479e-18, 
    1.714392e-18, 1.714469e-18, 1.714382e-18, 1.714342e-18, 1.714789e-18, 
    1.714536e-18, 1.714919e-18, 1.714898e-18, 1.714723e-18, 1.7149e-18, 
    1.713203e-18, 1.713156e-18, 1.712985e-18, 1.713119e-18, 1.712868e-18, 
    1.71301e-18, 1.713085e-18, 1.713385e-18, 1.713455e-18, 1.713515e-18, 
    1.713637e-18, 1.713791e-18, 1.714061e-18, 1.714299e-18, 1.714519e-18, 
    1.714504e-18, 1.714509e-18, 1.714556e-18, 1.714437e-18, 1.714576e-18, 
    1.714598e-18, 1.714538e-18, 1.714895e-18, 1.714793e-18, 1.714898e-18, 
    1.714832e-18, 1.713172e-18, 1.713253e-18, 1.713209e-18, 1.713291e-18, 
    1.713231e-18, 1.713489e-18, 1.713566e-18, 1.713934e-18, 1.713787e-18, 
    1.714025e-18, 1.713813e-18, 1.71385e-18, 1.714025e-18, 1.713826e-18, 
    1.714283e-18, 1.713966e-18, 1.714558e-18, 1.714234e-18, 1.714578e-18, 
    1.714518e-18, 1.714619e-18, 1.714707e-18, 1.714822e-18, 1.715028e-18, 
    1.714981e-18, 1.715156e-18, 1.713375e-18, 1.713478e-18, 1.713473e-18, 
    1.713583e-18, 1.713664e-18, 1.713845e-18, 1.714131e-18, 1.714024e-18, 
    1.714223e-18, 1.714262e-18, 1.713962e-18, 1.714143e-18, 1.71355e-18, 
    1.713642e-18, 1.71359e-18, 1.713381e-18, 1.714044e-18, 1.713701e-18, 
    1.714338e-18, 1.714153e-18, 1.714694e-18, 1.714421e-18, 1.714954e-18, 
    1.715174e-18, 1.715397e-18, 1.715639e-18, 1.713539e-18, 1.713468e-18, 
    1.713598e-18, 1.713771e-18, 1.713942e-18, 1.714163e-18, 1.714188e-18, 
    1.714228e-18, 1.714338e-18, 1.714428e-18, 1.714238e-18, 1.714451e-18, 
    1.713657e-18, 1.714075e-18, 1.713438e-18, 1.713625e-18, 1.713762e-18, 
    1.713705e-18, 1.714013e-18, 1.714084e-18, 1.714373e-18, 1.714226e-18, 
    1.715116e-18, 1.714721e-18, 1.715835e-18, 1.71552e-18, 1.713442e-18, 
    1.71354e-18, 1.713875e-18, 1.713716e-18, 1.71418e-18, 1.714293e-18, 
    1.714387e-18, 1.714503e-18, 1.714518e-18, 1.714587e-18, 1.714473e-18, 
    1.714583e-18, 1.714164e-18, 1.714352e-18, 1.713841e-18, 1.713963e-18, 
    1.713908e-18, 1.713845e-18, 1.714039e-18, 1.71424e-18, 1.71425e-18, 
    1.714313e-18, 1.714483e-18, 1.714182e-18, 1.715157e-18, 1.714545e-18, 
    1.713646e-18, 1.713827e-18, 1.71386e-18, 1.713788e-18, 1.714281e-18, 
    1.714102e-18, 1.714586e-18, 1.714456e-18, 1.71467e-18, 1.714563e-18, 
    1.714547e-18, 1.714411e-18, 1.714325e-18, 1.714109e-18, 1.713935e-18, 
    1.713799e-18, 1.713831e-18, 1.71398e-18, 1.714254e-18, 1.714517e-18, 
    1.714458e-18, 1.714654e-18, 1.714146e-18, 1.714356e-18, 1.714273e-18, 
    1.71449e-18, 1.71402e-18, 1.714404e-18, 1.713921e-18, 1.713964e-18, 
    1.714098e-18, 1.714366e-18, 1.714434e-18, 1.714496e-18, 1.714459e-18, 
    1.714262e-18, 1.714232e-18, 1.714096e-18, 1.714056e-18, 1.713955e-18, 
    1.713868e-18, 1.713946e-18, 1.714026e-18, 1.714264e-18, 1.714475e-18, 
    1.714708e-18, 1.714767e-18, 1.715025e-18, 1.714807e-18, 1.71516e-18, 
    1.714849e-18, 1.715393e-18, 1.714434e-18, 1.714851e-18, 1.714106e-18, 
    1.714188e-18, 1.714329e-18, 1.714665e-18, 1.714489e-18, 1.714698e-18, 
    1.714231e-18, 1.713982e-18, 1.713925e-18, 1.713806e-18, 1.713928e-18, 
    1.713918e-18, 1.714034e-18, 1.713997e-18, 1.714272e-18, 1.714124e-18, 
    1.714545e-18, 1.714698e-18, 1.715136e-18, 1.715402e-18, 1.715681e-18, 
    1.715802e-18, 1.71584e-18, 1.715855e-18 ;

 MEG_acetic_acid =
  2.569353e-19, 2.569735e-19, 2.569666e-19, 2.569958e-19, 2.569799e-19, 
    2.569988e-19, 2.569445e-19, 2.569746e-19, 2.569556e-19, 2.569391e-19, 
    2.570517e-19, 2.569972e-19, 2.571118e-19, 2.570764e-19, 2.571663e-19, 
    2.571058e-19, 2.571787e-19, 2.571654e-19, 2.572075e-19, 2.571955e-19, 
    2.572477e-19, 2.572131e-19, 2.572761e-19, 2.572398e-19, 2.572452e-19, 
    2.572118e-19, 2.570089e-19, 2.570446e-19, 2.570066e-19, 2.570118e-19, 
    2.570096e-19, 2.569799e-19, 2.569644e-19, 2.569331e-19, 2.569386e-19, 
    2.569624e-19, 2.570141e-19, 2.569971e-19, 2.570416e-19, 2.570406e-19, 
    2.570898e-19, 2.570675e-19, 2.571509e-19, 2.571274e-19, 2.57196e-19, 
    2.571786e-19, 2.57195e-19, 2.571901e-19, 2.571951e-19, 2.571696e-19, 
    2.571805e-19, 2.571584e-19, 2.570715e-19, 2.570968e-19, 2.570212e-19, 
    2.569746e-19, 2.569457e-19, 2.569232e-19, 2.569262e-19, 2.569317e-19, 
    2.569625e-19, 2.569908e-19, 2.570122e-19, 2.570263e-19, 2.570404e-19, 
    2.570811e-19, 2.571044e-19, 2.571552e-19, 2.571467e-19, 2.571616e-19, 
    2.571769e-19, 2.572016e-19, 2.571976e-19, 2.572083e-19, 2.571617e-19, 
    2.571925e-19, 2.571417e-19, 2.571555e-19, 2.570415e-19, 2.570018e-19, 
    2.569826e-19, 2.569678e-19, 2.569284e-19, 2.569559e-19, 2.569455e-19, 
    2.569707e-19, 2.569863e-19, 2.569787e-19, 2.570267e-19, 2.57008e-19, 
    2.571058e-19, 2.570636e-19, 2.571751e-19, 2.571485e-19, 2.571816e-19, 
    2.571648e-19, 2.571933e-19, 2.571677e-19, 2.572126e-19, 2.57222e-19, 
    2.572155e-19, 2.572415e-19, 2.571662e-19, 2.571948e-19, 2.569784e-19, 
    2.569796e-19, 2.569856e-19, 2.569591e-19, 2.569576e-19, 2.569328e-19, 
    2.569553e-19, 2.569641e-19, 2.569875e-19, 2.570008e-19, 2.570137e-19, 
    2.57042e-19, 2.570732e-19, 2.571178e-19, 2.571502e-19, 2.571718e-19, 
    2.571587e-19, 2.571703e-19, 2.571573e-19, 2.571513e-19, 2.572183e-19, 
    2.571804e-19, 2.572378e-19, 2.572347e-19, 2.572085e-19, 2.572351e-19, 
    2.569805e-19, 2.569734e-19, 2.569477e-19, 2.569678e-19, 2.569303e-19, 
    2.569515e-19, 2.569628e-19, 2.570078e-19, 2.570183e-19, 2.570272e-19, 
    2.570455e-19, 2.570686e-19, 2.571092e-19, 2.571449e-19, 2.571779e-19, 
    2.571755e-19, 2.571763e-19, 2.571834e-19, 2.571655e-19, 2.571864e-19, 
    2.571897e-19, 2.571807e-19, 2.572343e-19, 2.57219e-19, 2.572346e-19, 
    2.572248e-19, 2.569758e-19, 2.569879e-19, 2.569813e-19, 2.569936e-19, 
    2.569847e-19, 2.570233e-19, 2.570349e-19, 2.5709e-19, 2.57068e-19, 
    2.571038e-19, 2.570719e-19, 2.570774e-19, 2.571038e-19, 2.570739e-19, 
    2.571424e-19, 2.570949e-19, 2.571837e-19, 2.571351e-19, 2.571867e-19, 
    2.571777e-19, 2.571928e-19, 2.572061e-19, 2.572232e-19, 2.572542e-19, 
    2.572471e-19, 2.572734e-19, 2.570063e-19, 2.570218e-19, 2.570209e-19, 
    2.570375e-19, 2.570497e-19, 2.570768e-19, 2.571196e-19, 2.571036e-19, 
    2.571335e-19, 2.571393e-19, 2.570943e-19, 2.571214e-19, 2.570325e-19, 
    2.570463e-19, 2.570385e-19, 2.570072e-19, 2.571066e-19, 2.570552e-19, 
    2.571507e-19, 2.571229e-19, 2.572041e-19, 2.571632e-19, 2.572431e-19, 
    2.57276e-19, 2.573095e-19, 2.573458e-19, 2.570308e-19, 2.570202e-19, 
    2.570396e-19, 2.570656e-19, 2.570912e-19, 2.571245e-19, 2.571282e-19, 
    2.571342e-19, 2.571506e-19, 2.571642e-19, 2.571357e-19, 2.571676e-19, 
    2.570485e-19, 2.571113e-19, 2.570157e-19, 2.570437e-19, 2.570643e-19, 
    2.570558e-19, 2.57102e-19, 2.571126e-19, 2.571559e-19, 2.571338e-19, 
    2.572674e-19, 2.572082e-19, 2.573752e-19, 2.573281e-19, 2.570164e-19, 
    2.57031e-19, 2.570813e-19, 2.570574e-19, 2.57127e-19, 2.571439e-19, 
    2.571581e-19, 2.571754e-19, 2.571776e-19, 2.57188e-19, 2.57171e-19, 
    2.571875e-19, 2.571245e-19, 2.571527e-19, 2.570762e-19, 2.570945e-19, 
    2.570862e-19, 2.570768e-19, 2.571059e-19, 2.57136e-19, 2.571375e-19, 
    2.57147e-19, 2.571724e-19, 2.571273e-19, 2.572736e-19, 2.571817e-19, 
    2.570469e-19, 2.570741e-19, 2.570789e-19, 2.570682e-19, 2.571421e-19, 
    2.571153e-19, 2.571878e-19, 2.571684e-19, 2.572005e-19, 2.571845e-19, 
    2.571821e-19, 2.571617e-19, 2.571488e-19, 2.571163e-19, 2.570902e-19, 
    2.570698e-19, 2.570747e-19, 2.57097e-19, 2.57138e-19, 2.571775e-19, 
    2.571687e-19, 2.571981e-19, 2.571219e-19, 2.571534e-19, 2.571409e-19, 
    2.571736e-19, 2.57103e-19, 2.571606e-19, 2.570881e-19, 2.570946e-19, 
    2.571147e-19, 2.57155e-19, 2.571651e-19, 2.571744e-19, 2.571688e-19, 
    2.571392e-19, 2.571347e-19, 2.571144e-19, 2.571084e-19, 2.570932e-19, 
    2.570803e-19, 2.570919e-19, 2.57104e-19, 2.571396e-19, 2.571713e-19, 
    2.572062e-19, 2.57215e-19, 2.572538e-19, 2.572211e-19, 2.572739e-19, 
    2.572273e-19, 2.57309e-19, 2.571651e-19, 2.572276e-19, 2.571159e-19, 
    2.571281e-19, 2.571493e-19, 2.571998e-19, 2.571734e-19, 2.572047e-19, 
    2.571346e-19, 2.570974e-19, 2.570887e-19, 2.570709e-19, 2.570892e-19, 
    2.570877e-19, 2.571051e-19, 2.570995e-19, 2.571408e-19, 2.571186e-19, 
    2.571818e-19, 2.572047e-19, 2.572704e-19, 2.573102e-19, 2.573522e-19, 
    2.573703e-19, 2.573759e-19, 2.573782e-19 ;

 MEG_acetone =
  8.551299e-17, 8.552143e-17, 8.551989e-17, 8.552635e-17, 8.552284e-17, 
    8.552701e-17, 8.551504e-17, 8.552169e-17, 8.551749e-17, 8.551383e-17, 
    8.553867e-17, 8.552666e-17, 8.555192e-17, 8.554413e-17, 8.556397e-17, 
    8.555061e-17, 8.556669e-17, 8.556376e-17, 8.557304e-17, 8.557039e-17, 
    8.55819e-17, 8.557426e-17, 8.558817e-17, 8.558017e-17, 8.558136e-17, 
    8.557399e-17, 8.552924e-17, 8.553712e-17, 8.552873e-17, 8.552987e-17, 
    8.55294e-17, 8.552285e-17, 8.551943e-17, 8.55125e-17, 8.551373e-17, 
    8.551897e-17, 8.553038e-17, 8.552662e-17, 8.553644e-17, 8.553623e-17, 
    8.554707e-17, 8.554217e-17, 8.556055e-17, 8.555536e-17, 8.55705e-17, 
    8.556667e-17, 8.557029e-17, 8.556921e-17, 8.557031e-17, 8.556469e-17, 
    8.556708e-17, 8.55622e-17, 8.554305e-17, 8.554863e-17, 8.553194e-17, 
    8.552167e-17, 8.55153e-17, 8.551033e-17, 8.551098e-17, 8.55122e-17, 
    8.5519e-17, 8.552525e-17, 8.552996e-17, 8.553308e-17, 8.553619e-17, 
    8.554516e-17, 8.555029e-17, 8.55615e-17, 8.555963e-17, 8.556293e-17, 
    8.556629e-17, 8.557174e-17, 8.557086e-17, 8.557323e-17, 8.556295e-17, 
    8.556972e-17, 8.555853e-17, 8.556157e-17, 8.553644e-17, 8.552766e-17, 
    8.552343e-17, 8.552017e-17, 8.551148e-17, 8.551754e-17, 8.551527e-17, 
    8.552081e-17, 8.552426e-17, 8.552258e-17, 8.553317e-17, 8.552903e-17, 
    8.555059e-17, 8.554129e-17, 8.55659e-17, 8.556003e-17, 8.556733e-17, 
    8.556363e-17, 8.556992e-17, 8.556426e-17, 8.557416e-17, 8.557625e-17, 
    8.557481e-17, 8.558054e-17, 8.556393e-17, 8.557023e-17, 8.552251e-17, 
    8.552278e-17, 8.55241e-17, 8.551825e-17, 8.551793e-17, 8.551243e-17, 
    8.551742e-17, 8.551935e-17, 8.552451e-17, 8.552745e-17, 8.553028e-17, 
    8.553653e-17, 8.554342e-17, 8.555325e-17, 8.55604e-17, 8.556518e-17, 
    8.556229e-17, 8.556483e-17, 8.556197e-17, 8.556064e-17, 8.557543e-17, 
    8.556707e-17, 8.557972e-17, 8.557904e-17, 8.557326e-17, 8.557912e-17, 
    8.552298e-17, 8.55214e-17, 8.551575e-17, 8.552018e-17, 8.551187e-17, 
    8.551659e-17, 8.551907e-17, 8.552899e-17, 8.553131e-17, 8.553328e-17, 
    8.553731e-17, 8.554241e-17, 8.555135e-17, 8.555923e-17, 8.556651e-17, 
    8.556598e-17, 8.556617e-17, 8.556773e-17, 8.556377e-17, 8.556839e-17, 
    8.556911e-17, 8.556714e-17, 8.557894e-17, 8.557558e-17, 8.557902e-17, 
    8.557684e-17, 8.552193e-17, 8.552461e-17, 8.552315e-17, 8.552586e-17, 
    8.55239e-17, 8.553242e-17, 8.553498e-17, 8.554713e-17, 8.554228e-17, 
    8.555016e-17, 8.554313e-17, 8.554435e-17, 8.555016e-17, 8.554356e-17, 
    8.555868e-17, 8.55482e-17, 8.556779e-17, 8.555707e-17, 8.556845e-17, 
    8.556648e-17, 8.556981e-17, 8.557273e-17, 8.557651e-17, 8.558334e-17, 
    8.558178e-17, 8.558758e-17, 8.552866e-17, 8.553208e-17, 8.553188e-17, 
    8.553554e-17, 8.553823e-17, 8.554421e-17, 8.555365e-17, 8.555013e-17, 
    8.555671e-17, 8.555799e-17, 8.554806e-17, 8.555405e-17, 8.553445e-17, 
    8.55375e-17, 8.553576e-17, 8.552886e-17, 8.555078e-17, 8.553945e-17, 
    8.55605e-17, 8.555438e-17, 8.55723e-17, 8.556326e-17, 8.558089e-17, 
    8.558816e-17, 8.559553e-17, 8.560355e-17, 8.553406e-17, 8.553173e-17, 
    8.553601e-17, 8.554174e-17, 8.55474e-17, 8.555473e-17, 8.555554e-17, 
    8.555688e-17, 8.556049e-17, 8.556348e-17, 8.55572e-17, 8.556424e-17, 
    8.553797e-17, 8.555182e-17, 8.553074e-17, 8.553692e-17, 8.554145e-17, 
    8.553958e-17, 8.554976e-17, 8.555211e-17, 8.556166e-17, 8.555679e-17, 
    8.558627e-17, 8.557318e-17, 8.561004e-17, 8.559964e-17, 8.553089e-17, 
    8.553411e-17, 8.554521e-17, 8.553993e-17, 8.555528e-17, 8.5559e-17, 
    8.556214e-17, 8.556596e-17, 8.556645e-17, 8.556874e-17, 8.556499e-17, 
    8.556863e-17, 8.555474e-17, 8.556096e-17, 8.554407e-17, 8.554811e-17, 
    8.554629e-17, 8.554421e-17, 8.555062e-17, 8.555726e-17, 8.555759e-17, 
    8.555969e-17, 8.55653e-17, 8.555534e-17, 8.558762e-17, 8.556734e-17, 
    8.553762e-17, 8.55436e-17, 8.554468e-17, 8.554231e-17, 8.555863e-17, 
    8.555269e-17, 8.55687e-17, 8.556441e-17, 8.55715e-17, 8.556796e-17, 
    8.556743e-17, 8.556293e-17, 8.556008e-17, 8.555293e-17, 8.554716e-17, 
    8.554268e-17, 8.554375e-17, 8.554867e-17, 8.555771e-17, 8.556642e-17, 
    8.556449e-17, 8.557096e-17, 8.555416e-17, 8.55611e-17, 8.555835e-17, 
    8.556555e-17, 8.555e-17, 8.556269e-17, 8.554669e-17, 8.554813e-17, 
    8.555258e-17, 8.556145e-17, 8.556369e-17, 8.556575e-17, 8.556452e-17, 
    8.555798e-17, 8.555699e-17, 8.555251e-17, 8.555119e-17, 8.554783e-17, 
    8.554497e-17, 8.554754e-17, 8.55502e-17, 8.555806e-17, 8.556504e-17, 
    8.557274e-17, 8.55747e-17, 8.558325e-17, 8.557604e-17, 8.55877e-17, 
    8.55774e-17, 8.559543e-17, 8.556369e-17, 8.557747e-17, 8.555284e-17, 
    8.555553e-17, 8.556021e-17, 8.557134e-17, 8.556552e-17, 8.557242e-17, 
    8.555696e-17, 8.554875e-17, 8.554685e-17, 8.554292e-17, 8.554693e-17, 
    8.554662e-17, 8.555044e-17, 8.554922e-17, 8.555832e-17, 8.555344e-17, 
    8.556737e-17, 8.557241e-17, 8.558691e-17, 8.55957e-17, 8.560497e-17, 
    8.560896e-17, 8.56102e-17, 8.561071e-17 ;

 MEG_carene_3 =
  3.305598e-17, 3.305931e-17, 3.305871e-17, 3.306125e-17, 3.305987e-17, 
    3.306152e-17, 3.305679e-17, 3.305941e-17, 3.305776e-17, 3.305631e-17, 
    3.306611e-17, 3.306138e-17, 3.307135e-17, 3.306827e-17, 3.30761e-17, 
    3.307083e-17, 3.307718e-17, 3.307602e-17, 3.307968e-17, 3.307864e-17, 
    3.308318e-17, 3.308016e-17, 3.308565e-17, 3.308249e-17, 3.308296e-17, 
    3.308005e-17, 3.30624e-17, 3.30655e-17, 3.30622e-17, 3.306264e-17, 
    3.306246e-17, 3.305987e-17, 3.305852e-17, 3.305579e-17, 3.305627e-17, 
    3.305834e-17, 3.306285e-17, 3.306136e-17, 3.306524e-17, 3.306515e-17, 
    3.306943e-17, 3.30675e-17, 3.307475e-17, 3.30727e-17, 3.307868e-17, 
    3.307716e-17, 3.30786e-17, 3.307817e-17, 3.30786e-17, 3.307638e-17, 
    3.307733e-17, 3.30754e-17, 3.306785e-17, 3.307005e-17, 3.306346e-17, 
    3.305941e-17, 3.305689e-17, 3.305493e-17, 3.305519e-17, 3.305567e-17, 
    3.305835e-17, 3.306082e-17, 3.306268e-17, 3.306391e-17, 3.306514e-17, 
    3.306868e-17, 3.30707e-17, 3.307513e-17, 3.307439e-17, 3.307569e-17, 
    3.307702e-17, 3.307916e-17, 3.307882e-17, 3.307975e-17, 3.30757e-17, 
    3.307837e-17, 3.307395e-17, 3.307515e-17, 3.306523e-17, 3.306177e-17, 
    3.30601e-17, 3.305882e-17, 3.305538e-17, 3.305778e-17, 3.305688e-17, 
    3.305907e-17, 3.306043e-17, 3.305977e-17, 3.306394e-17, 3.306231e-17, 
    3.307082e-17, 3.306715e-17, 3.307686e-17, 3.307455e-17, 3.307742e-17, 
    3.307597e-17, 3.307845e-17, 3.307622e-17, 3.308012e-17, 3.308094e-17, 
    3.308038e-17, 3.308264e-17, 3.307608e-17, 3.307857e-17, 3.305974e-17, 
    3.305984e-17, 3.306037e-17, 3.305806e-17, 3.305793e-17, 3.305576e-17, 
    3.305773e-17, 3.305849e-17, 3.306053e-17, 3.306169e-17, 3.306281e-17, 
    3.306527e-17, 3.306799e-17, 3.307187e-17, 3.307469e-17, 3.307658e-17, 
    3.307544e-17, 3.307644e-17, 3.307531e-17, 3.307479e-17, 3.308062e-17, 
    3.307732e-17, 3.308231e-17, 3.308205e-17, 3.307977e-17, 3.308208e-17, 
    3.305992e-17, 3.30593e-17, 3.305707e-17, 3.305882e-17, 3.305554e-17, 
    3.30574e-17, 3.305838e-17, 3.306229e-17, 3.306321e-17, 3.306399e-17, 
    3.306558e-17, 3.306759e-17, 3.307112e-17, 3.307423e-17, 3.30771e-17, 
    3.30769e-17, 3.307697e-17, 3.307759e-17, 3.307602e-17, 3.307784e-17, 
    3.307813e-17, 3.307735e-17, 3.308201e-17, 3.308068e-17, 3.308204e-17, 
    3.308118e-17, 3.305951e-17, 3.306057e-17, 3.305999e-17, 3.306106e-17, 
    3.306029e-17, 3.306365e-17, 3.306466e-17, 3.306945e-17, 3.306754e-17, 
    3.307065e-17, 3.306788e-17, 3.306836e-17, 3.307065e-17, 3.306804e-17, 
    3.307401e-17, 3.306988e-17, 3.307761e-17, 3.307338e-17, 3.307787e-17, 
    3.307709e-17, 3.30784e-17, 3.307955e-17, 3.308105e-17, 3.308374e-17, 
    3.308313e-17, 3.308542e-17, 3.306216e-17, 3.306351e-17, 3.306344e-17, 
    3.306488e-17, 3.306594e-17, 3.30683e-17, 3.307203e-17, 3.307064e-17, 
    3.307324e-17, 3.307374e-17, 3.306982e-17, 3.307219e-17, 3.306445e-17, 
    3.306565e-17, 3.306497e-17, 3.306224e-17, 3.30709e-17, 3.306642e-17, 
    3.307473e-17, 3.307232e-17, 3.307939e-17, 3.307582e-17, 3.308278e-17, 
    3.308565e-17, 3.308856e-17, 3.309172e-17, 3.30643e-17, 3.306338e-17, 
    3.306507e-17, 3.306733e-17, 3.306956e-17, 3.307245e-17, 3.307277e-17, 
    3.30733e-17, 3.307473e-17, 3.307591e-17, 3.307343e-17, 3.307621e-17, 
    3.306584e-17, 3.307131e-17, 3.306298e-17, 3.306543e-17, 3.306722e-17, 
    3.306648e-17, 3.307049e-17, 3.307142e-17, 3.307519e-17, 3.307327e-17, 
    3.30849e-17, 3.307974e-17, 3.309428e-17, 3.309018e-17, 3.306304e-17, 
    3.306431e-17, 3.30687e-17, 3.306661e-17, 3.307267e-17, 3.307414e-17, 
    3.307538e-17, 3.307688e-17, 3.307708e-17, 3.307798e-17, 3.30765e-17, 
    3.307794e-17, 3.307246e-17, 3.307491e-17, 3.306825e-17, 3.306984e-17, 
    3.306912e-17, 3.30683e-17, 3.307083e-17, 3.307345e-17, 3.307358e-17, 
    3.307441e-17, 3.307662e-17, 3.30727e-17, 3.308543e-17, 3.307743e-17, 
    3.30657e-17, 3.306806e-17, 3.306849e-17, 3.306755e-17, 3.307399e-17, 
    3.307165e-17, 3.307797e-17, 3.307628e-17, 3.307907e-17, 3.307768e-17, 
    3.307747e-17, 3.307569e-17, 3.307457e-17, 3.307174e-17, 3.306947e-17, 
    3.30677e-17, 3.306812e-17, 3.307006e-17, 3.307363e-17, 3.307707e-17, 
    3.30763e-17, 3.307886e-17, 3.307223e-17, 3.307497e-17, 3.307388e-17, 
    3.307673e-17, 3.307058e-17, 3.307559e-17, 3.306928e-17, 3.306985e-17, 
    3.30716e-17, 3.30751e-17, 3.307599e-17, 3.30768e-17, 3.307632e-17, 
    3.307373e-17, 3.307334e-17, 3.307158e-17, 3.307105e-17, 3.306973e-17, 
    3.30686e-17, 3.306962e-17, 3.307067e-17, 3.307377e-17, 3.307652e-17, 
    3.307956e-17, 3.308033e-17, 3.308371e-17, 3.308086e-17, 3.308546e-17, 
    3.30814e-17, 3.308851e-17, 3.307599e-17, 3.308143e-17, 3.307171e-17, 
    3.307277e-17, 3.307461e-17, 3.307901e-17, 3.307671e-17, 3.307944e-17, 
    3.307333e-17, 3.307009e-17, 3.306934e-17, 3.306779e-17, 3.306938e-17, 
    3.306925e-17, 3.307076e-17, 3.307028e-17, 3.307387e-17, 3.307194e-17, 
    3.307744e-17, 3.307943e-17, 3.308515e-17, 3.308862e-17, 3.309228e-17, 
    3.309386e-17, 3.309434e-17, 3.309454e-17 ;

 MEG_ethanol =
  1.712902e-18, 1.713157e-18, 1.71311e-18, 1.713305e-18, 1.713199e-18, 
    1.713325e-18, 1.712964e-18, 1.713164e-18, 1.713037e-18, 1.712927e-18, 
    1.713678e-18, 1.713315e-18, 1.714078e-18, 1.713843e-18, 1.714442e-18, 
    1.714039e-18, 1.714525e-18, 1.714436e-18, 1.714717e-18, 1.714637e-18, 
    1.714985e-18, 1.714754e-18, 1.715174e-18, 1.714932e-18, 1.714968e-18, 
    1.714745e-18, 1.713393e-18, 1.713631e-18, 1.713378e-18, 1.713412e-18, 
    1.713398e-18, 1.7132e-18, 1.713096e-18, 1.712887e-18, 1.712924e-18, 
    1.713082e-18, 1.713427e-18, 1.713314e-18, 1.713611e-18, 1.713604e-18, 
    1.713932e-18, 1.713784e-18, 1.714339e-18, 1.714182e-18, 1.71464e-18, 
    1.714524e-18, 1.714634e-18, 1.714601e-18, 1.714634e-18, 1.714464e-18, 
    1.714537e-18, 1.714389e-18, 1.71381e-18, 1.713979e-18, 1.713474e-18, 
    1.713164e-18, 1.712971e-18, 1.712821e-18, 1.712841e-18, 1.712878e-18, 
    1.713083e-18, 1.713272e-18, 1.713414e-18, 1.713509e-18, 1.713603e-18, 
    1.713874e-18, 1.714029e-18, 1.714368e-18, 1.714311e-18, 1.714411e-18, 
    1.714513e-18, 1.714677e-18, 1.714651e-18, 1.714722e-18, 1.714412e-18, 
    1.714616e-18, 1.714278e-18, 1.71437e-18, 1.71361e-18, 1.713345e-18, 
    1.713217e-18, 1.713119e-18, 1.712856e-18, 1.713039e-18, 1.71297e-18, 
    1.713138e-18, 1.713242e-18, 1.713192e-18, 1.713512e-18, 1.713386e-18, 
    1.714038e-18, 1.713757e-18, 1.714501e-18, 1.714323e-18, 1.714544e-18, 
    1.714432e-18, 1.714622e-18, 1.714451e-18, 1.71475e-18, 1.714814e-18, 
    1.71477e-18, 1.714944e-18, 1.714441e-18, 1.714632e-18, 1.713189e-18, 
    1.713197e-18, 1.713238e-18, 1.713061e-18, 1.713051e-18, 1.712885e-18, 
    1.713035e-18, 1.713094e-18, 1.71325e-18, 1.713339e-18, 1.713424e-18, 
    1.713613e-18, 1.713821e-18, 1.714119e-18, 1.714335e-18, 1.714479e-18, 
    1.714392e-18, 1.714469e-18, 1.714382e-18, 1.714342e-18, 1.714789e-18, 
    1.714536e-18, 1.714919e-18, 1.714898e-18, 1.714723e-18, 1.7149e-18, 
    1.713203e-18, 1.713156e-18, 1.712985e-18, 1.713119e-18, 1.712868e-18, 
    1.71301e-18, 1.713085e-18, 1.713385e-18, 1.713455e-18, 1.713515e-18, 
    1.713637e-18, 1.713791e-18, 1.714061e-18, 1.714299e-18, 1.714519e-18, 
    1.714504e-18, 1.714509e-18, 1.714556e-18, 1.714437e-18, 1.714576e-18, 
    1.714598e-18, 1.714538e-18, 1.714895e-18, 1.714793e-18, 1.714898e-18, 
    1.714832e-18, 1.713172e-18, 1.713253e-18, 1.713209e-18, 1.713291e-18, 
    1.713231e-18, 1.713489e-18, 1.713566e-18, 1.713934e-18, 1.713787e-18, 
    1.714025e-18, 1.713813e-18, 1.71385e-18, 1.714025e-18, 1.713826e-18, 
    1.714283e-18, 1.713966e-18, 1.714558e-18, 1.714234e-18, 1.714578e-18, 
    1.714518e-18, 1.714619e-18, 1.714707e-18, 1.714822e-18, 1.715028e-18, 
    1.714981e-18, 1.715156e-18, 1.713375e-18, 1.713478e-18, 1.713473e-18, 
    1.713583e-18, 1.713664e-18, 1.713845e-18, 1.714131e-18, 1.714024e-18, 
    1.714223e-18, 1.714262e-18, 1.713962e-18, 1.714143e-18, 1.71355e-18, 
    1.713642e-18, 1.71359e-18, 1.713381e-18, 1.714044e-18, 1.713701e-18, 
    1.714338e-18, 1.714153e-18, 1.714694e-18, 1.714421e-18, 1.714954e-18, 
    1.715174e-18, 1.715397e-18, 1.715639e-18, 1.713539e-18, 1.713468e-18, 
    1.713598e-18, 1.713771e-18, 1.713942e-18, 1.714163e-18, 1.714188e-18, 
    1.714228e-18, 1.714338e-18, 1.714428e-18, 1.714238e-18, 1.714451e-18, 
    1.713657e-18, 1.714075e-18, 1.713438e-18, 1.713625e-18, 1.713762e-18, 
    1.713705e-18, 1.714013e-18, 1.714084e-18, 1.714373e-18, 1.714226e-18, 
    1.715116e-18, 1.714721e-18, 1.715835e-18, 1.71552e-18, 1.713442e-18, 
    1.71354e-18, 1.713875e-18, 1.713716e-18, 1.71418e-18, 1.714293e-18, 
    1.714387e-18, 1.714503e-18, 1.714518e-18, 1.714587e-18, 1.714473e-18, 
    1.714583e-18, 1.714164e-18, 1.714352e-18, 1.713841e-18, 1.713963e-18, 
    1.713908e-18, 1.713845e-18, 1.714039e-18, 1.71424e-18, 1.71425e-18, 
    1.714313e-18, 1.714483e-18, 1.714182e-18, 1.715157e-18, 1.714545e-18, 
    1.713646e-18, 1.713827e-18, 1.71386e-18, 1.713788e-18, 1.714281e-18, 
    1.714102e-18, 1.714586e-18, 1.714456e-18, 1.71467e-18, 1.714563e-18, 
    1.714547e-18, 1.714411e-18, 1.714325e-18, 1.714109e-18, 1.713935e-18, 
    1.713799e-18, 1.713831e-18, 1.71398e-18, 1.714254e-18, 1.714517e-18, 
    1.714458e-18, 1.714654e-18, 1.714146e-18, 1.714356e-18, 1.714273e-18, 
    1.71449e-18, 1.71402e-18, 1.714404e-18, 1.713921e-18, 1.713964e-18, 
    1.714098e-18, 1.714366e-18, 1.714434e-18, 1.714496e-18, 1.714459e-18, 
    1.714262e-18, 1.714232e-18, 1.714096e-18, 1.714056e-18, 1.713955e-18, 
    1.713868e-18, 1.713946e-18, 1.714026e-18, 1.714264e-18, 1.714475e-18, 
    1.714708e-18, 1.714767e-18, 1.715025e-18, 1.714807e-18, 1.71516e-18, 
    1.714849e-18, 1.715393e-18, 1.714434e-18, 1.714851e-18, 1.714106e-18, 
    1.714188e-18, 1.714329e-18, 1.714665e-18, 1.714489e-18, 1.714698e-18, 
    1.714231e-18, 1.713982e-18, 1.713925e-18, 1.713806e-18, 1.713928e-18, 
    1.713918e-18, 1.714034e-18, 1.713997e-18, 1.714272e-18, 1.714124e-18, 
    1.714545e-18, 1.714698e-18, 1.715136e-18, 1.715402e-18, 1.715681e-18, 
    1.715802e-18, 1.71584e-18, 1.715855e-18 ;

 MEG_formaldehyde =
  3.425804e-19, 3.426313e-19, 3.426221e-19, 3.426611e-19, 3.426398e-19, 
    3.426651e-19, 3.425927e-19, 3.426329e-19, 3.426075e-19, 3.425855e-19, 
    3.427355e-19, 3.42663e-19, 3.428157e-19, 3.427685e-19, 3.428885e-19, 
    3.428077e-19, 3.42905e-19, 3.428872e-19, 3.429433e-19, 3.429273e-19, 
    3.429969e-19, 3.429507e-19, 3.430348e-19, 3.429864e-19, 3.429936e-19, 
    3.42949e-19, 3.426786e-19, 3.427262e-19, 3.426755e-19, 3.426823e-19, 
    3.426795e-19, 3.426399e-19, 3.426192e-19, 3.425774e-19, 3.425849e-19, 
    3.426165e-19, 3.426854e-19, 3.426627e-19, 3.427221e-19, 3.427208e-19, 
    3.427864e-19, 3.427567e-19, 3.428678e-19, 3.428365e-19, 3.42928e-19, 
    3.429048e-19, 3.429267e-19, 3.429202e-19, 3.429268e-19, 3.428928e-19, 
    3.429073e-19, 3.428778e-19, 3.42762e-19, 3.427957e-19, 3.426949e-19, 
    3.426328e-19, 3.425943e-19, 3.425643e-19, 3.425682e-19, 3.425756e-19, 
    3.426166e-19, 3.426544e-19, 3.426829e-19, 3.427018e-19, 3.427206e-19, 
    3.427748e-19, 3.428058e-19, 3.428736e-19, 3.428623e-19, 3.428822e-19, 
    3.429025e-19, 3.429355e-19, 3.429302e-19, 3.429445e-19, 3.428823e-19, 
    3.429233e-19, 3.428556e-19, 3.42874e-19, 3.42722e-19, 3.42669e-19, 
    3.426434e-19, 3.426237e-19, 3.425712e-19, 3.426078e-19, 3.42594e-19, 
    3.426276e-19, 3.426485e-19, 3.426383e-19, 3.427023e-19, 3.426773e-19, 
    3.428077e-19, 3.427514e-19, 3.429001e-19, 3.428647e-19, 3.429088e-19, 
    3.428864e-19, 3.429244e-19, 3.428903e-19, 3.429501e-19, 3.429627e-19, 
    3.42954e-19, 3.429887e-19, 3.428883e-19, 3.429264e-19, 3.426378e-19, 
    3.426395e-19, 3.426475e-19, 3.426121e-19, 3.426102e-19, 3.42577e-19, 
    3.42607e-19, 3.426188e-19, 3.4265e-19, 3.426677e-19, 3.426849e-19, 
    3.427226e-19, 3.427643e-19, 3.428237e-19, 3.428669e-19, 3.428958e-19, 
    3.428783e-19, 3.428937e-19, 3.428764e-19, 3.428684e-19, 3.429577e-19, 
    3.429073e-19, 3.429837e-19, 3.429796e-19, 3.429447e-19, 3.429801e-19, 
    3.426407e-19, 3.426312e-19, 3.42597e-19, 3.426237e-19, 3.425737e-19, 
    3.426021e-19, 3.42617e-19, 3.42677e-19, 3.426911e-19, 3.42703e-19, 
    3.427273e-19, 3.427582e-19, 3.428122e-19, 3.428598e-19, 3.429039e-19, 
    3.429007e-19, 3.429018e-19, 3.429112e-19, 3.428873e-19, 3.429152e-19, 
    3.429196e-19, 3.429077e-19, 3.42979e-19, 3.429587e-19, 3.429795e-19, 
    3.429663e-19, 3.426343e-19, 3.426505e-19, 3.426417e-19, 3.426581e-19, 
    3.426463e-19, 3.426978e-19, 3.427132e-19, 3.427867e-19, 3.427574e-19, 
    3.42805e-19, 3.427625e-19, 3.427699e-19, 3.42805e-19, 3.427651e-19, 
    3.428565e-19, 3.427932e-19, 3.429116e-19, 3.428468e-19, 3.429156e-19, 
    3.429037e-19, 3.429238e-19, 3.429414e-19, 3.429643e-19, 3.430055e-19, 
    3.429962e-19, 3.430312e-19, 3.42675e-19, 3.426957e-19, 3.426945e-19, 
    3.427167e-19, 3.427329e-19, 3.42769e-19, 3.428261e-19, 3.428049e-19, 
    3.428446e-19, 3.428524e-19, 3.427924e-19, 3.428285e-19, 3.427101e-19, 
    3.427284e-19, 3.42718e-19, 3.426762e-19, 3.428088e-19, 3.427402e-19, 
    3.428675e-19, 3.428305e-19, 3.429388e-19, 3.428842e-19, 3.429908e-19, 
    3.430347e-19, 3.430793e-19, 3.431277e-19, 3.427077e-19, 3.426936e-19, 
    3.427195e-19, 3.427541e-19, 3.427883e-19, 3.428326e-19, 3.428375e-19, 
    3.428457e-19, 3.428675e-19, 3.428855e-19, 3.428475e-19, 3.428901e-19, 
    3.427314e-19, 3.428151e-19, 3.426876e-19, 3.42725e-19, 3.427524e-19, 
    3.427411e-19, 3.428026e-19, 3.428169e-19, 3.428746e-19, 3.428451e-19, 
    3.430233e-19, 3.429442e-19, 3.43167e-19, 3.431041e-19, 3.426885e-19, 
    3.42708e-19, 3.427751e-19, 3.427432e-19, 3.42836e-19, 3.428585e-19, 
    3.428774e-19, 3.429005e-19, 3.429035e-19, 3.429173e-19, 3.428946e-19, 
    3.429167e-19, 3.428327e-19, 3.428703e-19, 3.427682e-19, 3.427926e-19, 
    3.427816e-19, 3.427691e-19, 3.428078e-19, 3.42848e-19, 3.428499e-19, 
    3.428626e-19, 3.428965e-19, 3.428364e-19, 3.430314e-19, 3.429089e-19, 
    3.427292e-19, 3.427654e-19, 3.427719e-19, 3.427576e-19, 3.428562e-19, 
    3.428203e-19, 3.429171e-19, 3.428912e-19, 3.42934e-19, 3.429126e-19, 
    3.429094e-19, 3.428822e-19, 3.42865e-19, 3.428218e-19, 3.427869e-19, 
    3.427598e-19, 3.427662e-19, 3.42796e-19, 3.428507e-19, 3.429033e-19, 
    3.428916e-19, 3.429308e-19, 3.428292e-19, 3.428712e-19, 3.428546e-19, 
    3.428981e-19, 3.42804e-19, 3.428808e-19, 3.427841e-19, 3.427928e-19, 
    3.428196e-19, 3.428733e-19, 3.428868e-19, 3.428993e-19, 3.428918e-19, 
    3.428523e-19, 3.428463e-19, 3.428192e-19, 3.428112e-19, 3.42791e-19, 
    3.427737e-19, 3.427892e-19, 3.428053e-19, 3.428528e-19, 3.42895e-19, 
    3.429415e-19, 3.429533e-19, 3.430051e-19, 3.429614e-19, 3.430319e-19, 
    3.429697e-19, 3.430786e-19, 3.428868e-19, 3.429701e-19, 3.428212e-19, 
    3.428375e-19, 3.428658e-19, 3.429331e-19, 3.428979e-19, 3.429396e-19, 
    3.428462e-19, 3.427965e-19, 3.42785e-19, 3.427612e-19, 3.427855e-19, 
    3.427836e-19, 3.428067e-19, 3.427994e-19, 3.428544e-19, 3.428248e-19, 
    3.42909e-19, 3.429395e-19, 3.430271e-19, 3.430803e-19, 3.431363e-19, 
    3.431605e-19, 3.431679e-19, 3.43171e-19 ;

 MEG_isoprene =
  2.357687e-19, 2.358107e-19, 2.358031e-19, 2.358351e-19, 2.358177e-19, 
    2.358384e-19, 2.357791e-19, 2.35812e-19, 2.357912e-19, 2.357728e-19, 
    2.358961e-19, 2.358366e-19, 2.359617e-19, 2.359231e-19, 2.360213e-19, 
    2.359552e-19, 2.360348e-19, 2.360203e-19, 2.360662e-19, 2.360531e-19, 
    2.361101e-19, 2.360723e-19, 2.361411e-19, 2.361015e-19, 2.361074e-19, 
    2.360709e-19, 2.358494e-19, 2.358884e-19, 2.358469e-19, 2.358525e-19, 
    2.358502e-19, 2.358177e-19, 2.358008e-19, 2.357662e-19, 2.357723e-19, 
    2.357986e-19, 2.35855e-19, 2.358364e-19, 2.358851e-19, 2.35884e-19, 
    2.359377e-19, 2.359134e-19, 2.360044e-19, 2.359787e-19, 2.360537e-19, 
    2.360347e-19, 2.360526e-19, 2.360473e-19, 2.360527e-19, 2.360249e-19, 
    2.360367e-19, 2.360126e-19, 2.359178e-19, 2.359454e-19, 2.358628e-19, 
    2.35812e-19, 2.357804e-19, 2.357554e-19, 2.357587e-19, 2.357647e-19, 
    2.357987e-19, 2.358296e-19, 2.358529e-19, 2.358684e-19, 2.358838e-19, 
    2.359282e-19, 2.359536e-19, 2.360091e-19, 2.359999e-19, 2.360162e-19, 
    2.360328e-19, 2.360598e-19, 2.360555e-19, 2.360672e-19, 2.360163e-19, 
    2.360498e-19, 2.359944e-19, 2.360094e-19, 2.35885e-19, 2.358416e-19, 
    2.358206e-19, 2.358045e-19, 2.357611e-19, 2.357915e-19, 2.357802e-19, 
    2.358077e-19, 2.358247e-19, 2.358164e-19, 2.358689e-19, 2.358483e-19, 
    2.359551e-19, 2.359091e-19, 2.360309e-19, 2.360018e-19, 2.36038e-19, 
    2.360197e-19, 2.360507e-19, 2.360228e-19, 2.360718e-19, 2.360821e-19, 
    2.36075e-19, 2.361034e-19, 2.360212e-19, 2.360523e-19, 2.358161e-19, 
    2.358174e-19, 2.35824e-19, 2.35795e-19, 2.357934e-19, 2.357659e-19, 
    2.357909e-19, 2.358004e-19, 2.35826e-19, 2.358405e-19, 2.358546e-19, 
    2.358855e-19, 2.359196e-19, 2.359683e-19, 2.360037e-19, 2.360273e-19, 
    2.36013e-19, 2.360256e-19, 2.360114e-19, 2.360049e-19, 2.36078e-19, 
    2.360367e-19, 2.360993e-19, 2.360959e-19, 2.360673e-19, 2.360963e-19, 
    2.358184e-19, 2.358106e-19, 2.357826e-19, 2.358045e-19, 2.357631e-19, 
    2.357867e-19, 2.35799e-19, 2.358481e-19, 2.358596e-19, 2.358694e-19, 
    2.358893e-19, 2.359146e-19, 2.359589e-19, 2.359979e-19, 2.360339e-19, 
    2.360313e-19, 2.360322e-19, 2.360399e-19, 2.360203e-19, 2.360432e-19, 
    2.360467e-19, 2.36037e-19, 2.360954e-19, 2.360788e-19, 2.360958e-19, 
    2.36085e-19, 2.358132e-19, 2.358265e-19, 2.358192e-19, 2.358326e-19, 
    2.35823e-19, 2.358651e-19, 2.358778e-19, 2.35938e-19, 2.35914e-19, 
    2.35953e-19, 2.359181e-19, 2.359242e-19, 2.35953e-19, 2.359203e-19, 
    2.359951e-19, 2.359433e-19, 2.360403e-19, 2.359872e-19, 2.360435e-19, 
    2.360337e-19, 2.360502e-19, 2.360647e-19, 2.360834e-19, 2.361172e-19, 
    2.361095e-19, 2.361382e-19, 2.358465e-19, 2.358634e-19, 2.358625e-19, 
    2.358806e-19, 2.358939e-19, 2.359235e-19, 2.359702e-19, 2.359528e-19, 
    2.359854e-19, 2.359918e-19, 2.359426e-19, 2.359722e-19, 2.358752e-19, 
    2.358902e-19, 2.358817e-19, 2.358475e-19, 2.359561e-19, 2.358999e-19, 
    2.360041e-19, 2.359738e-19, 2.360625e-19, 2.360178e-19, 2.361051e-19, 
    2.36141e-19, 2.361775e-19, 2.362172e-19, 2.358733e-19, 2.358617e-19, 
    2.358829e-19, 2.359113e-19, 2.359393e-19, 2.359756e-19, 2.359796e-19, 
    2.359863e-19, 2.360041e-19, 2.360189e-19, 2.359878e-19, 2.360227e-19, 
    2.358927e-19, 2.359612e-19, 2.358568e-19, 2.358874e-19, 2.359099e-19, 
    2.359006e-19, 2.35951e-19, 2.359627e-19, 2.360099e-19, 2.359858e-19, 
    2.361317e-19, 2.360669e-19, 2.362493e-19, 2.361978e-19, 2.358575e-19, 
    2.358735e-19, 2.359285e-19, 2.359023e-19, 2.359783e-19, 2.359968e-19, 
    2.360123e-19, 2.360312e-19, 2.360336e-19, 2.360449e-19, 2.360264e-19, 
    2.360444e-19, 2.359757e-19, 2.360064e-19, 2.359228e-19, 2.359428e-19, 
    2.359338e-19, 2.359235e-19, 2.359552e-19, 2.359881e-19, 2.359897e-19, 
    2.360002e-19, 2.360279e-19, 2.359786e-19, 2.361384e-19, 2.36038e-19, 
    2.358909e-19, 2.359205e-19, 2.359259e-19, 2.359141e-19, 2.359949e-19, 
    2.359655e-19, 2.360448e-19, 2.360235e-19, 2.360586e-19, 2.360411e-19, 
    2.360384e-19, 2.360162e-19, 2.360021e-19, 2.359667e-19, 2.359381e-19, 
    2.359159e-19, 2.359212e-19, 2.359456e-19, 2.359904e-19, 2.360335e-19, 
    2.360239e-19, 2.360559e-19, 2.359728e-19, 2.360071e-19, 2.359935e-19, 
    2.360292e-19, 2.359522e-19, 2.36015e-19, 2.359358e-19, 2.35943e-19, 
    2.359649e-19, 2.360089e-19, 2.360199e-19, 2.360301e-19, 2.36024e-19, 
    2.359917e-19, 2.359868e-19, 2.359646e-19, 2.359581e-19, 2.359415e-19, 
    2.359273e-19, 2.3594e-19, 2.359532e-19, 2.359921e-19, 2.360267e-19, 
    2.360647e-19, 2.360744e-19, 2.361168e-19, 2.36081e-19, 2.361387e-19, 
    2.360878e-19, 2.36177e-19, 2.3602e-19, 2.360881e-19, 2.359662e-19, 
    2.359796e-19, 2.360027e-19, 2.360578e-19, 2.36029e-19, 2.360632e-19, 
    2.359867e-19, 2.35946e-19, 2.359366e-19, 2.359171e-19, 2.35937e-19, 
    2.359354e-19, 2.359544e-19, 2.359483e-19, 2.359934e-19, 2.359692e-19, 
    2.360382e-19, 2.360631e-19, 2.361348e-19, 2.361784e-19, 2.362242e-19, 
    2.36244e-19, 2.362501e-19, 2.362526e-19 ;

 MEG_methanol =
  5.874186e-17, 5.874731e-17, 5.874632e-17, 5.875051e-17, 5.874823e-17, 
    5.875094e-17, 5.874316e-17, 5.874748e-17, 5.874475e-17, 5.87424e-17, 
    5.87585e-17, 5.875071e-17, 5.876711e-17, 5.876204e-17, 5.877491e-17, 
    5.876625e-17, 5.877669e-17, 5.877478e-17, 5.87808e-17, 5.877908e-17, 
    5.878655e-17, 5.87816e-17, 5.879062e-17, 5.878543e-17, 5.87862e-17, 
    5.878142e-17, 5.875238e-17, 5.87575e-17, 5.875206e-17, 5.875279e-17, 
    5.875249e-17, 5.874823e-17, 5.874602e-17, 5.874154e-17, 5.874234e-17, 
    5.874572e-17, 5.875312e-17, 5.875068e-17, 5.875706e-17, 5.875692e-17, 
    5.876396e-17, 5.876077e-17, 5.87727e-17, 5.876934e-17, 5.877916e-17, 
    5.877667e-17, 5.877902e-17, 5.877832e-17, 5.877903e-17, 5.877538e-17, 
    5.877694e-17, 5.877377e-17, 5.876134e-17, 5.876496e-17, 5.875414e-17, 
    5.874747e-17, 5.874334e-17, 5.874013e-17, 5.874056e-17, 5.874134e-17, 
    5.874574e-17, 5.874979e-17, 5.875285e-17, 5.875488e-17, 5.87569e-17, 
    5.876271e-17, 5.876605e-17, 5.877332e-17, 5.87721e-17, 5.877424e-17, 
    5.877642e-17, 5.877996e-17, 5.877939e-17, 5.878093e-17, 5.877426e-17, 
    5.877865e-17, 5.877139e-17, 5.877336e-17, 5.875705e-17, 5.875136e-17, 
    5.874861e-17, 5.874649e-17, 5.874087e-17, 5.874479e-17, 5.874331e-17, 
    5.874692e-17, 5.874915e-17, 5.874806e-17, 5.875494e-17, 5.875224e-17, 
    5.876624e-17, 5.87602e-17, 5.877617e-17, 5.877236e-17, 5.87771e-17, 
    5.87747e-17, 5.877878e-17, 5.877511e-17, 5.878153e-17, 5.878289e-17, 
    5.878195e-17, 5.878567e-17, 5.877489e-17, 5.877898e-17, 5.874801e-17, 
    5.874819e-17, 5.874905e-17, 5.874526e-17, 5.874504e-17, 5.87415e-17, 
    5.874471e-17, 5.874596e-17, 5.874931e-17, 5.875122e-17, 5.875306e-17, 
    5.875711e-17, 5.876159e-17, 5.876796e-17, 5.877261e-17, 5.87757e-17, 
    5.877383e-17, 5.877548e-17, 5.877362e-17, 5.877276e-17, 5.878235e-17, 
    5.877693e-17, 5.878514e-17, 5.87847e-17, 5.878095e-17, 5.878475e-17, 
    5.874832e-17, 5.87473e-17, 5.874363e-17, 5.87465e-17, 5.874114e-17, 
    5.874417e-17, 5.874578e-17, 5.875222e-17, 5.875373e-17, 5.8755e-17, 
    5.875762e-17, 5.876093e-17, 5.876674e-17, 5.877184e-17, 5.877657e-17, 
    5.877623e-17, 5.877634e-17, 5.877736e-17, 5.877479e-17, 5.877779e-17, 
    5.877825e-17, 5.877698e-17, 5.878464e-17, 5.878245e-17, 5.878469e-17, 
    5.878327e-17, 5.874764e-17, 5.874938e-17, 5.874843e-17, 5.875019e-17, 
    5.874892e-17, 5.875445e-17, 5.875611e-17, 5.876399e-17, 5.876085e-17, 
    5.876595e-17, 5.87614e-17, 5.876219e-17, 5.876596e-17, 5.876167e-17, 
    5.877149e-17, 5.876468e-17, 5.87774e-17, 5.877044e-17, 5.877783e-17, 
    5.877655e-17, 5.877871e-17, 5.87806e-17, 5.878306e-17, 5.878748e-17, 
    5.878648e-17, 5.879024e-17, 5.875201e-17, 5.875422e-17, 5.87541e-17, 
    5.875648e-17, 5.875822e-17, 5.87621e-17, 5.876822e-17, 5.876594e-17, 
    5.877021e-17, 5.877104e-17, 5.87646e-17, 5.876848e-17, 5.875576e-17, 
    5.875774e-17, 5.875662e-17, 5.875214e-17, 5.876637e-17, 5.875901e-17, 
    5.877266e-17, 5.876869e-17, 5.878032e-17, 5.877446e-17, 5.87859e-17, 
    5.879061e-17, 5.87954e-17, 5.88006e-17, 5.875551e-17, 5.8754e-17, 
    5.875678e-17, 5.87605e-17, 5.876417e-17, 5.876892e-17, 5.876945e-17, 
    5.877032e-17, 5.877266e-17, 5.87746e-17, 5.877052e-17, 5.877509e-17, 
    5.875805e-17, 5.876704e-17, 5.875336e-17, 5.875737e-17, 5.876031e-17, 
    5.875909e-17, 5.87657e-17, 5.876723e-17, 5.877343e-17, 5.877026e-17, 
    5.878939e-17, 5.87809e-17, 5.880481e-17, 5.879806e-17, 5.875345e-17, 
    5.875555e-17, 5.876275e-17, 5.875932e-17, 5.876928e-17, 5.87717e-17, 
    5.877373e-17, 5.877621e-17, 5.877654e-17, 5.877801e-17, 5.877558e-17, 
    5.877795e-17, 5.876893e-17, 5.877297e-17, 5.876201e-17, 5.876463e-17, 
    5.876345e-17, 5.87621e-17, 5.876626e-17, 5.877057e-17, 5.877078e-17, 
    5.877214e-17, 5.877578e-17, 5.876932e-17, 5.879026e-17, 5.877711e-17, 
    5.875782e-17, 5.876171e-17, 5.876241e-17, 5.876087e-17, 5.877145e-17, 
    5.87676e-17, 5.877799e-17, 5.877521e-17, 5.877981e-17, 5.877751e-17, 
    5.877716e-17, 5.877425e-17, 5.87724e-17, 5.876775e-17, 5.876402e-17, 
    5.87611e-17, 5.87618e-17, 5.876499e-17, 5.877086e-17, 5.877651e-17, 
    5.877525e-17, 5.877945e-17, 5.876856e-17, 5.877306e-17, 5.877128e-17, 
    5.877595e-17, 5.876586e-17, 5.877409e-17, 5.876371e-17, 5.876464e-17, 
    5.876753e-17, 5.877329e-17, 5.877474e-17, 5.877607e-17, 5.877527e-17, 
    5.877103e-17, 5.877039e-17, 5.876748e-17, 5.876662e-17, 5.876445e-17, 
    5.876259e-17, 5.876426e-17, 5.876599e-17, 5.877108e-17, 5.877562e-17, 
    5.878061e-17, 5.878188e-17, 5.878743e-17, 5.878275e-17, 5.879031e-17, 
    5.878364e-17, 5.879533e-17, 5.877474e-17, 5.878368e-17, 5.87677e-17, 
    5.876944e-17, 5.877248e-17, 5.877971e-17, 5.877593e-17, 5.87804e-17, 
    5.877038e-17, 5.876504e-17, 5.876381e-17, 5.876126e-17, 5.876386e-17, 
    5.876366e-17, 5.876614e-17, 5.876535e-17, 5.877126e-17, 5.876809e-17, 
    5.877712e-17, 5.878039e-17, 5.87898e-17, 5.879551e-17, 5.880152e-17, 
    5.880411e-17, 5.880491e-17, 5.880524e-17 ;

 MEG_pinene_a =
  4.866617e-17, 4.867125e-17, 4.867032e-17, 4.867422e-17, 4.86721e-17, 
    4.867462e-17, 4.86674e-17, 4.86714e-17, 4.866887e-17, 4.866668e-17, 
    4.868164e-17, 4.86744e-17, 4.868963e-17, 4.868493e-17, 4.869689e-17, 
    4.868884e-17, 4.869854e-17, 4.869677e-17, 4.870236e-17, 4.870076e-17, 
    4.87077e-17, 4.87031e-17, 4.871148e-17, 4.870666e-17, 4.870737e-17, 
    4.870293e-17, 4.867596e-17, 4.868071e-17, 4.867565e-17, 4.867634e-17, 
    4.867606e-17, 4.86721e-17, 4.867004e-17, 4.866587e-17, 4.866661e-17, 
    4.866977e-17, 4.867665e-17, 4.867438e-17, 4.86803e-17, 4.868017e-17, 
    4.868671e-17, 4.868375e-17, 4.869483e-17, 4.869171e-17, 4.870083e-17, 
    4.869852e-17, 4.870071e-17, 4.870006e-17, 4.870071e-17, 4.869733e-17, 
    4.869877e-17, 4.869582e-17, 4.868428e-17, 4.868764e-17, 4.867759e-17, 
    4.86714e-17, 4.866756e-17, 4.866456e-17, 4.866495e-17, 4.866569e-17, 
    4.866979e-17, 4.867355e-17, 4.867639e-17, 4.867828e-17, 4.868015e-17, 
    4.868555e-17, 4.868865e-17, 4.869541e-17, 4.869428e-17, 4.869626e-17, 
    4.869829e-17, 4.870158e-17, 4.870105e-17, 4.870248e-17, 4.869628e-17, 
    4.870036e-17, 4.869361e-17, 4.869545e-17, 4.86803e-17, 4.867501e-17, 
    4.867245e-17, 4.867049e-17, 4.866525e-17, 4.866891e-17, 4.866753e-17, 
    4.867088e-17, 4.867295e-17, 4.867195e-17, 4.867833e-17, 4.867583e-17, 
    4.868883e-17, 4.868323e-17, 4.869805e-17, 4.869452e-17, 4.869892e-17, 
    4.869669e-17, 4.870048e-17, 4.869707e-17, 4.870303e-17, 4.87043e-17, 
    4.870343e-17, 4.870689e-17, 4.869687e-17, 4.870067e-17, 4.86719e-17, 
    4.867206e-17, 4.867286e-17, 4.866934e-17, 4.866914e-17, 4.866583e-17, 
    4.866883e-17, 4.867e-17, 4.867311e-17, 4.867488e-17, 4.867659e-17, 
    4.868035e-17, 4.868451e-17, 4.869043e-17, 4.869474e-17, 4.869762e-17, 
    4.869588e-17, 4.869741e-17, 4.869569e-17, 4.869489e-17, 4.87038e-17, 
    4.869876e-17, 4.870639e-17, 4.870598e-17, 4.87025e-17, 4.870603e-17, 
    4.867218e-17, 4.867123e-17, 4.866783e-17, 4.867049e-17, 4.866549e-17, 
    4.866833e-17, 4.866982e-17, 4.86758e-17, 4.867721e-17, 4.867839e-17, 
    4.868082e-17, 4.86839e-17, 4.868929e-17, 4.869403e-17, 4.869843e-17, 
    4.869811e-17, 4.869822e-17, 4.869916e-17, 4.869677e-17, 4.869956e-17, 
    4.869999e-17, 4.869881e-17, 4.870592e-17, 4.870389e-17, 4.870597e-17, 
    4.870466e-17, 4.867155e-17, 4.867316e-17, 4.867229e-17, 4.867392e-17, 
    4.867274e-17, 4.867788e-17, 4.867941e-17, 4.868674e-17, 4.868382e-17, 
    4.868857e-17, 4.868433e-17, 4.868506e-17, 4.868857e-17, 4.868459e-17, 
    4.86937e-17, 4.868739e-17, 4.86992e-17, 4.869273e-17, 4.86996e-17, 
    4.869841e-17, 4.870041e-17, 4.870217e-17, 4.870446e-17, 4.870857e-17, 
    4.870763e-17, 4.871113e-17, 4.867561e-17, 4.867767e-17, 4.867755e-17, 
    4.867976e-17, 4.868138e-17, 4.868498e-17, 4.869067e-17, 4.868855e-17, 
    4.869252e-17, 4.869329e-17, 4.868731e-17, 4.869091e-17, 4.86791e-17, 
    4.868093e-17, 4.867989e-17, 4.867573e-17, 4.868895e-17, 4.868211e-17, 
    4.86948e-17, 4.869111e-17, 4.870191e-17, 4.869647e-17, 4.87071e-17, 
    4.871148e-17, 4.871592e-17, 4.872075e-17, 4.867887e-17, 4.867746e-17, 
    4.868004e-17, 4.86835e-17, 4.86869e-17, 4.869132e-17, 4.869181e-17, 
    4.869262e-17, 4.86948e-17, 4.86966e-17, 4.869281e-17, 4.869706e-17, 
    4.868122e-17, 4.868957e-17, 4.867686e-17, 4.868059e-17, 4.868332e-17, 
    4.868219e-17, 4.868833e-17, 4.868975e-17, 4.86955e-17, 4.869257e-17, 
    4.871033e-17, 4.870245e-17, 4.872467e-17, 4.871839e-17, 4.867695e-17, 
    4.867889e-17, 4.868558e-17, 4.86824e-17, 4.869165e-17, 4.86939e-17, 
    4.869579e-17, 4.869809e-17, 4.869839e-17, 4.869977e-17, 4.869751e-17, 
    4.86997e-17, 4.869133e-17, 4.869508e-17, 4.86849e-17, 4.868733e-17, 
    4.868624e-17, 4.868498e-17, 4.868885e-17, 4.869285e-17, 4.869305e-17, 
    4.869432e-17, 4.869769e-17, 4.86917e-17, 4.871115e-17, 4.869893e-17, 
    4.868101e-17, 4.868462e-17, 4.868527e-17, 4.868384e-17, 4.869367e-17, 
    4.869009e-17, 4.869975e-17, 4.869716e-17, 4.870143e-17, 4.86993e-17, 
    4.869898e-17, 4.869627e-17, 4.869455e-17, 4.869024e-17, 4.868677e-17, 
    4.868406e-17, 4.86847e-17, 4.868767e-17, 4.869312e-17, 4.869837e-17, 
    4.86972e-17, 4.870111e-17, 4.869098e-17, 4.869517e-17, 4.869351e-17, 
    4.869785e-17, 4.868847e-17, 4.869612e-17, 4.868648e-17, 4.868735e-17, 
    4.869002e-17, 4.869537e-17, 4.869672e-17, 4.869797e-17, 4.869722e-17, 
    4.869328e-17, 4.869268e-17, 4.868999e-17, 4.868919e-17, 4.868717e-17, 
    4.868544e-17, 4.868699e-17, 4.86886e-17, 4.869333e-17, 4.869754e-17, 
    4.870218e-17, 4.870336e-17, 4.870852e-17, 4.870417e-17, 4.871119e-17, 
    4.870499e-17, 4.871586e-17, 4.869673e-17, 4.870503e-17, 4.869018e-17, 
    4.869181e-17, 4.869463e-17, 4.870134e-17, 4.869783e-17, 4.870199e-17, 
    4.869267e-17, 4.868772e-17, 4.868657e-17, 4.86842e-17, 4.868663e-17, 
    4.868643e-17, 4.868874e-17, 4.8688e-17, 4.869349e-17, 4.869055e-17, 
    4.869894e-17, 4.870198e-17, 4.871072e-17, 4.871602e-17, 4.872161e-17, 
    4.872402e-17, 4.872476e-17, 4.872506e-17 ;

 MEG_thujene_a =
  1.227203e-18, 1.227327e-18, 1.227305e-18, 1.227399e-18, 1.227348e-18, 
    1.227409e-18, 1.227233e-18, 1.227331e-18, 1.227269e-18, 1.227216e-18, 
    1.22758e-18, 1.227404e-18, 1.227774e-18, 1.227659e-18, 1.22795e-18, 
    1.227754e-18, 1.22799e-18, 1.227947e-18, 1.228083e-18, 1.228044e-18, 
    1.228213e-18, 1.228101e-18, 1.228305e-18, 1.228188e-18, 1.228205e-18, 
    1.228097e-18, 1.227441e-18, 1.227557e-18, 1.227434e-18, 1.227451e-18, 
    1.227444e-18, 1.227348e-18, 1.227298e-18, 1.227196e-18, 1.227214e-18, 
    1.227291e-18, 1.227458e-18, 1.227403e-18, 1.227547e-18, 1.227544e-18, 
    1.227703e-18, 1.227631e-18, 1.2279e-18, 1.227824e-18, 1.228046e-18, 
    1.22799e-18, 1.228043e-18, 1.228027e-18, 1.228043e-18, 1.227961e-18, 
    1.227996e-18, 1.227924e-18, 1.227644e-18, 1.227725e-18, 1.227481e-18, 
    1.227331e-18, 1.227237e-18, 1.227164e-18, 1.227174e-18, 1.227192e-18, 
    1.227291e-18, 1.227383e-18, 1.227452e-18, 1.227498e-18, 1.227543e-18, 
    1.227675e-18, 1.22775e-18, 1.227914e-18, 1.227887e-18, 1.227935e-18, 
    1.227984e-18, 1.228064e-18, 1.228051e-18, 1.228086e-18, 1.227935e-18, 
    1.228035e-18, 1.227871e-18, 1.227915e-18, 1.227547e-18, 1.227418e-18, 
    1.227356e-18, 1.227308e-18, 1.227181e-18, 1.22727e-18, 1.227237e-18, 
    1.227318e-18, 1.227368e-18, 1.227344e-18, 1.227499e-18, 1.227438e-18, 
    1.227754e-18, 1.227618e-18, 1.227978e-18, 1.227892e-18, 1.227999e-18, 
    1.227945e-18, 1.228037e-18, 1.227954e-18, 1.228099e-18, 1.22813e-18, 
    1.228109e-18, 1.228193e-18, 1.22795e-18, 1.228042e-18, 1.227343e-18, 
    1.227347e-18, 1.227366e-18, 1.22728e-18, 1.227276e-18, 1.227195e-18, 
    1.227268e-18, 1.227297e-18, 1.227372e-18, 1.227415e-18, 1.227457e-18, 
    1.227548e-18, 1.227649e-18, 1.227793e-18, 1.227898e-18, 1.227968e-18, 
    1.227926e-18, 1.227963e-18, 1.227921e-18, 1.227902e-18, 1.228118e-18, 
    1.227996e-18, 1.228181e-18, 1.228171e-18, 1.228086e-18, 1.228172e-18, 
    1.22735e-18, 1.227327e-18, 1.227244e-18, 1.227309e-18, 1.227187e-18, 
    1.227256e-18, 1.227292e-18, 1.227438e-18, 1.227472e-18, 1.227501e-18, 
    1.22756e-18, 1.227634e-18, 1.227765e-18, 1.227881e-18, 1.227987e-18, 
    1.22798e-18, 1.227982e-18, 1.228005e-18, 1.227947e-18, 1.228015e-18, 
    1.228026e-18, 1.227997e-18, 1.22817e-18, 1.22812e-18, 1.228171e-18, 
    1.228139e-18, 1.227334e-18, 1.227373e-18, 1.227352e-18, 1.227392e-18, 
    1.227363e-18, 1.227488e-18, 1.227525e-18, 1.227704e-18, 1.227632e-18, 
    1.227748e-18, 1.227645e-18, 1.227663e-18, 1.227748e-18, 1.227651e-18, 
    1.227873e-18, 1.227719e-18, 1.228006e-18, 1.227849e-18, 1.228016e-18, 
    1.227987e-18, 1.228036e-18, 1.228079e-18, 1.228134e-18, 1.228234e-18, 
    1.228211e-18, 1.228296e-18, 1.227433e-18, 1.227483e-18, 1.22748e-18, 
    1.227534e-18, 1.227573e-18, 1.227661e-18, 1.227799e-18, 1.227747e-18, 
    1.227844e-18, 1.227863e-18, 1.227717e-18, 1.227805e-18, 1.227518e-18, 
    1.227562e-18, 1.227537e-18, 1.227436e-18, 1.227757e-18, 1.227591e-18, 
    1.227899e-18, 1.22781e-18, 1.228072e-18, 1.22794e-18, 1.228198e-18, 
    1.228305e-18, 1.228413e-18, 1.22853e-18, 1.227512e-18, 1.227478e-18, 
    1.227541e-18, 1.227625e-18, 1.227707e-18, 1.227815e-18, 1.227827e-18, 
    1.227846e-18, 1.227899e-18, 1.227943e-18, 1.227851e-18, 1.227954e-18, 
    1.227569e-18, 1.227772e-18, 1.227463e-18, 1.227554e-18, 1.22762e-18, 
    1.227593e-18, 1.227742e-18, 1.227777e-18, 1.227916e-18, 1.227845e-18, 
    1.228277e-18, 1.228085e-18, 1.228625e-18, 1.228473e-18, 1.227466e-18, 
    1.227513e-18, 1.227675e-18, 1.227598e-18, 1.227823e-18, 1.227877e-18, 
    1.227923e-18, 1.227979e-18, 1.227987e-18, 1.22802e-18, 1.227965e-18, 
    1.228018e-18, 1.227815e-18, 1.227906e-18, 1.227659e-18, 1.227718e-18, 
    1.227691e-18, 1.227661e-18, 1.227755e-18, 1.227852e-18, 1.227857e-18, 
    1.227888e-18, 1.22797e-18, 1.227824e-18, 1.228297e-18, 1.228e-18, 
    1.227564e-18, 1.227652e-18, 1.227668e-18, 1.227633e-18, 1.227872e-18, 
    1.227785e-18, 1.22802e-18, 1.227957e-18, 1.22806e-18, 1.228009e-18, 
    1.228001e-18, 1.227935e-18, 1.227893e-18, 1.227788e-18, 1.227704e-18, 
    1.227638e-18, 1.227654e-18, 1.227726e-18, 1.227859e-18, 1.227986e-18, 
    1.227958e-18, 1.228053e-18, 1.227806e-18, 1.227908e-18, 1.227868e-18, 
    1.227973e-18, 1.227746e-18, 1.227931e-18, 1.227697e-18, 1.227718e-18, 
    1.227783e-18, 1.227913e-18, 1.227946e-18, 1.227976e-18, 1.227958e-18, 
    1.227862e-18, 1.227848e-18, 1.227782e-18, 1.227763e-18, 1.227714e-18, 
    1.227672e-18, 1.22771e-18, 1.227749e-18, 1.227864e-18, 1.227966e-18, 
    1.228079e-18, 1.228107e-18, 1.228233e-18, 1.228127e-18, 1.228298e-18, 
    1.228147e-18, 1.228411e-18, 1.227946e-18, 1.228148e-18, 1.227787e-18, 
    1.227827e-18, 1.227895e-18, 1.228058e-18, 1.227973e-18, 1.228074e-18, 
    1.227848e-18, 1.227727e-18, 1.227699e-18, 1.227642e-18, 1.227701e-18, 
    1.227696e-18, 1.227752e-18, 1.227734e-18, 1.227867e-18, 1.227796e-18, 
    1.228e-18, 1.228074e-18, 1.228286e-18, 1.228415e-18, 1.228551e-18, 
    1.228609e-18, 1.228627e-18, 1.228635e-18 ;

 MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 M_LITR1C_TO_LEACHING =
  7.96638e-26, -2.939316e-25, 1.593275e-25, 1.730626e-25, 8.241157e-27, 
    -1.867976e-25, 8.515785e-26, 1.977859e-25, -3.488721e-25, -5.768744e-26, 
    2.060269e-25, -7.691661e-26, 2.334972e-25, -2.747016e-26, 8.790487e-26, 
    1.950388e-25, -1.867976e-25, -4.999584e-25, -1.373504e-26, 4.944653e-26, 
    -9.614578e-26, 2.225091e-25, -4.58753e-25, 3.049198e-25, 1.922926e-26, 
    3.57114e-26, -9.614578e-26, -3.571124e-26, 2.747107e-27, -1.922909e-26, 
    -4.395231e-26, -5.493967e-27, -9.065174e-26, 1.208692e-25, 2.692085e-25, 
    5.494132e-27, 9.614595e-26, -2.225089e-25, 2.719555e-25, -2.417381e-25, 
    1.675686e-25, 1.703156e-25, 4.120545e-26, -1.785565e-25, 5.494058e-26, 
    3.296438e-26, 4.752353e-25, -2.527262e-25, -7.691661e-26, 2.747033e-26, 
    4.697413e-25, -4.367769e-25, -3.159078e-25, -3.516191e-25, 8.790487e-26, 
    -1.922909e-26, -2.417381e-25, -7.966364e-26, 4.3403e-25, -4.779822e-25, 
    -1.373504e-26, -2.746942e-27, -3.845826e-26, -1.785565e-25, 
    -4.944644e-25, -1.895446e-25, -2.472314e-26, -3.214018e-25, 
    -8.240992e-27, 2.911847e-25, -4.395231e-26, 3.296438e-26, -2.966786e-25, 
    -1.730625e-25, 2.527264e-25, 1.895448e-25, 3.845843e-26, -3.928245e-25, 
    -2.060268e-25, 5.52152e-25, 1.648223e-26, -4.312828e-25, -1.867976e-25, 
    -4.669934e-26, 1.373521e-26, -1.785565e-25, 6.263217e-25, 5.76876e-26, 
    9.614595e-26, -4.944636e-26, -3.845826e-26, 2.472323e-25, 1.455924e-25, 
    7.416975e-26, 9.889298e-26, -5.219339e-26, -2.3075e-25, -2.3075e-25, 
    2.197628e-26, 3.378841e-25, -8.240992e-27, -1.922909e-26, -1.703155e-25, 
    -2.554732e-25, -2.692083e-25, -5.494041e-26, -2.005327e-25, 
    -2.609673e-25, -1.20869e-25, 3.763425e-25, 8.257326e-32, -2.087738e-25, 
    -5.219339e-26, -3.928245e-25, 2.856907e-25, -3.021727e-25, -1.263631e-25, 
    -2.142679e-25, 4.944653e-26, -8.790471e-26, 1.675686e-25, -1.703155e-25, 
    -1.977857e-25, -1.23616e-25, -2.060268e-25, 3.983187e-25, -3.296421e-26, 
    -4.944644e-25, 1.648223e-26, 1.263632e-25, 9.06519e-26, 4.862235e-25, 
    -5.493967e-27, -4.395239e-25, 6.592867e-26, 1.593275e-25, -3.653542e-25, 
    2.747026e-25, 3.406311e-25, -3.40631e-25, -5.164406e-25, -9.614578e-26, 
    1.153751e-25, -4.340298e-25, 1.785567e-25, -2.197612e-26, -4.093066e-25, 
    -2.36244e-25, 4.36777e-25, -4.56006e-25, -3.268959e-25, 2.747107e-27, 
    1.867978e-25, 4.477651e-25, 5.494058e-26, -2.3075e-25, 1.181221e-25, 
    1.593275e-25, -1.373512e-25, 1.703156e-25, -4.367769e-25, -2.28003e-25, 
    7.96638e-26, 1.977859e-25, 5.494058e-26, -1.23616e-25, 9.339892e-26, 
    1.208692e-25, 3.543663e-25, 1.538335e-25, 2.389912e-25, -3.488721e-25, 
    4.862235e-25, 2.472323e-25, -1.18122e-25, -4.065596e-25, -3.159078e-25, 
    -3.323899e-25, -3.598602e-25, -3.873304e-25, 2.197628e-26, -4.395231e-26, 
    4.120545e-26, -1.538333e-25, 3.406311e-25, 1.758097e-25, -9.339876e-26, 
    -1.758095e-25, -1.20869e-25, -3.735953e-25, -5.576459e-25, -3.543661e-25, 
    -1.840506e-25, -1.428452e-25, 8.241157e-27, 5.494058e-26, -7.142256e-26, 
    1.428454e-25, 1.428454e-25, 2.911847e-25, 2.911847e-25, 2.472323e-25, 
    2.197628e-26, 3.790895e-25, 2.637145e-25, -3.104137e-25, -1.785565e-25, 
    3.900776e-25, -3.845826e-26, -2.856905e-25, 2.747026e-25, -1.867976e-25, 
    -9.339876e-26, 3.790895e-25, 1.922926e-26, -2.472321e-25, 8.241083e-26, 
    -4.972114e-25, 2.554734e-25, -4.422709e-25, -1.098802e-26, 2.14268e-25, 
    -2.472321e-25, -2.609673e-25, -4.148007e-25, -1.15375e-25, 2.582204e-25, 
    -1.648214e-25, -6.043446e-26, -2.801964e-25, -2.582203e-25, 
    -1.428452e-25, -1.785565e-25, -1.758095e-25, 2.527264e-25, -1.016398e-25, 
    -1.648207e-26, -2.747016e-26, 1.593275e-25, 1.867978e-25, 1.455924e-25, 
    -3.021727e-25, 1.895448e-25, -2.225089e-25, 6.043463e-26, -9.339876e-26, 
    -5.219339e-26, -4.312828e-25, -3.571131e-25, -7.142256e-26, 7.691677e-26, 
    -1.538333e-25, -1.483393e-25, -3.653542e-25, 1.428454e-25, 5.494058e-26, 
    9.339892e-26, -1.18122e-25, 5.43911e-25, -5.823692e-25, 1.181221e-25, 
    -2.582203e-25, -8.241066e-26, -3.296429e-25, 1.318573e-25, -4.010655e-25, 
    -7.691661e-26, 6.592867e-26, 3.57114e-26, 1.04387e-25, 7.96638e-26, 
    8.25715e-32, -3.37884e-25, -2.911845e-25, -3.818364e-25, 1.538335e-25, 
    5.494132e-27, -1.593274e-25, 1.373521e-26, 3.845835e-25, 5.768753e-25, 
    4.944653e-26, -5.219339e-26, -1.071339e-25, -2.527262e-25, -5.054525e-25, 
    1.153751e-25, 2.005329e-25, 2.774496e-25, -1.455922e-25, 4.66995e-26, 
    -1.15375e-25, -4.065596e-25, 4.972116e-25, -3.955715e-25, -2.197612e-26, 
    5.76876e-26, 1.153751e-25, -1.950387e-25, 9.614595e-26, -2.060268e-25, 
    -9.065174e-26, 4.66995e-26, 3.21402e-25, 4.120545e-26, -3.159078e-25, 
    -1.016398e-25, 1.428454e-25, -4.202947e-25, 8.257051e-32, 2.444853e-25, 
    7.554319e-25, -1.758095e-25, 5.219355e-26, 1.236162e-25, -4.477649e-25, 
    2.444853e-25, 1.153751e-25, 7.416975e-26, -2.747016e-26, 3.076668e-25, 
    5.494058e-26, -1.483393e-25, 7.691677e-26, 3.708484e-25, 7.142273e-26, 
    -2.692083e-25, -2.746942e-27, 1.565805e-25, -3.241488e-25, -1.071339e-25, 
    -3.049197e-25, -5.494041e-26, -9.889281e-26, -3.296429e-25, 
    -3.296421e-26, -8.515768e-26, -7.142256e-26 ;

 M_LITR2C_TO_LEACHING =
  -2.747024e-25, 1.758096e-25, -9.889284e-26, -2.582203e-25, -1.291101e-25, 
    -8.790474e-26, 2.197625e-26, -1.895447e-25, 1.840507e-25, 1.510864e-25, 
    2.14268e-25, -2.060268e-25, -1.098809e-25, 7.691675e-26, -1.483393e-25, 
    -1.15375e-25, -9.889284e-26, 1.785567e-25, 1.291102e-25, -1.098809e-25, 
    -1.648209e-26, -1.263631e-25, 5.494103e-27, 1.373513e-25, 4.94465e-26, 
    -1.950387e-25, 2.829436e-25, -1.346042e-25, 4.120543e-26, -3.40631e-25, 
    8.515782e-26, -2.747024e-25, 1.126281e-25, -2.087738e-25, 3.84584e-26, 
    9.065187e-26, 2.334972e-25, -1.20869e-25, 1.04387e-25, 2.801966e-25, 
    -2.005328e-25, 1.153751e-25, 1.703156e-25, -3.186548e-25, -2.801965e-25, 
    -1.593274e-25, -5.493996e-27, -1.840506e-25, -7.142259e-26, 
    -2.994256e-25, 3.021733e-26, -4.669937e-26, 9.889295e-26, -1.840506e-25, 
    -6.867557e-26, -1.263631e-25, 3.159079e-25, 2.362442e-25, 1.098815e-26, 
    3.296435e-26, -6.592854e-26, -3.873304e-25, 8.241128e-27, 1.483394e-25, 
    -9.339879e-26, 1.0164e-25, -1.977857e-25, -1.922917e-25, 1.483394e-25, 
    3.84584e-26, -8.515771e-26, 1.922923e-26, -3.296429e-25, 1.428453e-25, 
    -2.3075e-25, -1.648214e-25, -4.395234e-26, -5.768747e-26, -3.818364e-25, 
    2.417382e-25, -3.571127e-26, 3.900776e-25, 7.14227e-26, 1.483394e-25, 
    -9.614581e-26, 2.032799e-25, -5.494044e-26, 1.318572e-25, -1.236161e-25, 
    -1.758095e-25, 4.285359e-25, -1.318571e-25, -1.043869e-25, 4.669947e-26, 
    1.510864e-25, -2.444852e-25, -4.395234e-26, -1.538333e-25, 8.790485e-26, 
    -1.071339e-25, -3.186548e-25, 5.219352e-26, -2.225089e-25, 5.494103e-27, 
    -6.867557e-26, 2.74703e-26, -9.339879e-26, -1.098805e-26, -1.648214e-25, 
    -1.867976e-25, -8.515771e-26, -1.15375e-25, 1.236162e-25, 9.614592e-26, 
    -7.691664e-26, 2.280031e-25, 6.04346e-26, 3.84584e-26, -4.944639e-26, 
    1.922923e-26, -1.15375e-25, 7.691675e-26, -1.016399e-25, 1.703156e-25, 
    -3.021722e-26, -1.12628e-25, -2.719554e-25, 1.181221e-25, 1.09881e-25, 
    1.153751e-25, -3.845829e-26, -9.339879e-26, -9.339879e-26, 1.09881e-25, 
    -2.142679e-25, 1.675686e-25, -5.493996e-27, 5.494103e-27, -1.15375e-25, 
    -8.241069e-26, 2.14268e-25, -1.813036e-25, 1.510864e-25, -6.043449e-26, 
    -1.318571e-25, -2.417381e-25, -1.20869e-25, -1.867976e-25, -1.428452e-25, 
    -1.016399e-25, -1.538333e-25, -2.197614e-26, -3.296424e-26, 
    -2.005328e-25, 1.09881e-25, -3.543661e-25, -2.719554e-25, 9.339889e-26, 
    -5.494044e-26, 2.527263e-25, 8.790485e-26, -8.241069e-26, -8.790474e-26, 
    4.120543e-26, -2.74702e-26, -3.241489e-25, -1.236161e-25, 1.64822e-26, 
    -2.005328e-25, -2.115208e-25, -2.197614e-26, -2.472322e-25, 
    -7.142259e-26, -6.318152e-26, -2.994256e-25, -2.637143e-25, 2.74703e-26, 
    -1.043869e-25, 4.669947e-26, -3.571127e-26, -3.296424e-26, -2.3075e-25, 
    -1.098809e-25, -5.494044e-26, -1.593274e-25, 8.241128e-27, -9.339879e-26, 
    2.74703e-26, 3.296435e-26, 2.994258e-25, 2.087739e-25, -6.043449e-26, 
    1.153751e-25, 1.977858e-25, -1.538333e-25, -3.076667e-25, 1.922918e-25, 
    1.236162e-25, 1.181221e-25, -1.043869e-25, 1.318572e-25, 1.318572e-25, 
    -1.016399e-25, -3.571127e-26, 3.296435e-26, -7.142259e-26, 1.840507e-25, 
    -3.296424e-26, -2.719554e-25, -3.626072e-25, -8.515771e-26, 
    -2.692084e-25, -1.263631e-25, 1.64822e-26, -4.944639e-26, -1.758095e-25, 
    -7.142259e-26, -2.28003e-25, -1.20869e-25, 6.592865e-26, 1.428453e-25, 
    -2.032798e-25, 1.04387e-25, 1.785567e-25, -9.889284e-26, 5.219352e-26, 
    -1.016399e-25, -2.087738e-25, -1.373512e-25, -3.296424e-26, -1.20869e-25, 
    -1.867976e-25, 1.373518e-26, 4.669947e-26, -1.510863e-25, -4.010656e-25, 
    -1.263631e-25, 5.494103e-27, -1.867976e-25, 1.977858e-25, 7.691675e-26, 
    -9.614581e-26, -1.15375e-25, -3.296424e-26, -3.598602e-25, -1.236161e-25, 
    -1.098805e-26, -1.758095e-25, 2.087739e-25, -6.592854e-26, -1.703155e-25, 
    3.131609e-25, 3.516192e-25, 1.09881e-25, -1.483393e-25, 8.24108e-26, 
    1.620745e-25, -1.867976e-25, -1.977857e-25, -2.692084e-25, -1.922917e-25, 
    5.494055e-26, 1.593275e-25, -1.510863e-25, -2.170149e-25, -1.510863e-25, 
    -1.922912e-26, 2.225091e-25, 1.922918e-25, -1.098809e-25, 4.175478e-25, 
    -1.373512e-25, -1.922912e-26, 5.494103e-27, 9.889295e-26, -1.263631e-25, 
    -5.493996e-27, -1.098809e-25, -9.339879e-26, -9.889284e-26, 
    -1.922912e-26, 1.758096e-25, 1.840507e-25, -1.648214e-25, -6.043449e-26, 
    -9.889284e-26, -1.648214e-25, 8.24108e-26, -2.197619e-25, -6.043449e-26, 
    1.538334e-25, -1.098805e-26, 9.339889e-26, -1.867976e-25, -1.263631e-25, 
    -1.098805e-26, 9.889295e-26, 1.181221e-25, -3.021727e-25, 6.04346e-26, 
    1.428453e-25, -3.845829e-26, -2.087738e-25, -6.592854e-26, 5.494055e-26, 
    1.318572e-25, 2.19762e-25, -4.944639e-26, -1.922912e-26, -4.669937e-26, 
    3.076668e-25, 1.346043e-25, 1.153751e-25, 1.263632e-25, 2.74703e-26, 
    -1.20869e-25, -1.291101e-25, -2.74702e-26, 1.64822e-26, 1.455924e-25, 
    -2.005328e-25, -1.648209e-26, -2.746971e-27, 1.04387e-25, 5.351395e-32, 
    -1.18122e-25, 8.24108e-26, 1.703156e-25, -5.219342e-26, -2.911846e-25, 
    4.395245e-26, -1.593274e-25, 3.84584e-26, 1.895448e-25, -1.648209e-26, 
    -6.592854e-26, -2.060268e-25, -4.669937e-26 ;

 M_LITR3C_TO_LEACHING =
  -2.609671e-26, -4.669939e-26, 2.060271e-26, -6.867535e-27, -1.208691e-25, 
    -1.002664e-25, -2.060266e-26, 1.510866e-26, 2.747052e-27, -4.120535e-26, 
    -7.279613e-26, -8.790477e-26, -8.241071e-26, -6.592857e-26, 2.087739e-25, 
    9.477238e-26, -5.356696e-26, -1.510863e-25, -2.747022e-26, 1.263632e-25, 
    -2.47232e-26, -7.416964e-26, -6.180803e-26, 1.648217e-26, -6.592857e-26, 
    4.532594e-26, 8.103726e-26, 9.889292e-26, -1.414718e-25, 4.944647e-26, 
    -5.494023e-27, -7.829018e-26, 7.554321e-26, 9.065185e-26, 7.416969e-26, 
    -6.730208e-26, 9.614614e-27, -1.071339e-25, 1.593275e-25, -5.494023e-27, 
    -8.653126e-26, 6.867565e-26, 1.098813e-26, 7.142267e-26, -7.142262e-26, 
    2.060271e-26, 1.373513e-25, -7.142262e-26, 4.395242e-26, -1.469658e-25, 
    -1.030134e-25, -1.194956e-25, -7.691667e-26, -1.634479e-25, 
    -2.060266e-26, 1.373515e-26, 1.373539e-27, -3.845832e-26, -1.648212e-26, 
    1.387248e-25, 2.884379e-26, -4.395237e-26, -1.12628e-25, 1.771831e-25, 
    7.142267e-26, 1.04387e-25, -4.807291e-26, -2.609671e-26, -1.895447e-25, 
    -3.159076e-26, -4.532588e-26, 2.747052e-27, 1.92292e-26, 3.571135e-26, 
    1.09881e-25, 1.648217e-26, 2.675693e-32, -7.691667e-26, -4.669939e-26, 
    5.631404e-26, 2.675704e-32, 1.346042e-25, -3.57113e-26, 4.944647e-26, 
    -5.494023e-27, 8.378428e-26, -3.296427e-26, -1.277366e-25, -7.691667e-26, 
    8.241101e-27, -2.747022e-26, -3.708481e-26, -1.373486e-27, 1.057605e-25, 
    -3.296427e-26, 4.944647e-26, 1.359778e-25, -3.296427e-26, 4.395242e-26, 
    8.241077e-26, 2.747052e-27, -5.494047e-26, -4.120535e-26, -5.356696e-26, 
    -7.691667e-26, 7.691672e-26, 7.142267e-26, -3.433778e-26, 2.334974e-26, 
    5.768755e-26, -4.669939e-26, -5.631398e-26, -1.922915e-26, -2.884373e-26, 
    -2.115209e-25, -8.378423e-26, -5.906101e-26, -6.867559e-26, -9.61456e-27, 
    1.112545e-25, 1.263632e-25, -9.889287e-26, -5.768749e-26, -1.263631e-25, 
    -1.09881e-25, 2.747052e-27, -5.494047e-26, 1.153751e-25, -5.494047e-26, 
    3.02173e-26, -2.746998e-27, 4.944647e-26, 1.085075e-25, -3.845832e-26, 
    5.494076e-27, -1.15375e-25, 4.257891e-26, -7.00491e-26, -1.552069e-25, 
    -6.180803e-26, -3.57113e-26, -2.170149e-25, -7.416964e-26, -2.074003e-25, 
    -1.346042e-25, 1.977858e-25, -4.807291e-26, -5.494023e-27, -6.592857e-26, 
    1.373539e-27, 2.334974e-26, -1.455923e-25, -3.57113e-26, 5.494076e-27, 
    -1.09881e-25, 6.455511e-26, -2.747022e-26, 1.373515e-26, -1.043869e-25, 
    9.477238e-26, -2.47232e-26, -3.57113e-26, -1.318572e-25, 8.241101e-27, 
    -3.296427e-26, -1.15375e-25, -8.927828e-26, 5.081998e-26, -6.043452e-26, 
    8.653131e-26, -1.236161e-25, 1.92292e-26, 4.944647e-26, 2.747052e-27, 
    7.966375e-26, 8.515779e-26, 3.02173e-26, -7.691667e-26, -6.592857e-26, 
    -5.219344e-26, 1.387248e-25, -5.631398e-26, 8.241077e-26, 2.197622e-26, 
    1.648217e-26, 8.241101e-27, 1.112545e-25, 3.708486e-26, 6.455511e-26, 
    -5.494047e-26, -5.768749e-26, -1.538334e-25, -1.194956e-25, 1.318572e-25, 
    7.691672e-26, 5.356701e-26, 1.016399e-25, 1.510866e-26, 8.241101e-27, 
    -6.592857e-26, 1.04387e-25, 4.944647e-26, -1.071339e-25, -1.112545e-25, 
    4.944647e-26, 1.785569e-26, 1.098813e-26, -3.708481e-26, -5.906101e-26, 
    -1.648212e-26, 1.194956e-25, -1.098807e-26, -7.142262e-26, -5.081993e-26, 
    2.060271e-26, 3.708486e-26, 3.433784e-26, 4.395242e-26, 1.346042e-25, 
    9.614589e-26, 3.708486e-26, -2.197617e-26, -2.334968e-26, -2.197617e-26, 
    6.043457e-26, -2.884373e-26, -1.085074e-25, -2.746998e-27, 5.494052e-26, 
    7.966375e-26, -8.927828e-26, -9.477233e-26, 2.197622e-26, 3.433784e-26, 
    1.098813e-26, -6.318154e-26, -5.494023e-27, -3.845832e-26, -1.016399e-25, 
    2.675693e-32, 6.867565e-26, -1.057604e-25, 9.614614e-27, -8.653126e-26, 
    -7.416964e-26, -6.867535e-27, 5.494076e-27, 2.197622e-26, 1.057605e-25, 
    -7.829018e-26, -6.592857e-26, -4.120535e-26, -5.356696e-26, 
    -2.197617e-26, -4.120535e-26, 2.472325e-26, -5.631398e-26, -1.895447e-25, 
    3.433784e-26, 1.153751e-25, 1.12628e-25, 1.92292e-26, 9.614614e-27, 
    -5.219344e-26, -9.614584e-26, -1.098807e-26, -1.12628e-25, 4.944647e-26, 
    -2.197617e-26, -1.236158e-26, -3.433778e-26, 1.346042e-25, -1.016399e-25, 
    -8.241047e-27, -3.296427e-26, 4.12054e-26, -2.197617e-26, -5.906101e-26, 
    -3.708481e-26, -4.944642e-26, -3.433778e-26, 2.675689e-32, -7.554316e-26, 
    -1.249896e-25, -1.12628e-25, 9.202536e-26, -1.813036e-25, 8.241101e-27, 
    5.494052e-26, -1.263631e-25, 9.065185e-26, -1.318572e-25, 3.296432e-26, 
    -1.428453e-25, 5.494076e-27, -5.219344e-26, -1.469658e-25, 3.296432e-26, 
    -1.37351e-26, 1.373515e-26, -5.906101e-26, 5.21935e-26, -5.219344e-26, 
    -9.065179e-26, 8.515779e-26, -2.47232e-26, -5.631398e-26, 2.675685e-32, 
    9.889292e-26, -1.922915e-26, -1.510861e-26, -1.977858e-25, -4.395237e-26, 
    -1.524598e-25, 5.21935e-26, 5.631404e-26, -1.002664e-25, 5.081998e-26, 
    -1.813036e-25, -3.57113e-26, -8.241047e-27, 1.263632e-25, -3.708481e-26, 
    -6.867559e-26, 6.043457e-26, 7.142267e-26, -5.219344e-26, -2.060266e-26, 
    2.609676e-26, -2.087739e-25, 1.648217e-26, -5.081993e-26, 9.065185e-26, 
    -1.222426e-25, 7.691672e-26, -2.719554e-25, -1.043869e-25, -8.790477e-26 ;

 M_SOIL1C_TO_LEACHING =
  5.610788e-21, 5.019039e-21, 1.348146e-20, -6.184819e-20, -2.989907e-20, 
    2.171035e-20, 8.483887e-21, 7.027556e-21, 4.748603e-20, -1.49392e-20, 
    -1.452642e-20, 1.540148e-20, -3.125759e-20, -8.829132e-21, 4.916692e-21, 
    -3.561248e-20, 1.523692e-20, 3.870132e-20, -1.50328e-20, -2.304961e-20, 
    -3.211085e-20, -3.822351e-22, -1.185857e-20, 9.967955e-21, 3.344677e-20, 
    -1.015146e-20, -1.643231e-20, -2.516135e-20, 1.910101e-20, 2.094497e-20, 
    1.189873e-20, 1.986552e-20, 1.949937e-20, -4.024961e-21, -1.941218e-21, 
    1.083537e-20, -1.696583e-20, -1.327421e-20, 1.732378e-20, 2.239804e-21, 
    1.348286e-20, 2.979415e-21, 4.430098e-21, -9.63801e-21, 2.639065e-20, 
    -4.865785e-21, 4.904446e-20, -3.050637e-20, -3.013515e-20, 4.407207e-21, 
    -1.23149e-20, -4.513063e-20, -1.587336e-20, -5.060334e-21, -6.926327e-21, 
    -1.6272e-20, 1.305623e-20, -1.151307e-20, -2.793351e-20, 7.88395e-21, 
    -5.709755e-21, 1.930513e-20, 5.897468e-21, 7.178375e-22, 6.918138e-21, 
    3.600151e-20, 3.212584e-20, -1.950077e-20, -7.969594e-21, 4.233132e-20, 
    -1.449559e-20, -4.661158e-20, -2.148953e-20, -2.527839e-20, 
    -1.071381e-20, -4.39758e-21, 1.777046e-20, -2.072981e-20, -6.670491e-21, 
    -2.736634e-20, 1.635899e-21, -2.143411e-20, -3.612366e-20, -1.222274e-20, 
    -7.925176e-22, -3.787175e-21, -3.122761e-20, -1.448627e-20, 1.211754e-20, 
    2.573101e-20, -4.308421e-20, 1.900657e-20, -6.512412e-21, -2.036511e-21, 
    1.549449e-20, 2.980575e-20, 1.108389e-20, 2.829003e-20, 2.297074e-20, 
    -2.826827e-20, 2.198796e-20, -1.974586e-21, 2.887829e-21, 1.499744e-20, 
    2.028001e-20, -1.77541e-20, -1.20087e-20, -6.180779e-21, 2.818402e-20, 
    -1.982309e-20, 2.33139e-21, 2.444717e-20, 3.585599e-21, 9.553762e-21, 
    3.03486e-20, 1.786518e-20, 9.222407e-21, 1.692342e-20, -8.315957e-21, 
    -1.240397e-20, -3.940975e-21, 4.690052e-20, -2.193087e-20, 1.651426e-21, 
    -1.954943e-20, -1.892626e-20, 1.554142e-20, -9.822916e-21, -4.731471e-20, 
    -2.418169e-20, -2.88227e-20, -5.823403e-21, 1.72446e-20, -5.172838e-21, 
    1.946318e-20, -1.61968e-20, -2.067666e-20, 3.778987e-21, 8.103652e-21, 
    -1.69938e-20, -2.088164e-20, 3.713078e-20, -6.254298e-21, 2.480455e-20, 
    2.307988e-20, 2.127183e-20, 2.243865e-20, 1.7354e-20, -9.081572e-21, 
    -2.704378e-20, 1.12934e-20, -6.535052e-21, -1.01475e-20, -4.617022e-20, 
    3.750113e-20, -9.188417e-22, -8.813007e-21, -6.012282e-21, -1.161176e-20, 
    -8.291643e-21, 4.870604e-21, 1.265136e-20, 3.295001e-20, -5.531903e-21, 
    1.310062e-20, 1.494487e-20, 6.599841e-20, 5.204517e-21, -6.038564e-21, 
    -7.877157e-21, 3.693171e-20, -1.912986e-20, -1.777528e-20, 1.835994e-20, 
    3.022341e-22, 3.702644e-21, 6.896103e-21, 1.633815e-20, -1.151393e-20, 
    -2.480969e-21, -3.06791e-21, -1.027983e-20, -3.354912e-20, 1.257501e-20, 
    2.609523e-20, 5.966298e-20, -8.578896e-21, -1.801898e-20, 8.252055e-21, 
    3.018687e-20, -2.882154e-21, -6.675855e-21, 4.758924e-21, -1.374553e-20, 
    4.817152e-21, -2.281637e-20, 3.251771e-20, -1.545662e-20, 2.436373e-20, 
    -1.440938e-20, 1.514731e-20, 2.235015e-20, -2.555461e-20, 4.55792e-21, 
    1.787563e-20, -7.239893e-21, 7.542127e-21, 2.583566e-20, 8.086167e-22, 
    3.123908e-21, -4.063889e-20, 5.025512e-20, 1.769725e-20, -4.95613e-20, 
    -5.092558e-21, 5.794575e-21, 1.847899e-20, -3.60629e-20, -1.299006e-20, 
    -3.450419e-20, -7.097107e-21, 1.625644e-20, 3.846524e-20, 2.694255e-20, 
    -1.363752e-20, 2.764908e-20, 9.636321e-21, 1.773287e-20, 7.266181e-21, 
    -1.418197e-21, -2.362613e-20, -1.789177e-20, -3.288668e-20, 1.138981e-20, 
    -4.189221e-20, 2.128228e-20, -6.476514e-21, 3.862038e-22, 2.324215e-22, 
    4.663304e-20, 5.439745e-21, 1.047379e-20, -3.106872e-20, 9.292792e-21, 
    -1.303613e-20, 7.798535e-21, -1.375034e-20, -4.052663e-20, -3.818478e-20, 
    -1.412918e-20, -5.960253e-21, -7.746555e-21, 7.143767e-21, 3.428404e-21, 
    -3.255933e-21, -8.316502e-21, 4.598671e-20, 7.910232e-21, -1.126061e-20, 
    2.749868e-20, 2.194585e-20, -2.069813e-20, 1.23166e-20, -6.378359e-22, 
    -1.532456e-20, -3.025814e-20, -2.012533e-20, -5.708048e-21, 
    -1.635397e-20, 3.820822e-21, -7.893282e-21, -8.335762e-21, -5.282288e-20, 
    -2.680713e-20, -2.136909e-20, 8.21107e-21, 2.201737e-20, -3.171947e-21, 
    1.442465e-20, -6.742009e-21, -2.011545e-20, 7.323308e-21, 2.665875e-21, 
    1.38244e-20, 5.279317e-20, -5.298544e-20, 2.131647e-20, 1.373505e-20, 
    -1.643119e-20, 5.130457e-21, 5.932543e-21, -2.003598e-20, -4.7442e-22, 
    2.134392e-20, -1.998457e-20, 9.228317e-21, 3.009528e-20, -3.46806e-20, 
    -1.737238e-20, -1.352781e-20, 1.1061e-20, -2.762302e-22, -1.955479e-20, 
    2.819702e-20, 2.279716e-20, 2.892053e-20, 1.084558e-20, 1.874672e-20, 
    -1.530956e-20, 8.324178e-21, -3.039187e-20, 8.433286e-21, -1.040533e-20, 
    1.991159e-20, 4.165469e-21, 3.063925e-20, -2.179742e-20, -1.660758e-21, 
    3.666198e-20, -4.862601e-20, -1.25066e-20, 1.771223e-20, -1.568109e-20, 
    8.757865e-21, 4.802171e-21, 1.494827e-20, 1.805745e-20, 1.115107e-21, 
    1.619934e-20, 3.506715e-21, -2.932739e-20, 8.060928e-21, 2.407253e-20, 
    1.898651e-20, -1.429231e-20, 3.310326e-20, -3.183842e-21, 5.509461e-20 ;

 M_SOIL2C_TO_LEACHING =
  -9.988594e-21, -2.797423e-20, -1.144219e-21, 8.032101e-21, -1.435792e-20, 
    4.694008e-20, -8.466081e-21, -2.075555e-20, 3.589352e-20, -2.209486e-20, 
    1.073445e-20, -2.137783e-20, -1.405285e-20, 3.006418e-20, -1.142218e-21, 
    6.796008e-21, 3.186928e-21, -1.146276e-20, 2.124608e-20, -7.811678e-22, 
    -4.755376e-22, -6.241285e-21, -4.562454e-20, -2.265435e-20, 
    -1.928395e-20, -8.077616e-21, 1.462143e-20, -4.247749e-21, -1.409125e-21, 
    5.336264e-21, 8.039172e-21, -8.695679e-21, -3.208825e-20, -2.844837e-20, 
    1.312238e-20, -3.565432e-20, -1.489935e-20, -6.032259e-20, -2.216638e-20, 
    -4.704131e-20, 1.0722e-20, 2.768501e-21, -9.744604e-21, -3.524237e-21, 
    -2.212508e-20, -1.293775e-20, 3.32938e-20, -8.515693e-22, -6.000404e-21, 
    4.043894e-21, 5.161253e-21, -2.431383e-23, -1.773966e-20, -1.422304e-20, 
    3.226074e-20, -1.836311e-20, 3.596906e-21, -1.579587e-20, 2.600558e-20, 
    2.73641e-20, -7.283702e-21, 2.245843e-20, -1.31744e-20, -4.743943e-21, 
    7.969888e-21, 1.049525e-20, 7.643046e-21, -9.906313e-21, 2.097153e-20, 
    -4.394477e-21, -1.180118e-20, 7.123111e-21, -1.144438e-20, -1.79192e-20, 
    2.897113e-20, -7.294742e-21, 3.715011e-22, 2.599849e-20, -6.129765e-22, 
    -2.510931e-21, 2.580852e-20, 2.372686e-21, 4.449326e-21, 2.289073e-20, 
    3.570464e-20, -1.277362e-21, 2.427725e-20, 3.055586e-20, 4.829047e-21, 
    -8.617581e-22, -3.243776e-21, -1.543313e-20, 6.075892e-21, 1.5686e-21, 
    1.55926e-20, 1.602829e-20, -2.607682e-20, 2.045981e-20, 1.826641e-20, 
    1.405086e-20, -1.036769e-21, 3.989925e-20, 3.388134e-20, -9.809053e-21, 
    3.167459e-20, -5.187819e-21, 2.93138e-20, 1.922598e-20, 3.618958e-21, 
    -2.753771e-20, 1.453518e-20, -1.785984e-20, -1.504135e-21, 1.078038e-21, 
    -1.798593e-20, -2.743705e-20, -5.148524e-21, -2.790893e-20, 5.773086e-21, 
    -3.361473e-20, 5.739155e-21, -1.075537e-20, 2.53652e-20, -1.473196e-20, 
    -1.074661e-20, 5.246357e-21, 4.62785e-20, 3.487736e-20, -2.180618e-20, 
    -1.490499e-20, 1.060351e-20, -6.474824e-21, 2.240982e-20, -2.920099e-20, 
    1.461917e-20, 1.490811e-20, 2.137868e-20, 1.717845e-20, 2.018726e-20, 
    2.263033e-20, -2.700417e-20, 1.167509e-20, 2.933034e-21, -1.366153e-20, 
    -2.325124e-20, -5.812979e-22, -2.685348e-20, 3.317621e-20, 3.348776e-20, 
    -4.871149e-21, -4.957485e-20, 1.452302e-20, -1.053905e-20, 4.207233e-20, 
    -3.842029e-20, -4.382864e-20, 1.669893e-20, 3.441769e-20, -2.717723e-20, 
    -3.347842e-20, 8.928907e-21, -2.383419e-20, 3.974082e-21, -8.395403e-21, 
    -1.752903e-20, -5.120619e-20, -1.300308e-20, 7.249085e-22, -2.315084e-20, 
    -1.652675e-20, 2.975473e-21, -3.688394e-20, 3.147584e-20, -1.09782e-21, 
    -1.494033e-20, 1.499744e-20, 2.272591e-21, -5.296103e-21, -1.912815e-20, 
    4.3497e-20, -2.169083e-20, 5.42531e-21, 2.990926e-20, 8.549496e-21, 
    -1.420865e-20, 1.219898e-20, 2.688261e-20, 7.033777e-21, -2.42306e-20, 
    -3.243204e-21, -1.642893e-20, -7.687737e-21, -8.951825e-21, 5.003486e-21, 
    -2.50084e-20, -2.927385e-21, -2.749868e-20, 3.008815e-21, -3.517728e-21, 
    -1.924068e-20, -1.180712e-20, -2.668866e-20, -1.144666e-20, 1.142219e-21, 
    -1.332782e-21, -2.138859e-20, 3.781354e-20, -3.593196e-20, -1.768055e-20, 
    6.770266e-21, 5.331681e-20, 8.936272e-21, 1.73413e-20, 1.866303e-21, 
    -1.376872e-20, -2.925896e-20, -1.790844e-20, 1.029311e-20, 3.096272e-20, 
    1.934049e-20, 8.81358e-21, 8.826281e-21, 2.449777e-20, 1.389508e-20, 
    1.205509e-20, 3.423007e-21, 3.324234e-20, 9.857965e-21, -3.036755e-20, 
    -4.931616e-20, -3.686838e-20, 1.628955e-20, 2.083895e-20, -1.485411e-20, 
    -2.774606e-20, -2.062889e-20, -1.407461e-20, -9.934879e-21, 3.638741e-21, 
    -2.440899e-20, 8.606606e-21, -2.64636e-20, 2.428655e-20, 1.414022e-20, 
    -3.244505e-20, -2.112451e-20, -3.201642e-20, -8.886804e-21, 2.57681e-20, 
    -2.176123e-20, -1.337516e-20, 1.158262e-20, 3.13014e-20, 1.869132e-20, 
    -1.709107e-20, -1.699608e-20, 2.782041e-20, -6.308868e-21, 4.308193e-20, 
    1.943095e-20, -2.479852e-21, 2.187882e-20, 7.751068e-21, 8.407575e-21, 
    -1.277122e-20, 3.808404e-21, 2.341266e-20, -1.877868e-20, -1.78898e-20, 
    2.198205e-20, -2.289695e-20, -2.279546e-20, 6.873185e-21, 2.085053e-20, 
    -5.227407e-21, 8.440078e-21, 3.989896e-21, 3.420082e-20, -6.486392e-21, 
    -1.805123e-20, -4.901138e-21, 2.863667e-20, -1.71824e-20, -8.677301e-21, 
    1.303362e-20, -1.564659e-20, -2.613278e-21, 1.758726e-20, -3.682625e-20, 
    -1.454734e-20, 1.994807e-20, 9.945037e-21, 1.736335e-20, 4.455272e-20, 
    1.798026e-20, 9.391759e-21, -1.310747e-21, -5.280549e-21, -5.885636e-20, 
    -2.295237e-20, 2.763213e-20, -1.857542e-21, 2.545566e-20, -1.000585e-20, 
    -3.514851e-20, -9.054451e-21, -1.560248e-20, -1.659147e-20, 2.73299e-20, 
    -3.412958e-20, 1.27845e-20, 2.007615e-20, -2.893382e-20, -1.564207e-20, 
    1.532145e-20, 1.844311e-20, -4.024644e-20, -4.672685e-21, 1.423859e-20, 
    9.53056e-21, 4.738268e-21, 5.153889e-21, 5.909079e-21, -8.941947e-21, 
    -1.898368e-20, -1.262479e-20, 1.221058e-20, -6.49717e-21, -4.832443e-21, 
    -2.151327e-20, 3.373685e-20, -2.093849e-20, -5.090558e-21, -7.889314e-21, 
    1.393662e-20, 9.648478e-21, 6.723606e-21, -1.544586e-20 ;

 M_SOIL3C_TO_LEACHING =
  1.231772e-20, -3.586995e-21, -2.724365e-20, 2.924845e-21, 4.012504e-21, 
    4.861445e-20, 5.754708e-21, 7.887608e-21, 4.869698e-20, -1.285887e-20, 
    -1.007906e-20, 4.923484e-21, -6.952069e-21, 2.476325e-20, 4.351961e-20, 
    3.386548e-20, -1.647303e-20, 3.229437e-20, -2.849415e-20, 6.8616e-21, 
    -1.45089e-20, -1.289451e-20, 2.745232e-20, -4.730358e-21, -2.757388e-20, 
    1.147743e-20, 8.104737e-21, 5.544649e-21, 2.365496e-20, -7.628921e-21, 
    -1.96784e-22, -1.767916e-20, 5.34093e-22, -2.18418e-20, 1.990877e-20, 
    -1.447582e-20, -1.510927e-21, -3.263589e-20, 3.956528e-21, 1.346448e-20, 
    -3.967289e-21, 8.244315e-22, 7.270428e-21, 3.049228e-21, 4.541506e-20, 
    -1.015429e-20, -3.293924e-20, 1.85904e-20, -4.652902e-21, -1.359342e-20, 
    -3.063417e-20, -3.533373e-20, 1.576225e-20, 3.436677e-20, -4.364772e-20, 
    9.261113e-21, -1.553379e-20, -6.732938e-21, 2.342168e-21, -1.872696e-20, 
    1.335917e-21, -1.549138e-20, 6.660302e-21, -8.553464e-21, 5.093954e-21, 
    -2.715659e-20, 6.049677e-20, -1.546253e-20, 3.150158e-20, 1.668734e-20, 
    -1.918048e-21, -1.273052e-20, -6.570378e-21, 1.988785e-20, -2.845147e-20, 
    -8.344506e-21, 5.492665e-20, -2.282739e-20, -9.362342e-21, -4.198777e-20, 
    -3.871234e-20, 1.038978e-20, 5.824831e-21, -1.218175e-20, 1.25086e-20, 
    -1.607494e-20, -1.780185e-20, -4.736955e-20, 1.033099e-20, -3.288157e-21, 
    -2.585969e-20, -5.12675e-21, 2.261027e-20, 3.937889e-21, 7.237069e-21, 
    1.393864e-20, -1.662146e-20, 2.660752e-20, -2.053307e-20, 4.648934e-21, 
    -1.160018e-20, 4.527566e-20, 2.523088e-21, -5.102715e-21, -3.939316e-20, 
    -3.153409e-20, -1.969983e-20, 5.669318e-20, 5.068523e-21, -3.774473e-21, 
    -3.530797e-20, -6.930294e-21, -1.536359e-21, 2.210984e-20, 5.404697e-21, 
    -2.3921e-20, -5.598058e-21, -1.603056e-20, -1.773569e-20, -1.715667e-20, 
    -2.907772e-20, 2.249972e-20, 9.90971e-21, -5.951445e-22, 2.061276e-20, 
    2.331963e-21, -3.474708e-22, 1.219304e-20, 3.932671e-20, -1.185829e-20, 
    3.445074e-20, 1.74538e-20, 1.706903e-20, 2.972623e-21, -6.840682e-21, 
    -3.447591e-20, 1.707243e-20, 8.471757e-21, -7.78272e-21, 7.148853e-21, 
    3.483073e-20, 2.455998e-20, -8.902341e-21, 3.339332e-20, 2.868024e-21, 
    2.947191e-21, 4.153884e-21, 5.010278e-21, 1.987427e-20, 3.700437e-20, 
    6.404129e-21, 2.213074e-20, -2.069053e-20, -2.746078e-20, 4.949488e-21, 
    -8.989414e-21, 2.703415e-20, 3.417168e-20, -2.837767e-20, 5.229244e-20, 
    -4.266521e-20, -1.935854e-21, -9.843293e-21, -4.007651e-20, 
    -3.228303e-20, -3.406144e-20, -2.059119e-21, 4.982846e-21, -4.892146e-20, 
    5.021007e-21, -3.59905e-20, 6.021616e-21, -1.494033e-20, 3.761155e-21, 
    2.047197e-20, 4.042204e-21, -1.925119e-21, -7.847757e-21, 3.655085e-20, 
    -2.110359e-20, -3.380415e-20, 5.127633e-21, -1.634664e-20, -4.300421e-20, 
    -4.632062e-20, -7.722502e-21, -3.837231e-21, 1.714336e-20, 2.94266e-20, 
    1.403818e-20, 2.836723e-20, -1.031035e-20, 1.104262e-20, -1.178169e-20, 
    1.057186e-20, -2.388197e-20, 7.480487e-21, 3.377776e-21, -1.146187e-21, 
    -8.945033e-21, 2.141425e-21, 1.359511e-20, -2.100378e-20, -4.188288e-20, 
    -1.815131e-20, -5.302388e-20, 6.548033e-21, -2.079456e-20, -1.438421e-20, 
    3.387109e-21, -1.049355e-20, -3.086458e-20, -4.400987e-20, -1.002592e-20, 
    2.353535e-20, 8.491251e-21, 9.221835e-21, -1.613147e-20, 2.823434e-20, 
    -4.838925e-21, -1.03652e-20, 1.164031e-20, 1.1454e-20, 4.333133e-20, 
    2.971784e-20, -1.307291e-20, -3.692193e-21, 8.334335e-21, -2.252233e-20, 
    3.601142e-20, -8.855126e-21, -5.298927e-21, -1.55875e-20, 2.835773e-21, 
    3.492347e-20, 2.872883e-20, -1.977149e-21, 1.249104e-20, -4.171128e-20, 
    -3.048682e-21, -1.622791e-20, -2.929118e-20, -1.692624e-20, 
    -2.054943e-20, -7.636409e-22, -9.312597e-21, -5.886162e-21, 
    -3.107609e-20, 1.174719e-20, 3.82562e-21, -1.903202e-20, -2.258678e-20, 
    2.571438e-21, -8.71489e-21, 6.740303e-21, 3.597756e-21, 2.02421e-20, 
    1.402173e-20, -7.513845e-21, -2.700079e-20, 8.722228e-21, -4.267791e-20, 
    2.998644e-20, -1.459182e-21, 3.103593e-20, 8.784441e-21, 5.086268e-20, 
    -1.443425e-20, -6.747096e-21, -2.98886e-20, 2.551616e-20, 7.53421e-20, 
    2.534343e-20, 1.379923e-20, 6.440894e-21, -1.660109e-20, 9.9018e-21, 
    4.97083e-20, 6.233921e-21, 2.623687e-20, -4.912446e-20, 3.89781e-20, 
    -1.260612e-20, -1.86803e-20, 2.505787e-20, 4.135615e-20, -1.150374e-20, 
    3.638831e-20, 8.149429e-21, 2.878212e-21, -1.281731e-20, -8.086098e-21, 
    9.179143e-21, 4.404945e-21, -7.490381e-21, 1.638624e-20, 2.126756e-20, 
    -2.908112e-20, 1.653494e-20, 1.235391e-20, -2.254467e-20, -3.863235e-21, 
    -6.829065e-21, -7.327822e-21, 2.82476e-21, 2.457043e-20, -3.801967e-20, 
    -1.242235e-20, -9.774877e-21, 2.474715e-20, -3.132562e-22, 1.098551e-20, 
    -5.7615e-21, -2.895161e-20, 1.028461e-20, -4.473361e-21, -2.685548e-20, 
    -1.344696e-20, 3.337947e-20, -9.365739e-21, 7.166069e-21, -9.330118e-21, 
    -9.707839e-21, 2.087062e-20, 2.752097e-21, -1.366409e-20, 2.023786e-20, 
    2.536547e-20, 1.976544e-20, 1.550553e-20, -1.397961e-20, -1.001913e-20, 
    1.200108e-20, -3.952046e-21, 7.697927e-21, -1.632289e-20, -3.442103e-20, 
    8.801657e-21 ;

 NBP =
  -7.624269e-08, -7.645139e-08, -7.641083e-08, -7.657911e-08, -7.648578e-08, 
    -7.659595e-08, -7.628502e-08, -7.645966e-08, -7.634819e-08, -7.62615e-08, 
    -7.690554e-08, -7.658662e-08, -7.723681e-08, -7.70335e-08, -7.754418e-08, 
    -7.720516e-08, -7.761253e-08, -7.753444e-08, -7.776953e-08, -7.77022e-08, 
    -7.800275e-08, -7.780061e-08, -7.815856e-08, -7.79545e-08, -7.798641e-08, 
    -7.779394e-08, -7.665084e-08, -7.686582e-08, -7.663809e-08, 
    -7.666875e-08, -7.6655e-08, -7.648769e-08, -7.640334e-08, -7.622676e-08, 
    -7.625883e-08, -7.638853e-08, -7.668255e-08, -7.658277e-08, 
    -7.683426e-08, -7.682858e-08, -7.710845e-08, -7.698227e-08, 
    -7.745253e-08, -7.731892e-08, -7.7705e-08, -7.760792e-08, -7.770044e-08, 
    -7.767239e-08, -7.77008e-08, -7.755842e-08, -7.761943e-08, -7.749413e-08, 
    -7.700589e-08, -7.71494e-08, -7.67213e-08, -7.646373e-08, -7.629267e-08, 
    -7.617125e-08, -7.618841e-08, -7.622113e-08, -7.638929e-08, 
    -7.654739e-08, -7.666784e-08, -7.674839e-08, -7.682777e-08, 
    -7.706788e-08, -7.719501e-08, -7.747953e-08, -7.742823e-08, 
    -7.751517e-08, -7.759827e-08, -7.773771e-08, -7.771477e-08, 
    -7.777619e-08, -7.75129e-08, -7.768788e-08, -7.739899e-08, -7.747801e-08, 
    -7.684923e-08, -7.66097e-08, -7.650777e-08, -7.641862e-08, -7.620162e-08, 
    -7.635147e-08, -7.629239e-08, -7.643295e-08, -7.652225e-08, 
    -7.647809e-08, -7.67506e-08, -7.664466e-08, -7.720254e-08, -7.696229e-08, 
    -7.758857e-08, -7.743876e-08, -7.762448e-08, -7.752973e-08, 
    -7.769207e-08, -7.754596e-08, -7.779906e-08, -7.785415e-08, -7.78165e-08, 
    -7.796114e-08, -7.753786e-08, -7.770043e-08, -7.647685e-08, 
    -7.648405e-08, -7.651761e-08, -7.637008e-08, -7.636106e-08, 
    -7.622587e-08, -7.634618e-08, -7.639739e-08, -7.652743e-08, 
    -7.660432e-08, -7.667741e-08, -7.683809e-08, -7.701749e-08, -7.72683e-08, 
    -7.744847e-08, -7.75692e-08, -7.749518e-08, -7.756054e-08, -7.748747e-08, 
    -7.745323e-08, -7.78335e-08, -7.761999e-08, -7.794034e-08, -7.792262e-08, 
    -7.777765e-08, -7.792462e-08, -7.648911e-08, -7.644767e-08, 
    -7.630373e-08, -7.641638e-08, -7.621115e-08, -7.632602e-08, 
    -7.639206e-08, -7.664685e-08, -7.670285e-08, -7.675474e-08, 
    -7.685723e-08, -7.698873e-08, -7.721936e-08, -7.741998e-08, -7.76031e-08, 
    -7.758969e-08, -7.759441e-08, -7.76353e-08, -7.7534e-08, -7.765193e-08, 
    -7.767171e-08, -7.761997e-08, -7.792025e-08, -7.783448e-08, 
    -7.792224e-08, -7.78664e-08, -7.646114e-08, -7.653087e-08, -7.649319e-08, 
    -7.656404e-08, -7.651412e-08, -7.673605e-08, -7.680259e-08, 
    -7.711383e-08, -7.698614e-08, -7.718939e-08, -7.70068e-08, -7.703915e-08, 
    -7.719597e-08, -7.701667e-08, -7.74089e-08, -7.714296e-08, -7.763688e-08, 
    -7.737135e-08, -7.765352e-08, -7.760231e-08, -7.768711e-08, 
    -7.776304e-08, -7.785858e-08, -7.803479e-08, -7.7994e-08, -7.814135e-08, 
    -7.663483e-08, -7.672524e-08, -7.671731e-08, -7.681193e-08, -7.68819e-08, 
    -7.703356e-08, -7.727672e-08, -7.71853e-08, -7.735314e-08, -7.738683e-08, 
    -7.713184e-08, -7.728839e-08, -7.678577e-08, -7.686698e-08, 
    -7.681864e-08, -7.664195e-08, -7.720634e-08, -7.691673e-08, 
    -7.745144e-08, -7.729462e-08, -7.775221e-08, -7.752466e-08, 
    -7.797154e-08, -7.816244e-08, -7.834216e-08, -7.855203e-08, 
    -7.677461e-08, -7.671318e-08, -7.682319e-08, -7.697533e-08, 
    -7.711654e-08, -7.730418e-08, -7.732339e-08, -7.735854e-08, 
    -7.744958e-08, -7.752611e-08, -7.736963e-08, -7.754529e-08, 
    -7.688577e-08, -7.723148e-08, -7.668994e-08, -7.685301e-08, 
    -7.696638e-08, -7.691667e-08, -7.717485e-08, -7.723568e-08, 
    -7.748282e-08, -7.735509e-08, -7.811531e-08, -7.777906e-08, 
    -7.871185e-08, -7.845127e-08, -7.669171e-08, -7.677441e-08, 
    -7.706215e-08, -7.692525e-08, -7.731672e-08, -7.741303e-08, 
    -7.749135e-08, -7.75914e-08, -7.760222e-08, -7.76615e-08, -7.756436e-08, 
    -7.765767e-08, -7.730458e-08, -7.74624e-08, -7.702928e-08, -7.713471e-08, 
    -7.708622e-08, -7.703301e-08, -7.719722e-08, -7.737208e-08, 
    -7.737585e-08, -7.743191e-08, -7.758979e-08, -7.731831e-08, 
    -7.815863e-08, -7.763973e-08, -7.686458e-08, -7.702379e-08, 
    -7.704657e-08, -7.698489e-08, -7.740338e-08, -7.725177e-08, 
    -7.766006e-08, -7.754974e-08, -7.77305e-08, -7.764068e-08, -7.762746e-08, 
    -7.75121e-08, -7.744025e-08, -7.725872e-08, -7.711099e-08, -7.699384e-08, 
    -7.702109e-08, -7.714976e-08, -7.738279e-08, -7.760318e-08, 
    -7.755491e-08, -7.771676e-08, -7.728835e-08, -7.7468e-08, -7.739856e-08, 
    -7.757962e-08, -7.718286e-08, -7.752063e-08, -7.709649e-08, 
    -7.713369e-08, -7.724876e-08, -7.748016e-08, -7.75314e-08, -7.758604e-08, 
    -7.755232e-08, -7.738871e-08, -7.736191e-08, -7.724597e-08, 
    -7.721394e-08, -7.71256e-08, -7.705243e-08, -7.711927e-08, -7.718945e-08, 
    -7.738879e-08, -7.756837e-08, -7.776411e-08, -7.781203e-08, 
    -7.804059e-08, -7.785449e-08, -7.816151e-08, -7.790043e-08, 
    -7.835236e-08, -7.754026e-08, -7.789281e-08, -7.725401e-08, 
    -7.732286e-08, -7.744735e-08, -7.773286e-08, -7.757877e-08, 
    -7.775899e-08, -7.736087e-08, -7.715419e-08, -7.710074e-08, 
    -7.700096e-08, -7.710302e-08, -7.709473e-08, -7.719238e-08, -7.7161e-08, 
    -7.739541e-08, -7.72695e-08, -7.762712e-08, -7.775758e-08, -7.812591e-08, 
    -7.835159e-08, -7.858132e-08, -7.86827e-08, -7.871355e-08, -7.872645e-08 ;

 NDEPLOY =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NDEP_TO_SMINN =
  3.989144e-10, 3.989147e-10, 3.989121e-10, 3.989123e-10, 3.989108e-10, 
    3.989089e-10, 3.989084e-10, 3.989066e-10, 3.98906e-10, 3.989042e-10, 
    3.989026e-10, 3.989029e-10, 3.989014e-10, 3.988995e-10, 3.988979e-10, 
    3.988982e-10, 3.988966e-10, 3.988948e-10, 3.988943e-10, 3.988924e-10, 
    3.988909e-10, 3.988911e-10, 3.988885e-10, 3.988888e-10, 3.988872e-10, 
    3.988854e-10, 3.989112e-10, 3.989115e-10, 3.989089e-10, 3.989092e-10, 
    3.989076e-10, 3.989057e-10, 3.989052e-10, 3.989034e-10, 3.989018e-10, 
    3.989021e-10, 3.989005e-10, 3.988987e-10, 3.988971e-10, 3.988974e-10, 
    3.988947e-10, 3.98895e-10, 3.988934e-10, 3.988916e-10, 3.988911e-10, 
    3.988892e-10, 3.988887e-10, 3.988869e-10, 3.988853e-10, 3.988856e-10, 
    3.98883e-10, 3.988832e-10, 3.989091e-10, 3.989072e-10, 3.989067e-10, 
    3.989049e-10, 3.989033e-10, 3.989036e-10, 3.98901e-10, 3.989012e-10, 
    3.988997e-10, 3.988978e-10, 3.988973e-10, 3.988955e-10, 3.988939e-10, 
    3.988942e-10, 3.988926e-10, 3.988908e-10, 3.988903e-10, 3.988884e-10, 
    3.988879e-10, 3.98886e-10, 3.988855e-10, 3.988837e-10, 3.988821e-10, 
    3.988824e-10, 3.988798e-10, 3.9888e-10, 3.989059e-10, 3.98904e-10, 
    3.989035e-10, 3.989017e-10, 3.989001e-10, 3.989004e-10, 3.988988e-10, 
    3.98897e-10, 3.988965e-10, 3.988946e-10, 3.988941e-10, 3.988923e-10, 
    3.988907e-10, 3.98891e-10, 3.988894e-10, 3.988876e-10, 3.98886e-10, 
    3.988863e-10, 3.988836e-10, 3.988839e-10, 3.988813e-10, 3.988816e-10, 
    3.988789e-10, 3.988792e-10, 3.988766e-10, 3.988768e-10, 3.989017e-10, 
    3.989019e-10, 3.989004e-10, 3.988985e-10, 3.98898e-10, 3.988962e-10, 
    3.988946e-10, 3.988949e-10, 3.988933e-10, 3.988914e-10, 3.988899e-10, 
    3.988901e-10, 3.988886e-10, 3.988867e-10, 3.988862e-10, 3.988844e-10, 
    3.988839e-10, 3.98882e-10, 3.988815e-10, 3.988797e-10, 3.988781e-10, 
    3.988784e-10, 3.988757e-10, 3.98876e-10, 3.988744e-10, 3.988726e-10, 
    3.988995e-10, 3.988977e-10, 3.988972e-10, 3.988953e-10, 3.988938e-10, 
    3.98894e-10, 3.988924e-10, 3.988906e-10, 3.98889e-10, 3.988893e-10, 
    3.988878e-10, 3.988859e-10, 3.988854e-10, 3.988835e-10, 3.98883e-10, 
    3.988812e-10, 3.988807e-10, 3.988788e-10, 3.988783e-10, 3.988765e-10, 
    3.988749e-10, 3.988752e-10, 3.988725e-10, 3.988728e-10, 3.988712e-10, 
    3.988694e-10, 3.988963e-10, 3.988945e-10, 3.988929e-10, 3.988932e-10, 
    3.988906e-10, 3.988908e-10, 3.988893e-10, 3.988874e-10, 3.988858e-10, 
    3.988861e-10, 3.988835e-10, 3.988838e-10, 3.988822e-10, 3.988803e-10, 
    3.988798e-10, 3.98878e-10, 3.988775e-10, 3.988756e-10, 3.988751e-10, 
    3.988733e-10, 3.988717e-10, 3.98872e-10, 3.988694e-10, 3.988696e-10, 
    3.98867e-10, 3.988673e-10, 3.988931e-10, 3.988913e-10, 3.988908e-10, 
    3.988889e-10, 3.988874e-10, 3.988876e-10, 3.988861e-10, 3.988842e-10, 
    3.988826e-10, 3.988829e-10, 3.988803e-10, 3.988806e-10, 3.98879e-10, 
    3.988772e-10, 3.988767e-10, 3.988748e-10, 3.988743e-10, 3.988724e-10, 
    3.988719e-10, 3.988701e-10, 3.988685e-10, 3.988688e-10, 3.988662e-10, 
    3.988664e-10, 3.988649e-10, 3.98863e-10, 3.988899e-10, 3.988881e-10, 
    3.988865e-10, 3.988868e-10, 3.988842e-10, 3.988845e-10, 3.988829e-10, 
    3.98881e-10, 3.988795e-10, 3.988797e-10, 3.988782e-10, 3.988763e-10, 
    3.988758e-10, 3.98874e-10, 3.988724e-10, 3.988727e-10, 3.9887e-10, 
    3.988703e-10, 3.988687e-10, 3.988669e-10, 3.988653e-10, 3.988656e-10, 
    3.98863e-10, 3.988632e-10, 3.988606e-10, 3.988609e-10, 3.988868e-10, 
    3.988849e-10, 3.988833e-10, 3.988836e-10, 3.98881e-10, 3.988813e-10, 
    3.988786e-10, 3.988789e-10, 3.988763e-10, 3.988765e-10, 3.988739e-10, 
    3.988742e-10, 3.988716e-10, 3.988719e-10, 3.988703e-10, 3.988684e-10, 
    3.988679e-10, 3.988661e-10, 3.988645e-10, 3.988648e-10, 3.988632e-10, 
    3.988614e-10, 3.988609e-10, 3.98859e-10, 3.988585e-10, 3.988566e-10, 
    3.988836e-10, 3.988817e-10, 3.988802e-10, 3.988804e-10, 3.988778e-10, 
    3.988781e-10, 3.988765e-10, 3.988747e-10, 3.988731e-10, 3.988734e-10, 
    3.988707e-10, 3.98871e-10, 3.988684e-10, 3.988687e-10, 3.98866e-10, 
    3.988663e-10, 3.988637e-10, 3.988639e-10, 3.988613e-10, 3.988616e-10, 
    3.9886e-10, 3.988582e-10, 3.988566e-10, 3.988569e-10, 3.988542e-10, 
    3.988545e-10, 3.988793e-10, 3.988796e-10, 3.98878e-10, 3.988762e-10, 
    3.988746e-10, 3.988749e-10, 3.988722e-10, 3.988725e-10, 3.988699e-10, 
    3.988702e-10, 3.988686e-10, 3.988667e-10, 3.988652e-10, 3.988655e-10, 
    3.988628e-10, 3.988631e-10, 3.988605e-10, 3.988607e-10, 3.988592e-10, 
    3.988573e-10, 3.988568e-10, 3.98855e-10, 3.988545e-10, 3.988526e-10, 
    3.988521e-10, 3.988503e-10, 3.988761e-10, 3.988764e-10, 3.988748e-10, 
    3.98873e-10, 3.988725e-10, 3.988706e-10, 3.98869e-10, 3.988693e-10, 
    3.988678e-10, 3.988659e-10, 3.988644e-10, 3.988646e-10, 3.98862e-10, 
    3.988623e-10, 3.988607e-10, 3.988589e-10, 3.988573e-10, 3.988576e-10, 
    3.988549e-10, 3.988552e-10, 3.988536e-10, 3.988518e-10, 3.988513e-10, 
    3.988494e-10, 3.988489e-10, 3.988476e-10 ;

 NEE =
  7.624269e-08, 7.645139e-08, 7.641083e-08, 7.657911e-08, 7.648578e-08, 
    7.659595e-08, 7.628502e-08, 7.645966e-08, 7.634819e-08, 7.62615e-08, 
    7.690554e-08, 7.658662e-08, 7.723681e-08, 7.70335e-08, 7.754418e-08, 
    7.720516e-08, 7.761253e-08, 7.753444e-08, 7.776953e-08, 7.77022e-08, 
    7.800275e-08, 7.780061e-08, 7.815856e-08, 7.79545e-08, 7.798641e-08, 
    7.779394e-08, 7.665084e-08, 7.686582e-08, 7.663809e-08, 7.666875e-08, 
    7.6655e-08, 7.648769e-08, 7.640334e-08, 7.622676e-08, 7.625883e-08, 
    7.638853e-08, 7.668255e-08, 7.658277e-08, 7.683426e-08, 7.682858e-08, 
    7.710845e-08, 7.698227e-08, 7.745253e-08, 7.731892e-08, 7.7705e-08, 
    7.760792e-08, 7.770044e-08, 7.767239e-08, 7.77008e-08, 7.755842e-08, 
    7.761943e-08, 7.749413e-08, 7.700589e-08, 7.71494e-08, 7.67213e-08, 
    7.646373e-08, 7.629267e-08, 7.617125e-08, 7.618841e-08, 7.622113e-08, 
    7.638929e-08, 7.654739e-08, 7.666784e-08, 7.674839e-08, 7.682777e-08, 
    7.706788e-08, 7.719501e-08, 7.747953e-08, 7.742823e-08, 7.751517e-08, 
    7.759827e-08, 7.773771e-08, 7.771477e-08, 7.777619e-08, 7.75129e-08, 
    7.768788e-08, 7.739899e-08, 7.747801e-08, 7.684923e-08, 7.66097e-08, 
    7.650777e-08, 7.641862e-08, 7.620162e-08, 7.635147e-08, 7.629239e-08, 
    7.643295e-08, 7.652225e-08, 7.647809e-08, 7.67506e-08, 7.664466e-08, 
    7.720254e-08, 7.696229e-08, 7.758857e-08, 7.743876e-08, 7.762448e-08, 
    7.752973e-08, 7.769207e-08, 7.754596e-08, 7.779906e-08, 7.785415e-08, 
    7.78165e-08, 7.796114e-08, 7.753786e-08, 7.770043e-08, 7.647685e-08, 
    7.648405e-08, 7.651761e-08, 7.637008e-08, 7.636106e-08, 7.622587e-08, 
    7.634618e-08, 7.639739e-08, 7.652743e-08, 7.660432e-08, 7.667741e-08, 
    7.683809e-08, 7.701749e-08, 7.72683e-08, 7.744847e-08, 7.75692e-08, 
    7.749518e-08, 7.756054e-08, 7.748747e-08, 7.745323e-08, 7.78335e-08, 
    7.761999e-08, 7.794034e-08, 7.792262e-08, 7.777765e-08, 7.792462e-08, 
    7.648911e-08, 7.644767e-08, 7.630373e-08, 7.641638e-08, 7.621115e-08, 
    7.632602e-08, 7.639206e-08, 7.664685e-08, 7.670285e-08, 7.675474e-08, 
    7.685723e-08, 7.698873e-08, 7.721936e-08, 7.741998e-08, 7.76031e-08, 
    7.758969e-08, 7.759441e-08, 7.76353e-08, 7.7534e-08, 7.765193e-08, 
    7.767171e-08, 7.761997e-08, 7.792025e-08, 7.783448e-08, 7.792224e-08, 
    7.78664e-08, 7.646114e-08, 7.653087e-08, 7.649319e-08, 7.656404e-08, 
    7.651412e-08, 7.673605e-08, 7.680259e-08, 7.711383e-08, 7.698614e-08, 
    7.718939e-08, 7.70068e-08, 7.703915e-08, 7.719597e-08, 7.701667e-08, 
    7.74089e-08, 7.714296e-08, 7.763688e-08, 7.737135e-08, 7.765352e-08, 
    7.760231e-08, 7.768711e-08, 7.776304e-08, 7.785858e-08, 7.803479e-08, 
    7.7994e-08, 7.814135e-08, 7.663483e-08, 7.672524e-08, 7.671731e-08, 
    7.681193e-08, 7.68819e-08, 7.703356e-08, 7.727672e-08, 7.71853e-08, 
    7.735314e-08, 7.738683e-08, 7.713184e-08, 7.728839e-08, 7.678577e-08, 
    7.686698e-08, 7.681864e-08, 7.664195e-08, 7.720634e-08, 7.691673e-08, 
    7.745144e-08, 7.729462e-08, 7.775221e-08, 7.752466e-08, 7.797154e-08, 
    7.816244e-08, 7.834216e-08, 7.855203e-08, 7.677461e-08, 7.671318e-08, 
    7.682319e-08, 7.697533e-08, 7.711654e-08, 7.730418e-08, 7.732339e-08, 
    7.735854e-08, 7.744958e-08, 7.752611e-08, 7.736963e-08, 7.754529e-08, 
    7.688577e-08, 7.723148e-08, 7.668994e-08, 7.685301e-08, 7.696638e-08, 
    7.691667e-08, 7.717485e-08, 7.723568e-08, 7.748282e-08, 7.735509e-08, 
    7.811531e-08, 7.777906e-08, 7.871185e-08, 7.845127e-08, 7.669171e-08, 
    7.677441e-08, 7.706215e-08, 7.692525e-08, 7.731672e-08, 7.741303e-08, 
    7.749135e-08, 7.75914e-08, 7.760222e-08, 7.76615e-08, 7.756436e-08, 
    7.765767e-08, 7.730458e-08, 7.74624e-08, 7.702928e-08, 7.713471e-08, 
    7.708622e-08, 7.703301e-08, 7.719722e-08, 7.737208e-08, 7.737585e-08, 
    7.743191e-08, 7.758979e-08, 7.731831e-08, 7.815863e-08, 7.763973e-08, 
    7.686458e-08, 7.702379e-08, 7.704657e-08, 7.698489e-08, 7.740338e-08, 
    7.725177e-08, 7.766006e-08, 7.754974e-08, 7.77305e-08, 7.764068e-08, 
    7.762746e-08, 7.75121e-08, 7.744025e-08, 7.725872e-08, 7.711099e-08, 
    7.699384e-08, 7.702109e-08, 7.714976e-08, 7.738279e-08, 7.760318e-08, 
    7.755491e-08, 7.771676e-08, 7.728835e-08, 7.7468e-08, 7.739856e-08, 
    7.757962e-08, 7.718286e-08, 7.752063e-08, 7.709649e-08, 7.713369e-08, 
    7.724876e-08, 7.748016e-08, 7.75314e-08, 7.758604e-08, 7.755232e-08, 
    7.738871e-08, 7.736191e-08, 7.724597e-08, 7.721394e-08, 7.71256e-08, 
    7.705243e-08, 7.711927e-08, 7.718945e-08, 7.738879e-08, 7.756837e-08, 
    7.776411e-08, 7.781203e-08, 7.804059e-08, 7.785449e-08, 7.816151e-08, 
    7.790043e-08, 7.835236e-08, 7.754026e-08, 7.789281e-08, 7.725401e-08, 
    7.732286e-08, 7.744735e-08, 7.773286e-08, 7.757877e-08, 7.775899e-08, 
    7.736087e-08, 7.715419e-08, 7.710074e-08, 7.700096e-08, 7.710302e-08, 
    7.709473e-08, 7.719238e-08, 7.7161e-08, 7.739541e-08, 7.72695e-08, 
    7.762712e-08, 7.775758e-08, 7.812591e-08, 7.835159e-08, 7.858132e-08, 
    7.86827e-08, 7.871355e-08, 7.872645e-08 ;

 NEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NEP =
  -7.624269e-08, -7.645139e-08, -7.641083e-08, -7.657911e-08, -7.648578e-08, 
    -7.659595e-08, -7.628502e-08, -7.645966e-08, -7.634819e-08, -7.62615e-08, 
    -7.690554e-08, -7.658662e-08, -7.723681e-08, -7.70335e-08, -7.754418e-08, 
    -7.720516e-08, -7.761253e-08, -7.753444e-08, -7.776953e-08, -7.77022e-08, 
    -7.800275e-08, -7.780061e-08, -7.815856e-08, -7.79545e-08, -7.798641e-08, 
    -7.779394e-08, -7.665084e-08, -7.686582e-08, -7.663809e-08, 
    -7.666875e-08, -7.6655e-08, -7.648769e-08, -7.640334e-08, -7.622676e-08, 
    -7.625883e-08, -7.638853e-08, -7.668255e-08, -7.658277e-08, 
    -7.683426e-08, -7.682858e-08, -7.710845e-08, -7.698227e-08, 
    -7.745253e-08, -7.731892e-08, -7.7705e-08, -7.760792e-08, -7.770044e-08, 
    -7.767239e-08, -7.77008e-08, -7.755842e-08, -7.761943e-08, -7.749413e-08, 
    -7.700589e-08, -7.71494e-08, -7.67213e-08, -7.646373e-08, -7.629267e-08, 
    -7.617125e-08, -7.618841e-08, -7.622113e-08, -7.638929e-08, 
    -7.654739e-08, -7.666784e-08, -7.674839e-08, -7.682777e-08, 
    -7.706788e-08, -7.719501e-08, -7.747953e-08, -7.742823e-08, 
    -7.751517e-08, -7.759827e-08, -7.773771e-08, -7.771477e-08, 
    -7.777619e-08, -7.75129e-08, -7.768788e-08, -7.739899e-08, -7.747801e-08, 
    -7.684923e-08, -7.66097e-08, -7.650777e-08, -7.641862e-08, -7.620162e-08, 
    -7.635147e-08, -7.629239e-08, -7.643295e-08, -7.652225e-08, 
    -7.647809e-08, -7.67506e-08, -7.664466e-08, -7.720254e-08, -7.696229e-08, 
    -7.758857e-08, -7.743876e-08, -7.762448e-08, -7.752973e-08, 
    -7.769207e-08, -7.754596e-08, -7.779906e-08, -7.785415e-08, -7.78165e-08, 
    -7.796114e-08, -7.753786e-08, -7.770043e-08, -7.647685e-08, 
    -7.648405e-08, -7.651761e-08, -7.637008e-08, -7.636106e-08, 
    -7.622587e-08, -7.634618e-08, -7.639739e-08, -7.652743e-08, 
    -7.660432e-08, -7.667741e-08, -7.683809e-08, -7.701749e-08, -7.72683e-08, 
    -7.744847e-08, -7.75692e-08, -7.749518e-08, -7.756054e-08, -7.748747e-08, 
    -7.745323e-08, -7.78335e-08, -7.761999e-08, -7.794034e-08, -7.792262e-08, 
    -7.777765e-08, -7.792462e-08, -7.648911e-08, -7.644767e-08, 
    -7.630373e-08, -7.641638e-08, -7.621115e-08, -7.632602e-08, 
    -7.639206e-08, -7.664685e-08, -7.670285e-08, -7.675474e-08, 
    -7.685723e-08, -7.698873e-08, -7.721936e-08, -7.741998e-08, -7.76031e-08, 
    -7.758969e-08, -7.759441e-08, -7.76353e-08, -7.7534e-08, -7.765193e-08, 
    -7.767171e-08, -7.761997e-08, -7.792025e-08, -7.783448e-08, 
    -7.792224e-08, -7.78664e-08, -7.646114e-08, -7.653087e-08, -7.649319e-08, 
    -7.656404e-08, -7.651412e-08, -7.673605e-08, -7.680259e-08, 
    -7.711383e-08, -7.698614e-08, -7.718939e-08, -7.70068e-08, -7.703915e-08, 
    -7.719597e-08, -7.701667e-08, -7.74089e-08, -7.714296e-08, -7.763688e-08, 
    -7.737135e-08, -7.765352e-08, -7.760231e-08, -7.768711e-08, 
    -7.776304e-08, -7.785858e-08, -7.803479e-08, -7.7994e-08, -7.814135e-08, 
    -7.663483e-08, -7.672524e-08, -7.671731e-08, -7.681193e-08, -7.68819e-08, 
    -7.703356e-08, -7.727672e-08, -7.71853e-08, -7.735314e-08, -7.738683e-08, 
    -7.713184e-08, -7.728839e-08, -7.678577e-08, -7.686698e-08, 
    -7.681864e-08, -7.664195e-08, -7.720634e-08, -7.691673e-08, 
    -7.745144e-08, -7.729462e-08, -7.775221e-08, -7.752466e-08, 
    -7.797154e-08, -7.816244e-08, -7.834216e-08, -7.855203e-08, 
    -7.677461e-08, -7.671318e-08, -7.682319e-08, -7.697533e-08, 
    -7.711654e-08, -7.730418e-08, -7.732339e-08, -7.735854e-08, 
    -7.744958e-08, -7.752611e-08, -7.736963e-08, -7.754529e-08, 
    -7.688577e-08, -7.723148e-08, -7.668994e-08, -7.685301e-08, 
    -7.696638e-08, -7.691667e-08, -7.717485e-08, -7.723568e-08, 
    -7.748282e-08, -7.735509e-08, -7.811531e-08, -7.777906e-08, 
    -7.871185e-08, -7.845127e-08, -7.669171e-08, -7.677441e-08, 
    -7.706215e-08, -7.692525e-08, -7.731672e-08, -7.741303e-08, 
    -7.749135e-08, -7.75914e-08, -7.760222e-08, -7.76615e-08, -7.756436e-08, 
    -7.765767e-08, -7.730458e-08, -7.74624e-08, -7.702928e-08, -7.713471e-08, 
    -7.708622e-08, -7.703301e-08, -7.719722e-08, -7.737208e-08, 
    -7.737585e-08, -7.743191e-08, -7.758979e-08, -7.731831e-08, 
    -7.815863e-08, -7.763973e-08, -7.686458e-08, -7.702379e-08, 
    -7.704657e-08, -7.698489e-08, -7.740338e-08, -7.725177e-08, 
    -7.766006e-08, -7.754974e-08, -7.77305e-08, -7.764068e-08, -7.762746e-08, 
    -7.75121e-08, -7.744025e-08, -7.725872e-08, -7.711099e-08, -7.699384e-08, 
    -7.702109e-08, -7.714976e-08, -7.738279e-08, -7.760318e-08, 
    -7.755491e-08, -7.771676e-08, -7.728835e-08, -7.7468e-08, -7.739856e-08, 
    -7.757962e-08, -7.718286e-08, -7.752063e-08, -7.709649e-08, 
    -7.713369e-08, -7.724876e-08, -7.748016e-08, -7.75314e-08, -7.758604e-08, 
    -7.755232e-08, -7.738871e-08, -7.736191e-08, -7.724597e-08, 
    -7.721394e-08, -7.71256e-08, -7.705243e-08, -7.711927e-08, -7.718945e-08, 
    -7.738879e-08, -7.756837e-08, -7.776411e-08, -7.781203e-08, 
    -7.804059e-08, -7.785449e-08, -7.816151e-08, -7.790043e-08, 
    -7.835236e-08, -7.754026e-08, -7.789281e-08, -7.725401e-08, 
    -7.732286e-08, -7.744735e-08, -7.773286e-08, -7.757877e-08, 
    -7.775899e-08, -7.736087e-08, -7.715419e-08, -7.710074e-08, 
    -7.700096e-08, -7.710302e-08, -7.709473e-08, -7.719238e-08, -7.7161e-08, 
    -7.739541e-08, -7.72695e-08, -7.762712e-08, -7.775758e-08, -7.812591e-08, 
    -7.835159e-08, -7.858132e-08, -7.86827e-08, -7.871355e-08, -7.872645e-08 ;

 NET_NMIN =
  1.074108e-08, 1.077048e-08, 1.076477e-08, 1.078847e-08, 1.077532e-08, 
    1.079084e-08, 1.074704e-08, 1.077164e-08, 1.075594e-08, 1.074373e-08, 
    1.083445e-08, 1.078953e-08, 1.088112e-08, 1.085248e-08, 1.092442e-08, 
    1.087666e-08, 1.093404e-08, 1.092304e-08, 1.095616e-08, 1.094667e-08, 
    1.098901e-08, 1.096054e-08, 1.101096e-08, 1.098222e-08, 1.098671e-08, 
    1.09596e-08, 1.079858e-08, 1.082886e-08, 1.079678e-08, 1.08011e-08, 
    1.079916e-08, 1.077559e-08, 1.076371e-08, 1.073884e-08, 1.074335e-08, 
    1.076162e-08, 1.080304e-08, 1.078899e-08, 1.082441e-08, 1.082361e-08, 
    1.086304e-08, 1.084526e-08, 1.091151e-08, 1.089268e-08, 1.094707e-08, 
    1.093339e-08, 1.094643e-08, 1.094248e-08, 1.094648e-08, 1.092642e-08, 
    1.093501e-08, 1.091737e-08, 1.084859e-08, 1.086881e-08, 1.08085e-08, 
    1.077222e-08, 1.074812e-08, 1.073102e-08, 1.073343e-08, 1.073804e-08, 
    1.076173e-08, 1.0784e-08, 1.080097e-08, 1.081232e-08, 1.08235e-08, 
    1.085732e-08, 1.087523e-08, 1.091531e-08, 1.090808e-08, 1.092033e-08, 
    1.093203e-08, 1.095168e-08, 1.094845e-08, 1.09571e-08, 1.092001e-08, 
    1.094466e-08, 1.090396e-08, 1.091509e-08, 1.082652e-08, 1.079278e-08, 
    1.077842e-08, 1.076586e-08, 1.073529e-08, 1.07564e-08, 1.074808e-08, 
    1.076788e-08, 1.078046e-08, 1.077424e-08, 1.081263e-08, 1.07977e-08, 
    1.087629e-08, 1.084245e-08, 1.093067e-08, 1.090957e-08, 1.093573e-08, 
    1.092238e-08, 1.094525e-08, 1.092467e-08, 1.096032e-08, 1.096808e-08, 
    1.096278e-08, 1.098315e-08, 1.092353e-08, 1.094643e-08, 1.077407e-08, 
    1.077508e-08, 1.077981e-08, 1.075903e-08, 1.075775e-08, 1.073871e-08, 
    1.075566e-08, 1.076287e-08, 1.078119e-08, 1.079202e-08, 1.080232e-08, 
    1.082495e-08, 1.085022e-08, 1.088555e-08, 1.091093e-08, 1.092794e-08, 
    1.091751e-08, 1.092672e-08, 1.091643e-08, 1.09116e-08, 1.096517e-08, 
    1.093509e-08, 1.098022e-08, 1.097773e-08, 1.09573e-08, 1.097801e-08, 
    1.077579e-08, 1.076995e-08, 1.074968e-08, 1.076555e-08, 1.073664e-08, 
    1.075282e-08, 1.076212e-08, 1.079801e-08, 1.08059e-08, 1.081321e-08, 
    1.082765e-08, 1.084617e-08, 1.087866e-08, 1.090692e-08, 1.093272e-08, 
    1.093083e-08, 1.093149e-08, 1.093725e-08, 1.092298e-08, 1.093959e-08, 
    1.094238e-08, 1.093509e-08, 1.097739e-08, 1.096531e-08, 1.097767e-08, 
    1.096981e-08, 1.077185e-08, 1.078168e-08, 1.077637e-08, 1.078635e-08, 
    1.077932e-08, 1.081058e-08, 1.081995e-08, 1.086379e-08, 1.084581e-08, 
    1.087444e-08, 1.084872e-08, 1.085327e-08, 1.087537e-08, 1.085011e-08, 
    1.090536e-08, 1.08679e-08, 1.093747e-08, 1.090007e-08, 1.093982e-08, 
    1.09326e-08, 1.094455e-08, 1.095525e-08, 1.09687e-08, 1.099353e-08, 
    1.098778e-08, 1.100854e-08, 1.079632e-08, 1.080906e-08, 1.080794e-08, 
    1.082127e-08, 1.083112e-08, 1.085249e-08, 1.088674e-08, 1.087386e-08, 
    1.089751e-08, 1.090225e-08, 1.086633e-08, 1.088838e-08, 1.081758e-08, 
    1.082902e-08, 1.082221e-08, 1.079732e-08, 1.087682e-08, 1.083603e-08, 
    1.091135e-08, 1.088926e-08, 1.095372e-08, 1.092167e-08, 1.098461e-08, 
    1.101151e-08, 1.103682e-08, 1.106639e-08, 1.081601e-08, 1.080736e-08, 
    1.082285e-08, 1.084429e-08, 1.086418e-08, 1.089061e-08, 1.089331e-08, 
    1.089826e-08, 1.091109e-08, 1.092187e-08, 1.089983e-08, 1.092457e-08, 
    1.083167e-08, 1.088037e-08, 1.080408e-08, 1.082705e-08, 1.084302e-08, 
    1.083602e-08, 1.087239e-08, 1.088096e-08, 1.091577e-08, 1.089778e-08, 
    1.100487e-08, 1.09575e-08, 1.10889e-08, 1.105219e-08, 1.080433e-08, 
    1.081598e-08, 1.085651e-08, 1.083723e-08, 1.089237e-08, 1.090594e-08, 
    1.091697e-08, 1.093107e-08, 1.093259e-08, 1.094094e-08, 1.092726e-08, 
    1.09404e-08, 1.089067e-08, 1.091289e-08, 1.085188e-08, 1.086674e-08, 
    1.08599e-08, 1.085241e-08, 1.087554e-08, 1.090017e-08, 1.09007e-08, 
    1.09086e-08, 1.093084e-08, 1.08926e-08, 1.101097e-08, 1.093787e-08, 
    1.082868e-08, 1.085111e-08, 1.085432e-08, 1.084563e-08, 1.090458e-08, 
    1.088323e-08, 1.094074e-08, 1.09252e-08, 1.095066e-08, 1.093801e-08, 
    1.093615e-08, 1.09199e-08, 1.090978e-08, 1.08842e-08, 1.086339e-08, 
    1.084689e-08, 1.085073e-08, 1.086886e-08, 1.090168e-08, 1.093273e-08, 
    1.092593e-08, 1.094873e-08, 1.088838e-08, 1.091368e-08, 1.09039e-08, 
    1.092941e-08, 1.087352e-08, 1.09211e-08, 1.086135e-08, 1.086659e-08, 
    1.08828e-08, 1.09154e-08, 1.092261e-08, 1.093031e-08, 1.092556e-08, 
    1.090252e-08, 1.089874e-08, 1.088241e-08, 1.08779e-08, 1.086545e-08, 
    1.085515e-08, 1.086456e-08, 1.087445e-08, 1.090253e-08, 1.092782e-08, 
    1.09554e-08, 1.096215e-08, 1.099434e-08, 1.096813e-08, 1.101138e-08, 
    1.09746e-08, 1.103826e-08, 1.092386e-08, 1.097353e-08, 1.088354e-08, 
    1.089324e-08, 1.091078e-08, 1.095099e-08, 1.092929e-08, 1.095467e-08, 
    1.089859e-08, 1.086948e-08, 1.086195e-08, 1.08479e-08, 1.086227e-08, 
    1.08611e-08, 1.087486e-08, 1.087044e-08, 1.090346e-08, 1.088572e-08, 
    1.09361e-08, 1.095448e-08, 1.100636e-08, 1.103815e-08, 1.107051e-08, 
    1.108479e-08, 1.108914e-08, 1.109096e-08 ;

 NFIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NFIX_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 OCDEP =
  6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14 ;

 O_SCALAR =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 PARVEGLN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PBOT =
  100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5 ;

 PCH4 =
  0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627 ;

 PCO2 =
  28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399 ;

 PCT_LANDUNIT =
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PCT_NAT_PFT =
  13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892,
  55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_CTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_NTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PLANT_NDEMAND =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 POTENTIAL_IMMOB =
  5.20049e-14, 5.213718e-14, 5.211149e-14, 5.221808e-14, 5.215898e-14, 
    5.222874e-14, 5.203175e-14, 5.214241e-14, 5.207179e-14, 5.201684e-14, 
    5.242459e-14, 5.222284e-14, 5.263398e-14, 5.250555e-14, 5.282794e-14, 
    5.261398e-14, 5.287104e-14, 5.282182e-14, 5.297001e-14, 5.292758e-14, 
    5.311679e-14, 5.298958e-14, 5.321482e-14, 5.308646e-14, 5.310653e-14, 
    5.298538e-14, 5.226351e-14, 5.239947e-14, 5.225544e-14, 5.227484e-14, 
    5.226615e-14, 5.216018e-14, 5.210672e-14, 5.199481e-14, 5.201514e-14, 
    5.209735e-14, 5.228357e-14, 5.222042e-14, 5.237959e-14, 5.2376e-14, 
    5.255292e-14, 5.247318e-14, 5.277016e-14, 5.268585e-14, 5.292935e-14, 
    5.286815e-14, 5.292647e-14, 5.290879e-14, 5.29267e-14, 5.283694e-14, 
    5.28754e-14, 5.27964e-14, 5.248811e-14, 5.257879e-14, 5.23081e-14, 
    5.214496e-14, 5.203659e-14, 5.19596e-14, 5.197049e-14, 5.199123e-14, 
    5.209783e-14, 5.219801e-14, 5.227428e-14, 5.232526e-14, 5.237548e-14, 
    5.252724e-14, 5.260758e-14, 5.278718e-14, 5.275483e-14, 5.280965e-14, 
    5.286207e-14, 5.294995e-14, 5.29355e-14, 5.297419e-14, 5.280824e-14, 
    5.291854e-14, 5.273639e-14, 5.278623e-14, 5.238897e-14, 5.223747e-14, 
    5.217287e-14, 5.211642e-14, 5.197886e-14, 5.207386e-14, 5.203642e-14, 
    5.212552e-14, 5.218208e-14, 5.215412e-14, 5.232666e-14, 5.225961e-14, 
    5.261234e-14, 5.246054e-14, 5.285596e-14, 5.276147e-14, 5.28786e-14, 
    5.281885e-14, 5.292119e-14, 5.282909e-14, 5.29886e-14, 5.302328e-14, 
    5.299958e-14, 5.309065e-14, 5.282398e-14, 5.292645e-14, 5.215333e-14, 
    5.215789e-14, 5.217915e-14, 5.208566e-14, 5.207994e-14, 5.199425e-14, 
    5.207052e-14, 5.210297e-14, 5.218537e-14, 5.223406e-14, 5.228033e-14, 
    5.2382e-14, 5.249542e-14, 5.265388e-14, 5.27676e-14, 5.284375e-14, 
    5.279707e-14, 5.283828e-14, 5.279221e-14, 5.277061e-14, 5.301028e-14, 
    5.287575e-14, 5.307756e-14, 5.306641e-14, 5.29751e-14, 5.306766e-14, 
    5.216109e-14, 5.213484e-14, 5.204361e-14, 5.211501e-14, 5.198491e-14, 
    5.205773e-14, 5.209958e-14, 5.226097e-14, 5.229644e-14, 5.232927e-14, 
    5.239412e-14, 5.247727e-14, 5.262297e-14, 5.274961e-14, 5.286512e-14, 
    5.285667e-14, 5.285964e-14, 5.288541e-14, 5.282154e-14, 5.28959e-14, 
    5.290836e-14, 5.287575e-14, 5.306491e-14, 5.301091e-14, 5.306617e-14, 
    5.303102e-14, 5.214338e-14, 5.218755e-14, 5.216368e-14, 5.220855e-14, 
    5.217693e-14, 5.231742e-14, 5.235951e-14, 5.25563e-14, 5.247562e-14, 
    5.260404e-14, 5.248868e-14, 5.250912e-14, 5.260816e-14, 5.249493e-14, 
    5.27426e-14, 5.257469e-14, 5.288642e-14, 5.271889e-14, 5.28969e-14, 
    5.286462e-14, 5.291808e-14, 5.296591e-14, 5.302609e-14, 5.313698e-14, 
    5.311132e-14, 5.320402e-14, 5.225338e-14, 5.23106e-14, 5.230559e-14, 
    5.236546e-14, 5.240972e-14, 5.250561e-14, 5.26592e-14, 5.260147e-14, 
    5.270746e-14, 5.272871e-14, 5.256771e-14, 5.266656e-14, 5.23489e-14, 
    5.240025e-14, 5.23697e-14, 5.225788e-14, 5.261474e-14, 5.243172e-14, 
    5.276947e-14, 5.26705e-14, 5.295909e-14, 5.281563e-14, 5.309718e-14, 
    5.321724e-14, 5.333024e-14, 5.346198e-14, 5.234185e-14, 5.230298e-14, 
    5.237259e-14, 5.246877e-14, 5.255804e-14, 5.267654e-14, 5.268867e-14, 
    5.271085e-14, 5.27683e-14, 5.281657e-14, 5.271783e-14, 5.282868e-14, 
    5.241209e-14, 5.263062e-14, 5.228825e-14, 5.239142e-14, 5.246312e-14, 
    5.24317e-14, 5.259488e-14, 5.26333e-14, 5.278925e-14, 5.270868e-14, 
    5.318759e-14, 5.297597e-14, 5.356227e-14, 5.339874e-14, 5.228939e-14, 
    5.234173e-14, 5.252365e-14, 5.243713e-14, 5.268446e-14, 5.274524e-14, 
    5.279465e-14, 5.285774e-14, 5.286457e-14, 5.290192e-14, 5.284069e-14, 
    5.289952e-14, 5.267679e-14, 5.277638e-14, 5.250291e-14, 5.256951e-14, 
    5.253889e-14, 5.250527e-14, 5.260901e-14, 5.271937e-14, 5.272178e-14, 
    5.275714e-14, 5.285662e-14, 5.268546e-14, 5.321478e-14, 5.288811e-14, 
    5.239877e-14, 5.24994e-14, 5.251382e-14, 5.247485e-14, 5.273915e-14, 
    5.264345e-14, 5.290102e-14, 5.283148e-14, 5.294541e-14, 5.288881e-14, 
    5.288047e-14, 5.280774e-14, 5.276241e-14, 5.264783e-14, 5.255453e-14, 
    5.24805e-14, 5.249773e-14, 5.257902e-14, 5.272613e-14, 5.286516e-14, 
    5.283472e-14, 5.293676e-14, 5.266654e-14, 5.277991e-14, 5.273609e-14, 
    5.285031e-14, 5.259993e-14, 5.281303e-14, 5.254538e-14, 5.256888e-14, 
    5.264155e-14, 5.278756e-14, 5.281991e-14, 5.285435e-14, 5.283311e-14, 
    5.272988e-14, 5.271298e-14, 5.263979e-14, 5.261956e-14, 5.256377e-14, 
    5.251753e-14, 5.255976e-14, 5.260409e-14, 5.272994e-14, 5.284321e-14, 
    5.296658e-14, 5.299677e-14, 5.314058e-14, 5.302346e-14, 5.321659e-14, 
    5.305232e-14, 5.333657e-14, 5.282544e-14, 5.304758e-14, 5.264487e-14, 
    5.268834e-14, 5.276687e-14, 5.294686e-14, 5.284978e-14, 5.296333e-14, 
    5.271232e-14, 5.25818e-14, 5.254806e-14, 5.2485e-14, 5.254951e-14, 
    5.254426e-14, 5.260595e-14, 5.258614e-14, 5.273412e-14, 5.265465e-14, 
    5.288025e-14, 5.296245e-14, 5.319429e-14, 5.333613e-14, 5.34804e-14, 
    5.3544e-14, 5.356335e-14, 5.357144e-14 ;

 POT_F_DENIT =
  2.431536e-36, 2.080171e-35, 1.377042e-35, 7.51097e-35, 2.945023e-35, 
    8.881373e-35, 3.775778e-36, 2.262524e-35, 7.249973e-36, 2.95697e-36, 
    1.808846e-33, 8.093939e-35, 3.946951e-32, 6.045991e-33, 6.088165e-31, 
    2.958383e-32, 1.100823e-30, 5.589807e-31, 4.199307e-30, 2.372932e-30, 
    2.909635e-29, 5.454859e-30, 1.022441e-28, 1.959256e-29, 2.545516e-29, 
    5.157598e-30, 1.529097e-34, 1.237951e-33, 1.348288e-34, 1.824726e-34, 
    1.593225e-34, 3.003121e-35, 1.276494e-35, 2.058065e-36, 2.875827e-36, 
    1.096847e-35, 2.089805e-34, 7.787286e-35, 9.12848e-34, 8.643058e-34, 
    1.214609e-32, 3.736812e-33, 2.72498e-31, 8.287591e-32, 2.430399e-30, 
    1.057477e-30, 2.337914e-30, 1.840018e-30, 2.345202e-30, 6.887896e-31, 
    1.167867e-30, 3.928743e-31, 4.667509e-33, 1.773161e-32, 3.054395e-34, 
    2.358835e-35, 4.088082e-36, 1.149436e-36, 1.377033e-36, 1.940986e-36, 
    1.105402e-35, 5.469746e-35, 1.807634e-34, 3.977145e-34, 8.575428e-34, 
    8.34156e-33, 2.69561e-32, 3.457341e-31, 2.197837e-31, 4.725023e-31, 
    9.728318e-31, 3.209095e-30, 2.641e-30, 4.442478e-30, 4.630589e-31, 
    2.100941e-30, 1.695494e-31, 3.410151e-31, 1.055934e-33, 1.017697e-34, 
    3.678611e-35, 1.490986e-35, 1.581801e-36, 7.500951e-36, 4.076749e-36, 
    1.724691e-35, 4.25128e-35, 2.724771e-35, 4.063328e-34, 1.438516e-34, 
    2.887758e-32, 3.095547e-33, 8.94634e-31, 2.41262e-31, 1.219711e-30, 
    5.363627e-31, 2.177187e-30, 6.179375e-31, 5.384613e-30, 8.539326e-30, 
    6.233685e-30, 2.06851e-29, 5.758325e-31, 2.338045e-30, 2.691009e-35, 
    2.894075e-35, 4.057476e-35, 9.080108e-36, 8.27686e-36, 2.039305e-36, 
    7.101458e-36, 1.200639e-35, 4.477733e-35, 9.648016e-35, 1.986333e-34, 
    9.472638e-34, 5.205024e-33, 5.251311e-32, 2.62879e-31, 7.563291e-31, 
    3.964653e-31, 7.014704e-31, 3.705541e-31, 2.741184e-31, 7.187649e-30, 
    1.173657e-30, 1.743426e-29, 1.506449e-29, 4.497641e-30, 1.531475e-29, 
    3.04559e-35, 2.002432e-35, 4.583814e-36, 1.456866e-35, 1.747991e-36, 
    5.770927e-36, 1.137196e-35, 1.470528e-34, 2.549317e-34, 4.230895e-34, 
    1.138245e-33, 3.971221e-33, 3.365823e-32, 2.043549e-31, 1.014278e-30, 
    9.032062e-31, 9.408806e-31, 1.338794e-30, 5.567699e-31, 1.544329e-30, 
    1.829777e-30, 1.173308e-30, 1.477218e-29, 7.244453e-30, 1.501769e-29, 
    9.453937e-30, 2.295419e-35, 4.635668e-35, 3.173496e-35, 6.461318e-35, 
    3.918533e-35, 3.528461e-34, 6.730773e-34, 1.277267e-32, 3.875749e-33, 
    2.559798e-32, 4.706361e-33, 6.374028e-33, 2.720699e-32, 5.162966e-33, 
    1.852806e-31, 1.671785e-32, 1.357209e-30, 1.32692e-31, 1.565558e-30, 
    1.007367e-30, 2.086567e-30, 3.976023e-30, 8.858512e-30, 3.775103e-29, 
    2.707442e-29, 8.909693e-29, 1.30531e-34, 3.17464e-34, 2.936628e-34, 
    7.362291e-34, 1.441659e-33, 6.048335e-33, 5.665552e-32, 2.464709e-32, 
    1.126559e-31, 1.521901e-31, 1.507442e-32, 6.296677e-32, 5.718368e-34, 
    1.250379e-33, 7.855341e-34, 1.400796e-34, 2.989184e-32, 2.010164e-33, 
    2.698833e-31, 6.659578e-32, 3.628413e-30, 5.134083e-31, 2.252845e-29, 
    1.054976e-28, 4.337753e-28, 2.162218e-27, 5.131526e-34, 2.820386e-34, 
    8.205746e-34, 3.501788e-33, 1.309011e-32, 7.259584e-32, 8.627697e-32, 
    1.182309e-31, 2.654278e-31, 5.197211e-31, 1.305896e-31, 6.143558e-31, 
    1.497649e-33, 3.758781e-32, 2.246509e-34, 1.09386e-33, 3.217284e-33, 
    2.008247e-33, 2.239435e-32, 3.903964e-32, 3.558205e-31, 1.146259e-31, 
    7.23638e-29, 4.552815e-30, 7.106188e-27, 1.00624e-27, 2.285472e-34, 
    5.120692e-34, 7.901357e-33, 2.178861e-33, 8.125475e-32, 1.921216e-31, 
    3.833498e-31, 9.169636e-31, 1.006659e-30, 1.676492e-30, 7.251408e-31, 
    1.62218e-30, 7.285792e-32, 2.972194e-31, 5.810477e-33, 1.548275e-32, 
    9.881065e-33, 6.016816e-33, 2.748668e-32, 1.334958e-31, 1.379941e-31, 
    2.271224e-31, 9.0572e-31, 8.242193e-32, 1.024441e-28, 1.392712e-30, 
    1.22124e-33, 5.522901e-33, 6.830898e-33, 3.829655e-33, 1.76336e-31, 
    4.519103e-32, 1.655817e-30, 6.386244e-31, 3.018376e-30, 1.402101e-30, 
    1.25149e-30, 4.59802e-31, 2.444659e-31, 4.81349e-32, 1.243548e-32, 
    4.166146e-33, 5.380952e-33, 1.778853e-32, 1.468531e-31, 1.015282e-30, 
    6.682074e-31, 2.686088e-30, 6.2921e-32, 3.123257e-31, 1.689693e-31, 
    8.278788e-31, 2.41056e-32, 4.962282e-31, 1.086891e-32, 1.533495e-32, 
    4.397302e-32, 3.477105e-31, 5.442648e-31, 8.753326e-31, 6.531403e-31, 
    1.547918e-31, 1.218636e-31, 4.286784e-32, 3.203159e-32, 1.422964e-32, 
    7.213664e-33, 1.34234e-32, 2.560963e-32, 1.548728e-31, 7.510358e-31, 
    4.012579e-30, 6.003471e-30, 3.959985e-29, 8.568919e-30, 1.048367e-28, 
    1.256413e-29, 4.701216e-28, 5.885199e-31, 1.178497e-29, 4.611026e-32, 
    8.586307e-32, 2.603937e-31, 3.081409e-30, 8.217949e-31, 3.843672e-30, 
    1.207228e-31, 1.853259e-32, 1.130717e-32, 4.455016e-33, 1.154876e-32, 
    1.069319e-32, 2.629645e-32, 1.971957e-32, 1.642661e-31, 5.306551e-32, 
    1.247989e-30, 3.797551e-30, 7.874024e-29, 4.669595e-28, 2.693259e-27, 
    5.730218e-27, 7.194341e-27, 7.90995e-27 ;

 POT_F_NIT =
  5.751129e-11, 5.782231e-11, 5.77618e-11, 5.801307e-11, 5.787363e-11, 
    5.803824e-11, 5.757428e-11, 5.783463e-11, 5.766837e-11, 5.753924e-11, 
    5.850205e-11, 5.802427e-11, 5.900044e-11, 5.86943e-11, 5.946479e-11, 
    5.895273e-11, 5.956829e-11, 5.945003e-11, 5.98064e-11, 5.97042e-11, 
    6.016099e-11, 5.985359e-11, 6.039847e-11, 6.008753e-11, 6.013609e-11, 
    5.984342e-11, 5.812035e-11, 5.844249e-11, 5.810127e-11, 5.814715e-11, 
    5.812656e-11, 5.787647e-11, 5.77506e-11, 5.748753e-11, 5.753525e-11, 
    5.77285e-11, 5.816776e-11, 5.80185e-11, 5.839507e-11, 5.838655e-11, 
    5.880704e-11, 5.861727e-11, 5.932612e-11, 5.912426e-11, 5.970846e-11, 
    5.956128e-11, 5.970153e-11, 5.965898e-11, 5.970206e-11, 5.948629e-11, 
    5.957868e-11, 5.938899e-11, 5.865284e-11, 5.886876e-11, 5.822581e-11, 
    5.784069e-11, 5.758565e-11, 5.740496e-11, 5.743048e-11, 5.747915e-11, 
    5.772962e-11, 5.79656e-11, 5.814573e-11, 5.826634e-11, 5.838532e-11, 
    5.874599e-11, 5.89374e-11, 5.936694e-11, 5.928936e-11, 5.942084e-11, 
    5.954665e-11, 5.975806e-11, 5.972325e-11, 5.981646e-11, 5.941738e-11, 
    5.968245e-11, 5.924514e-11, 5.936459e-11, 5.841757e-11, 5.805878e-11, 
    5.790644e-11, 5.777337e-11, 5.745011e-11, 5.767324e-11, 5.758522e-11, 
    5.779474e-11, 5.792804e-11, 5.786209e-11, 5.826964e-11, 5.811103e-11, 
    5.894874e-11, 5.858724e-11, 5.953196e-11, 5.930527e-11, 5.958635e-11, 
    5.944285e-11, 5.968881e-11, 5.946742e-11, 5.985118e-11, 5.993488e-11, 
    5.987766e-11, 6.009759e-11, 5.945513e-11, 5.970146e-11, 5.786027e-11, 
    5.787102e-11, 5.792112e-11, 5.770098e-11, 5.768752e-11, 5.748619e-11, 
    5.766532e-11, 5.774168e-11, 5.793577e-11, 5.805068e-11, 5.816003e-11, 
    5.840078e-11, 5.867018e-11, 5.904788e-11, 5.931994e-11, 5.950262e-11, 
    5.939058e-11, 5.948948e-11, 5.937891e-11, 5.932712e-11, 5.990348e-11, 
    5.957952e-11, 6.006592e-11, 6.003897e-11, 5.981864e-11, 6.004199e-11, 
    5.787856e-11, 5.781669e-11, 5.76021e-11, 5.777e-11, 5.746427e-11, 
    5.763529e-11, 5.773371e-11, 5.81143e-11, 5.819811e-11, 5.827582e-11, 
    5.842948e-11, 5.862694e-11, 5.897407e-11, 5.927687e-11, 5.955395e-11, 
    5.953362e-11, 5.954078e-11, 5.960272e-11, 5.944929e-11, 5.962792e-11, 
    5.96579e-11, 5.957948e-11, 6.003534e-11, 5.990495e-11, 6.003838e-11, 
    5.995345e-11, 5.78368e-11, 5.794092e-11, 5.788463e-11, 5.799048e-11, 
    5.791588e-11, 5.824784e-11, 5.834754e-11, 5.881512e-11, 5.862304e-11, 
    5.89289e-11, 5.865408e-11, 5.870273e-11, 5.893881e-11, 5.866892e-11, 
    5.926011e-11, 5.885894e-11, 5.960512e-11, 5.920338e-11, 5.963033e-11, 
    5.955271e-11, 5.968125e-11, 5.979645e-11, 5.994157e-11, 6.02097e-11, 
    6.014756e-11, 6.037214e-11, 5.809632e-11, 5.823166e-11, 5.821976e-11, 
    5.836154e-11, 5.846651e-11, 5.869434e-11, 5.906056e-11, 5.892273e-11, 
    5.91759e-11, 5.922678e-11, 5.884219e-11, 5.907815e-11, 5.832228e-11, 
    5.844406e-11, 5.837156e-11, 5.81069e-11, 5.895439e-11, 5.851873e-11, 
    5.932438e-11, 5.908751e-11, 5.978e-11, 5.943512e-11, 6.011336e-11, 
    6.04043e-11, 6.067884e-11, 6.100024e-11, 5.83056e-11, 5.821357e-11, 
    5.837842e-11, 5.860681e-11, 5.881918e-11, 5.910199e-11, 5.913098e-11, 
    5.918403e-11, 5.932159e-11, 5.943736e-11, 5.920077e-11, 5.946638e-11, 
    5.847227e-11, 5.899228e-11, 5.81787e-11, 5.84231e-11, 5.859329e-11, 
    5.851863e-11, 5.890693e-11, 5.89986e-11, 5.937181e-11, 5.917876e-11, 
    6.033238e-11, 5.982073e-11, 6.124556e-11, 6.084582e-11, 5.818141e-11, 
    5.830528e-11, 5.873731e-11, 5.853158e-11, 5.91209e-11, 5.926637e-11, 
    5.938476e-11, 5.953622e-11, 5.955259e-11, 5.964243e-11, 5.949524e-11, 
    5.963662e-11, 5.910255e-11, 5.934093e-11, 5.868784e-11, 5.884647e-11, 
    5.877347e-11, 5.869343e-11, 5.894061e-11, 5.920443e-11, 5.921012e-11, 
    5.929481e-11, 5.953371e-11, 5.912321e-11, 6.039846e-11, 5.960935e-11, 
    5.84405e-11, 5.867962e-11, 5.871387e-11, 5.862115e-11, 5.925176e-11, 
    5.90229e-11, 5.964024e-11, 5.947311e-11, 5.974706e-11, 5.961086e-11, 
    5.959081e-11, 5.941612e-11, 5.930744e-11, 5.903334e-11, 5.881075e-11, 
    5.863454e-11, 5.867549e-11, 5.886912e-11, 5.922059e-11, 5.955399e-11, 
    5.948087e-11, 5.972616e-11, 5.907799e-11, 5.934936e-11, 5.924438e-11, 
    5.951827e-11, 5.891904e-11, 5.942908e-11, 5.878897e-11, 5.884496e-11, 
    5.901835e-11, 5.936782e-11, 5.944533e-11, 5.952806e-11, 5.9477e-11, 
    5.922957e-11, 5.918908e-11, 5.901411e-11, 5.896582e-11, 5.883273e-11, 
    5.872262e-11, 5.88232e-11, 5.89289e-11, 5.922964e-11, 5.950125e-11, 
    5.979802e-11, 5.987078e-11, 6.021847e-11, 5.99353e-11, 6.040284e-11, 
    6.000513e-11, 6.069439e-11, 5.945876e-11, 5.999364e-11, 5.902626e-11, 
    5.913014e-11, 5.93182e-11, 5.975063e-11, 5.951704e-11, 5.979029e-11, 
    5.91875e-11, 5.887579e-11, 5.879532e-11, 5.864523e-11, 5.879874e-11, 
    5.878625e-11, 5.89333e-11, 5.888603e-11, 5.923963e-11, 5.904957e-11, 
    5.959024e-11, 5.978808e-11, 6.034851e-11, 6.069321e-11, 6.104511e-11, 
    6.120073e-11, 6.124814e-11, 6.126796e-11 ;

 PROD100C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHA =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHADE_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Q2M =
  0.0005836726, 0.0005836753, 0.0005836748, 0.000583677, 0.0005836758, 
    0.0005836772, 0.0005836732, 0.0005836755, 0.0005836741, 0.0005836729, 
    0.0005836812, 0.0005836771, 0.0005836816, 0.000583679, 0.0005836857, 
    0.0005836812, 0.0005836866, 0.0005836856, 0.0005836887, 0.0005836879, 
    0.0005836917, 0.0005836891, 0.0005836939, 0.0005836911, 0.0005836915, 
    0.0005836891, 0.000583678, 0.0005836806, 0.0005836778, 0.0005836782, 
    0.000583678, 0.0005836758, 0.0005836747, 0.0005836725, 0.0005836729, 
    0.0005836745, 0.0005836784, 0.0005836771, 0.0005836804, 0.0005836803, 
    0.00058368, 0.0005836823, 0.0005836845, 0.0005836828, 0.0005836879, 
    0.0005836866, 0.0005836878, 0.0005836874, 0.0005836878, 0.0005836859, 
    0.0005836867, 0.0005836851, 0.0005836826, 0.0005836805, 0.0005836789, 
    0.0005836755, 0.0005836733, 0.0005836717, 0.000583672, 0.0005836724, 
    0.0005836745, 0.0005836766, 0.0005836782, 0.0005836793, 0.0005836803, 
    0.0005836794, 0.0005836811, 0.0005836849, 0.0005836842, 0.0005836854, 
    0.0005836865, 0.0005836883, 0.000583688, 0.0005836888, 0.0005836854, 
    0.0005836876, 0.0005836838, 0.0005836849, 0.0005836804, 0.0005836774, 
    0.000583676, 0.0005836749, 0.0005836721, 0.0005836741, 0.0005836733, 
    0.0005836752, 0.0005836763, 0.0005836757, 0.0005836793, 0.0005836779, 
    0.0005836812, 0.000583682, 0.0005836863, 0.0005836844, 0.0005836868, 
    0.0005836856, 0.0005836877, 0.0005836858, 0.0005836891, 0.0005836898, 
    0.0005836893, 0.0005836912, 0.0005836857, 0.0005836878, 0.0005836757, 
    0.0005836758, 0.0005836763, 0.0005836743, 0.0005836742, 0.0005836724, 
    0.000583674, 0.0005836746, 0.0005836764, 0.0005836774, 0.0005836783, 
    0.0005836804, 0.0005836827, 0.0005836821, 0.0005836845, 0.0005836861, 
    0.0005836851, 0.000583686, 0.000583685, 0.0005836846, 0.0005836895, 
    0.0005836867, 0.000583691, 0.0005836908, 0.0005836888, 0.0005836908, 
    0.0005836759, 0.0005836753, 0.0005836734, 0.0005836749, 0.0005836723, 
    0.0005836737, 0.0005836746, 0.0005836779, 0.0005836787, 0.0005836794, 
    0.0005836807, 0.0005836824, 0.0005836815, 0.0005836841, 0.0005836865, 
    0.0005836863, 0.0005836864, 0.0005836869, 0.0005836856, 0.0005836872, 
    0.0005836874, 0.0005836867, 0.0005836907, 0.0005836896, 0.0005836908, 
    0.00058369, 0.0005836755, 0.0005836764, 0.0005836759, 0.0005836769, 
    0.0005836762, 0.0005836791, 0.0005836799, 0.0005836801, 0.0005836824, 
    0.000583681, 0.0005836827, 0.0005836791, 0.000583681, 0.0005836788, 
    0.0005836839, 0.0005836804, 0.000583687, 0.0005836834, 0.0005836872, 
    0.0005836865, 0.0005836876, 0.0005836886, 0.0005836899, 0.0005836922, 
    0.0005836917, 0.0005836936, 0.0005836778, 0.0005836789, 0.0005836789, 
    0.0005836801, 0.000583681, 0.0005836791, 0.0005836822, 0.000583681, 
    0.0005836833, 0.0005836837, 0.0005836803, 0.0005836824, 0.0005836797, 
    0.0005836808, 0.0005836802, 0.0005836778, 0.0005836813, 0.0005836814, 
    0.0005836845, 0.0005836824, 0.0005836885, 0.0005836855, 0.0005836914, 
    0.0005836939, 0.0005836963, 0.000583699, 0.0005836796, 0.0005836788, 
    0.0005836802, 0.0005836822, 0.0005836801, 0.0005836826, 0.0005836828, 
    0.0005836833, 0.0005836845, 0.0005836855, 0.0005836834, 0.0005836858, 
    0.0005836809, 0.0005836816, 0.0005836785, 0.0005836806, 0.0005836821, 
    0.0005836815, 0.0005836809, 0.0005836817, 0.0005836849, 0.0005836833, 
    0.0005836932, 0.0005836888, 0.0005837012, 0.0005836977, 0.0005836785, 
    0.0005836796, 0.0005836794, 0.0005836816, 0.0005836828, 0.000583684, 
    0.0005836851, 0.0005836863, 0.0005836865, 0.0005836873, 0.0005836861, 
    0.0005836873, 0.0005836826, 0.0005836847, 0.000583679, 0.0005836803, 
    0.0005836798, 0.0005836791, 0.0005836812, 0.0005836834, 0.0005836835, 
    0.0005836842, 0.0005836862, 0.0005836828, 0.0005836936, 0.0005836868, 
    0.0005836808, 0.0005836788, 0.0005836792, 0.0005836824, 0.0005836839, 
    0.0005836819, 0.0005836873, 0.0005836858, 0.0005836882, 0.000583687, 
    0.0005836869, 0.0005836854, 0.0005836844, 0.000583682, 0.0005836801, 
    0.0005836825, 0.0005836789, 0.0005836805, 0.0005836836, 0.0005836865, 
    0.0005836859, 0.000583688, 0.0005836824, 0.0005836847, 0.0005836838, 
    0.0005836862, 0.000583681, 0.0005836852, 0.0005836799, 0.0005836803, 
    0.0005836819, 0.0005836848, 0.0005836856, 0.0005836863, 0.0005836859, 
    0.0005836837, 0.0005836833, 0.0005836819, 0.0005836814, 0.0005836803, 
    0.0005836793, 0.0005836802, 0.000583681, 0.0005836837, 0.0005836861, 
    0.0005836886, 0.0005836893, 0.0005836922, 0.0005836897, 0.0005836937, 
    0.0005836902, 0.0005836963, 0.0005836856, 0.0005836902, 0.000583682, 
    0.0005836828, 0.0005836844, 0.0005836881, 0.0005836862, 0.0005836886, 
    0.0005836833, 0.0005836806, 0.0005836799, 0.0005836826, 0.0005836799, 
    0.0005836799, 0.0005836812, 0.0005836808, 0.0005836838, 0.0005836822, 
    0.0005836868, 0.0005836886, 0.0005836934, 0.0005836964, 0.0005836995, 
    0.0005837008, 0.0005837012, 0.0005837014 ;

 QBOT =
  0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045 ;

 QCHARGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_PERCH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_XS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRIP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLOOD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_ICE_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_LIQ_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINFL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QIRRIG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRGWL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QRUNOFF_NODYNLNDUSE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QRUNOFF_R =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QRUNOFF_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QSNOMELT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSOIL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QVEGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QVEGT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RETRANSN =
  4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07 ;

 RETRANSN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RH2M =
  81.18176, 81.18085, 81.18102, 81.1803, 81.18069, 81.18022, 81.18156, 
    81.18082, 81.18129, 81.18166, 81.17892, 81.18027, 81.17705, 81.17792, 
    81.1757, 81.17719, 81.1754, 81.17573, 81.17469, 81.17499, 81.17371, 
    81.17456, 81.17301, 81.1739, 81.17377, 81.17459, 81.17998, 81.1791, 
    81.18003, 81.17991, 81.17996, 81.18069, 81.18107, 81.18181, 81.18167, 
    81.18112, 81.17985, 81.18027, 81.17918, 81.1792, 81.17759, 81.17854, 
    81.17609, 81.17667, 81.17498, 81.17541, 81.175, 81.17512, 81.175, 
    81.17562, 81.17535, 81.1759, 81.17844, 81.17741, 81.17967, 81.18082, 
    81.18153, 81.18205, 81.18198, 81.18184, 81.18112, 81.18042, 81.17989, 
    81.17955, 81.1792, 81.1778, 81.17723, 81.17598, 81.17619, 81.17582, 
    81.17545, 81.17484, 81.17493, 81.17467, 81.17582, 81.17506, 81.17631, 
    81.17597, 81.17918, 81.18015, 81.18063, 81.18098, 81.18192, 81.18128, 
    81.18153, 81.18092, 81.18053, 81.18072, 81.17953, 81.18, 81.17719, 
    81.17863, 81.17549, 81.17614, 81.17533, 81.17574, 81.17504, 81.17567, 
    81.17457, 81.17434, 81.1745, 81.17386, 81.1757, 81.175, 81.18073, 
    81.18069, 81.18055, 81.1812, 81.18124, 81.18182, 81.1813, 81.18108, 
    81.1805, 81.18018, 81.17986, 81.17916, 81.1784, 81.1769, 81.1761, 
    81.17557, 81.17589, 81.17561, 81.17593, 81.17607, 81.17443, 81.17536, 
    81.17395, 81.17403, 81.17467, 81.17402, 81.18067, 81.18085, 81.18148, 
    81.18098, 81.18188, 81.18139, 81.18111, 81.18001, 81.17975, 81.17953, 
    81.17908, 81.1785, 81.17711, 81.17623, 81.17542, 81.17548, 81.17546, 
    81.17529, 81.17573, 81.17521, 81.17513, 81.17535, 81.17403, 81.17441, 
    81.17403, 81.17427, 81.18079, 81.1805, 81.18066, 81.18035, 81.18057, 
    81.17962, 81.17934, 81.17758, 81.17852, 81.17725, 81.17843, 81.17789, 
    81.17725, 81.17798, 81.17629, 81.17746, 81.17528, 81.17648, 81.1752, 
    81.17542, 81.17506, 81.17473, 81.17431, 81.17355, 81.17372, 81.17307, 
    81.18004, 81.17966, 81.17968, 81.17928, 81.17897, 81.17791, 81.17686, 
    81.17725, 81.17651, 81.17637, 81.17747, 81.17681, 81.1794, 81.17905, 
    81.17924, 81.18002, 81.17718, 81.17884, 81.17609, 81.17677, 81.17477, 
    81.17578, 81.17382, 81.17301, 81.17219, 81.1713, 81.17944, 81.1797, 
    81.17922, 81.17858, 81.17755, 81.17673, 81.17664, 81.17649, 81.17609, 
    81.17576, 81.17646, 81.17567, 81.179, 81.17706, 81.17981, 81.17912, 
    81.17861, 81.17883, 81.17729, 81.17702, 81.17596, 81.17651, 81.17322, 
    81.17467, 81.17057, 81.17173, 81.17979, 81.17944, 81.1778, 81.17879, 
    81.17667, 81.17625, 81.17591, 81.17548, 81.17543, 81.17517, 81.17559, 
    81.17519, 81.17673, 81.17604, 81.17793, 81.17747, 81.17767, 81.17791, 
    81.17719, 81.17645, 81.17641, 81.17618, 81.17556, 81.17667, 81.17307, 
    81.17533, 81.17904, 81.17797, 81.17786, 81.17852, 81.1763, 81.17696, 
    81.17518, 81.17565, 81.17487, 81.17526, 81.17532, 81.17582, 81.17614, 
    81.17693, 81.17757, 81.17847, 81.17796, 81.17741, 81.1764, 81.17543, 
    81.17564, 81.17493, 81.1768, 81.17603, 81.17633, 81.17553, 81.17726, 
    81.17585, 81.17763, 81.17747, 81.17697, 81.17599, 81.17574, 81.17551, 
    81.17564, 81.17637, 81.17648, 81.17698, 81.17713, 81.17751, 81.17782, 
    81.17754, 81.17724, 81.17636, 81.17558, 81.17473, 81.17451, 81.17355, 
    81.17436, 81.17307, 81.17421, 81.1722, 81.17574, 81.1742, 81.17694, 
    81.17664, 81.17612, 81.17488, 81.17553, 81.17477, 81.17648, 81.1774, 
    81.17761, 81.17845, 81.1776, 81.17764, 81.17722, 81.17735, 81.17633, 
    81.17688, 81.17532, 81.17477, 81.17315, 81.17217, 81.17113, 81.17069, 
    81.17056, 81.1705 ;

 RH2M_R =
  81.18176, 81.18085, 81.18102, 81.1803, 81.18069, 81.18022, 81.18156, 
    81.18082, 81.18129, 81.18166, 81.17892, 81.18027, 81.17705, 81.17792, 
    81.1757, 81.17719, 81.1754, 81.17573, 81.17469, 81.17499, 81.17371, 
    81.17456, 81.17301, 81.1739, 81.17377, 81.17459, 81.17998, 81.1791, 
    81.18003, 81.17991, 81.17996, 81.18069, 81.18107, 81.18181, 81.18167, 
    81.18112, 81.17985, 81.18027, 81.17918, 81.1792, 81.17759, 81.17854, 
    81.17609, 81.17667, 81.17498, 81.17541, 81.175, 81.17512, 81.175, 
    81.17562, 81.17535, 81.1759, 81.17844, 81.17741, 81.17967, 81.18082, 
    81.18153, 81.18205, 81.18198, 81.18184, 81.18112, 81.18042, 81.17989, 
    81.17955, 81.1792, 81.1778, 81.17723, 81.17598, 81.17619, 81.17582, 
    81.17545, 81.17484, 81.17493, 81.17467, 81.17582, 81.17506, 81.17631, 
    81.17597, 81.17918, 81.18015, 81.18063, 81.18098, 81.18192, 81.18128, 
    81.18153, 81.18092, 81.18053, 81.18072, 81.17953, 81.18, 81.17719, 
    81.17863, 81.17549, 81.17614, 81.17533, 81.17574, 81.17504, 81.17567, 
    81.17457, 81.17434, 81.1745, 81.17386, 81.1757, 81.175, 81.18073, 
    81.18069, 81.18055, 81.1812, 81.18124, 81.18182, 81.1813, 81.18108, 
    81.1805, 81.18018, 81.17986, 81.17916, 81.1784, 81.1769, 81.1761, 
    81.17557, 81.17589, 81.17561, 81.17593, 81.17607, 81.17443, 81.17536, 
    81.17395, 81.17403, 81.17467, 81.17402, 81.18067, 81.18085, 81.18148, 
    81.18098, 81.18188, 81.18139, 81.18111, 81.18001, 81.17975, 81.17953, 
    81.17908, 81.1785, 81.17711, 81.17623, 81.17542, 81.17548, 81.17546, 
    81.17529, 81.17573, 81.17521, 81.17513, 81.17535, 81.17403, 81.17441, 
    81.17403, 81.17427, 81.18079, 81.1805, 81.18066, 81.18035, 81.18057, 
    81.17962, 81.17934, 81.17758, 81.17852, 81.17725, 81.17843, 81.17789, 
    81.17725, 81.17798, 81.17629, 81.17746, 81.17528, 81.17648, 81.1752, 
    81.17542, 81.17506, 81.17473, 81.17431, 81.17355, 81.17372, 81.17307, 
    81.18004, 81.17966, 81.17968, 81.17928, 81.17897, 81.17791, 81.17686, 
    81.17725, 81.17651, 81.17637, 81.17747, 81.17681, 81.1794, 81.17905, 
    81.17924, 81.18002, 81.17718, 81.17884, 81.17609, 81.17677, 81.17477, 
    81.17578, 81.17382, 81.17301, 81.17219, 81.1713, 81.17944, 81.1797, 
    81.17922, 81.17858, 81.17755, 81.17673, 81.17664, 81.17649, 81.17609, 
    81.17576, 81.17646, 81.17567, 81.179, 81.17706, 81.17981, 81.17912, 
    81.17861, 81.17883, 81.17729, 81.17702, 81.17596, 81.17651, 81.17322, 
    81.17467, 81.17057, 81.17173, 81.17979, 81.17944, 81.1778, 81.17879, 
    81.17667, 81.17625, 81.17591, 81.17548, 81.17543, 81.17517, 81.17559, 
    81.17519, 81.17673, 81.17604, 81.17793, 81.17747, 81.17767, 81.17791, 
    81.17719, 81.17645, 81.17641, 81.17618, 81.17556, 81.17667, 81.17307, 
    81.17533, 81.17904, 81.17797, 81.17786, 81.17852, 81.1763, 81.17696, 
    81.17518, 81.17565, 81.17487, 81.17526, 81.17532, 81.17582, 81.17614, 
    81.17693, 81.17757, 81.17847, 81.17796, 81.17741, 81.1764, 81.17543, 
    81.17564, 81.17493, 81.1768, 81.17603, 81.17633, 81.17553, 81.17726, 
    81.17585, 81.17763, 81.17747, 81.17697, 81.17599, 81.17574, 81.17551, 
    81.17564, 81.17637, 81.17648, 81.17698, 81.17713, 81.17751, 81.17782, 
    81.17754, 81.17724, 81.17636, 81.17558, 81.17473, 81.17451, 81.17355, 
    81.17436, 81.17307, 81.17421, 81.1722, 81.17574, 81.1742, 81.17694, 
    81.17664, 81.17612, 81.17488, 81.17553, 81.17477, 81.17648, 81.1774, 
    81.17761, 81.17845, 81.1776, 81.17764, 81.17722, 81.17735, 81.17633, 
    81.17688, 81.17532, 81.17477, 81.17315, 81.17217, 81.17113, 81.17069, 
    81.17056, 81.1705 ;

 RH2M_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 RR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RSCANOPY =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 SABG =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 SABG_PEN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN =
  0.0005333776, 0.000534783, 0.0005345098, 0.000535643, 0.0005350144, 
    0.0005357562, 0.0005336624, 0.0005348384, 0.0005340877, 0.0005335038, 
    0.0005378405, 0.0005356931, 0.0005400709, 0.0005387019, 0.00054214, 
    0.0005398577, 0.0005426001, 0.0005420743, 0.0005436569, 0.0005432035, 
    0.0005452267, 0.000543866, 0.0005462753, 0.0005449018, 0.0005451165, 
    0.0005438208, 0.0005361259, 0.0005375736, 0.00053604, 0.0005362465, 
    0.0005361538, 0.0005350271, 0.0005344591, 0.0005332698, 0.0005334857, 
    0.0005343592, 0.000536339, 0.000535667, 0.0005373603, 0.0005373221, 
    0.0005392063, 0.0005383568, 0.0005415229, 0.0005406232, 0.0005432224, 
    0.0005425687, 0.0005431915, 0.0005430026, 0.0005431938, 0.0005422353, 
    0.0005426459, 0.0005418024, 0.0005385165, 0.0005394827, 0.0005366001, 
    0.0005348657, 0.0005337137, 0.000532896, 0.0005330115, 0.0005332318, 
    0.0005343642, 0.0005354287, 0.0005362397, 0.0005367821, 0.0005373164, 
    0.0005389332, 0.0005397891, 0.0005417045, 0.000541359, 0.0005419443, 
    0.0005425037, 0.0005434423, 0.0005432878, 0.0005437012, 0.0005419287, 
    0.0005431067, 0.0005411617, 0.0005416937, 0.0005374616, 0.0005358486, 
    0.0005351622, 0.0005345618, 0.0005331003, 0.0005341095, 0.0005337116, 
    0.0005346581, 0.0005352593, 0.0005349619, 0.0005367969, 0.0005360834, 
    0.0005398397, 0.0005382221, 0.0005424385, 0.0005414299, 0.00054268, 
    0.0005420421, 0.0005431349, 0.0005421513, 0.0005438551, 0.0005442259, 
    0.0005439724, 0.000544946, 0.0005420964, 0.0005431909, 0.0005349538, 
    0.0005350024, 0.0005352282, 0.0005342347, 0.000534174, 0.0005332635, 
    0.0005340736, 0.0005344185, 0.0005352941, 0.0005358118, 0.0005363039, 
    0.0005373858, 0.0005385936, 0.0005402822, 0.0005414952, 0.0005423079, 
    0.0005418095, 0.0005422494, 0.0005417575, 0.0005415269, 0.0005440867, 
    0.0005426495, 0.0005448058, 0.0005446866, 0.0005437106, 0.0005446998, 
    0.0005350363, 0.0005347572, 0.0005337879, 0.0005345463, 0.0005331642, 
    0.0005339378, 0.0005343825, 0.0005360981, 0.0005364751, 0.0005368245, 
    0.0005375145, 0.0005383999, 0.0005399527, 0.0005413032, 0.000542536, 
    0.0005424456, 0.0005424774, 0.0005427526, 0.0005420705, 0.0005428644, 
    0.0005429975, 0.0005426492, 0.0005446704, 0.0005440931, 0.0005446838, 
    0.0005443078, 0.0005348478, 0.0005353173, 0.0005350635, 0.0005355406, 
    0.0005352044, 0.0005366988, 0.0005371467, 0.0005392423, 0.0005383824, 
    0.0005397509, 0.0005385214, 0.0005387393, 0.0005397951, 0.0005385877, 
    0.0005412285, 0.000539438, 0.0005427632, 0.0005409755, 0.0005428751, 
    0.0005425302, 0.000543101, 0.0005436122, 0.0005442552, 0.0005454413, 
    0.0005451666, 0.0005461585, 0.0005360173, 0.000536626, 0.0005365725, 
    0.0005372096, 0.0005376806, 0.0005387018, 0.0005403389, 0.0005397233, 
    0.0005408532, 0.00054108, 0.0005393631, 0.0005404172, 0.000537033, 
    0.0005375797, 0.0005372542, 0.0005360644, 0.0005398645, 0.0005379145, 
    0.0005415145, 0.0005404587, 0.0005435391, 0.0005420073, 0.0005450154, 
    0.0005463004, 0.00054751, 0.0005489225, 0.0005369583, 0.0005365446, 
    0.0005372853, 0.0005383097, 0.0005392603, 0.0005405237, 0.0005406529, 
    0.0005408895, 0.0005415023, 0.0005420175, 0.000540964, 0.0005421465, 
    0.0005377062, 0.0005400337, 0.0005363874, 0.0005374855, 0.0005382486, 
    0.000537914, 0.0005396522, 0.0005400617, 0.0005417254, 0.0005408655, 
    0.000545983, 0.0005437196, 0.0005499979, 0.0005482442, 0.0005364, 
    0.0005369568, 0.0005388941, 0.0005379724, 0.0005406079, 0.0005412564, 
    0.0005417835, 0.0005424571, 0.0005425297, 0.0005429288, 0.0005422747, 
    0.000542903, 0.0005405258, 0.0005415882, 0.0005386722, 0.0005393819, 
    0.0005390554, 0.0005386971, 0.0005398026, 0.0005409799, 0.0005410052, 
    0.0005413825, 0.0005424455, 0.0005406176, 0.0005462745, 0.0005427814, 
    0.0005375638, 0.0005386358, 0.000538789, 0.0005383738, 0.0005411912, 
    0.0005401705, 0.0005429192, 0.0005421764, 0.0005433931, 0.0005427885, 
    0.0005426994, 0.0005419228, 0.000541439, 0.0005402169, 0.0005392222, 
    0.0005384334, 0.0005386167, 0.0005394831, 0.0005410518, 0.0005425356, 
    0.0005422105, 0.0005433, 0.0005404158, 0.0005416253, 0.0005411577, 
    0.0005423766, 0.0005397066, 0.0005419807, 0.000539125, 0.0005393754, 
    0.0005401501, 0.000541708, 0.0005420528, 0.0005424207, 0.0005421935, 
    0.0005410921, 0.0005409116, 0.0005401309, 0.0005399152, 0.0005393204, 
    0.0005388277, 0.0005392777, 0.0005397502, 0.0005410922, 0.0005423011, 
    0.0005436187, 0.0005439413, 0.0005454797, 0.000544227, 0.0005462936, 
    0.0005445362, 0.0005475781, 0.0005421126, 0.000544486, 0.0005401854, 
    0.0005406489, 0.000541487, 0.000543409, 0.0005423715, 0.0005435848, 
    0.0005409045, 0.000539513, 0.0005391531, 0.0005384812, 0.0005391683, 
    0.0005391124, 0.0005397699, 0.0005395585, 0.0005411366, 0.000540289, 
    0.0005426964, 0.0005435746, 0.0005460539, 0.0005475729, 0.000549119, 
    0.0005498012, 0.0005500088, 0.0005500956 ;

 SMINN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_PLANT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_SOIL1N_L1 =
  3.610095e-14, 3.619275e-14, 3.617492e-14, 3.624889e-14, 3.620788e-14, 
    3.625629e-14, 3.611958e-14, 3.619638e-14, 3.614737e-14, 3.610924e-14, 
    3.63922e-14, 3.625219e-14, 3.65375e-14, 3.644839e-14, 3.667211e-14, 
    3.652362e-14, 3.670202e-14, 3.666786e-14, 3.67707e-14, 3.674125e-14, 
    3.687256e-14, 3.678428e-14, 3.694059e-14, 3.68515e-14, 3.686543e-14, 
    3.678136e-14, 3.628042e-14, 3.637477e-14, 3.627482e-14, 3.628828e-14, 
    3.628225e-14, 3.620871e-14, 3.617161e-14, 3.609395e-14, 3.610806e-14, 
    3.616511e-14, 3.629434e-14, 3.625051e-14, 3.636097e-14, 3.635848e-14, 
    3.648126e-14, 3.642592e-14, 3.663201e-14, 3.65735e-14, 3.674248e-14, 
    3.670001e-14, 3.674048e-14, 3.672822e-14, 3.674064e-14, 3.667835e-14, 
    3.670504e-14, 3.665022e-14, 3.643628e-14, 3.649921e-14, 3.631136e-14, 
    3.619815e-14, 3.612295e-14, 3.606952e-14, 3.607707e-14, 3.609147e-14, 
    3.616544e-14, 3.623496e-14, 3.628789e-14, 3.632327e-14, 3.635812e-14, 
    3.646343e-14, 3.651919e-14, 3.664382e-14, 3.662137e-14, 3.665942e-14, 
    3.669579e-14, 3.675678e-14, 3.674675e-14, 3.67736e-14, 3.665844e-14, 
    3.673498e-14, 3.660857e-14, 3.664316e-14, 3.636748e-14, 3.626234e-14, 
    3.621752e-14, 3.617835e-14, 3.608288e-14, 3.614881e-14, 3.612282e-14, 
    3.618466e-14, 3.622391e-14, 3.620451e-14, 3.632424e-14, 3.627771e-14, 
    3.652249e-14, 3.641715e-14, 3.669155e-14, 3.662598e-14, 3.670726e-14, 
    3.66658e-14, 3.673682e-14, 3.667291e-14, 3.678359e-14, 3.680766e-14, 
    3.679121e-14, 3.685442e-14, 3.666936e-14, 3.674047e-14, 3.620396e-14, 
    3.620712e-14, 3.622187e-14, 3.615699e-14, 3.615303e-14, 3.609356e-14, 
    3.614649e-14, 3.616901e-14, 3.622619e-14, 3.625998e-14, 3.629209e-14, 
    3.636265e-14, 3.644136e-14, 3.655131e-14, 3.663023e-14, 3.668308e-14, 
    3.665069e-14, 3.667928e-14, 3.664731e-14, 3.663232e-14, 3.679864e-14, 
    3.670529e-14, 3.684533e-14, 3.683759e-14, 3.677423e-14, 3.683846e-14, 
    3.620934e-14, 3.619113e-14, 3.612782e-14, 3.617737e-14, 3.608708e-14, 
    3.613762e-14, 3.616665e-14, 3.627865e-14, 3.630327e-14, 3.632605e-14, 
    3.637105e-14, 3.642875e-14, 3.652987e-14, 3.661775e-14, 3.669791e-14, 
    3.669204e-14, 3.669411e-14, 3.671199e-14, 3.666767e-14, 3.671926e-14, 
    3.672791e-14, 3.670529e-14, 3.683655e-14, 3.679908e-14, 3.683743e-14, 
    3.681303e-14, 3.619705e-14, 3.62277e-14, 3.621114e-14, 3.624228e-14, 
    3.622033e-14, 3.631783e-14, 3.634704e-14, 3.64836e-14, 3.642761e-14, 
    3.651673e-14, 3.643668e-14, 3.645086e-14, 3.651959e-14, 3.644101e-14, 
    3.661289e-14, 3.649636e-14, 3.671268e-14, 3.659643e-14, 3.671996e-14, 
    3.669756e-14, 3.673466e-14, 3.676785e-14, 3.680961e-14, 3.688657e-14, 
    3.686876e-14, 3.693309e-14, 3.627339e-14, 3.63131e-14, 3.630962e-14, 
    3.635117e-14, 3.638188e-14, 3.644842e-14, 3.655501e-14, 3.651495e-14, 
    3.65885e-14, 3.660324e-14, 3.649152e-14, 3.656011e-14, 3.633967e-14, 
    3.637531e-14, 3.635411e-14, 3.627651e-14, 3.652416e-14, 3.639715e-14, 
    3.663153e-14, 3.656285e-14, 3.676312e-14, 3.666357e-14, 3.685895e-14, 
    3.694226e-14, 3.702068e-14, 3.71121e-14, 3.633478e-14, 3.630781e-14, 
    3.635611e-14, 3.642286e-14, 3.64848e-14, 3.656704e-14, 3.657546e-14, 
    3.659085e-14, 3.663072e-14, 3.666422e-14, 3.65957e-14, 3.667262e-14, 
    3.638353e-14, 3.653518e-14, 3.629759e-14, 3.636918e-14, 3.641894e-14, 
    3.639713e-14, 3.651038e-14, 3.653703e-14, 3.664526e-14, 3.658935e-14, 
    3.692169e-14, 3.677483e-14, 3.71817e-14, 3.706821e-14, 3.629837e-14, 
    3.633469e-14, 3.646094e-14, 3.640091e-14, 3.657254e-14, 3.661472e-14, 
    3.664901e-14, 3.669278e-14, 3.669752e-14, 3.672345e-14, 3.668096e-14, 
    3.672178e-14, 3.656722e-14, 3.663633e-14, 3.644655e-14, 3.649277e-14, 
    3.647152e-14, 3.644818e-14, 3.652018e-14, 3.659677e-14, 3.659844e-14, 
    3.662297e-14, 3.669201e-14, 3.657324e-14, 3.694056e-14, 3.671386e-14, 
    3.637428e-14, 3.644411e-14, 3.645412e-14, 3.642708e-14, 3.661049e-14, 
    3.654408e-14, 3.672282e-14, 3.667456e-14, 3.675363e-14, 3.671434e-14, 
    3.670856e-14, 3.665809e-14, 3.662663e-14, 3.654712e-14, 3.648237e-14, 
    3.6431e-14, 3.644295e-14, 3.649937e-14, 3.660146e-14, 3.669794e-14, 
    3.667681e-14, 3.674762e-14, 3.656011e-14, 3.663877e-14, 3.660837e-14, 
    3.668763e-14, 3.651388e-14, 3.666176e-14, 3.647602e-14, 3.649233e-14, 
    3.654276e-14, 3.664408e-14, 3.666653e-14, 3.669043e-14, 3.667569e-14, 
    3.660405e-14, 3.659233e-14, 3.654154e-14, 3.65275e-14, 3.648878e-14, 
    3.64567e-14, 3.648601e-14, 3.651676e-14, 3.66041e-14, 3.66827e-14, 
    3.676832e-14, 3.678927e-14, 3.688906e-14, 3.680779e-14, 3.694181e-14, 
    3.682781e-14, 3.702507e-14, 3.667037e-14, 3.682453e-14, 3.654506e-14, 
    3.657523e-14, 3.662972e-14, 3.675463e-14, 3.668726e-14, 3.676606e-14, 
    3.659187e-14, 3.65013e-14, 3.647789e-14, 3.643412e-14, 3.647889e-14, 
    3.647525e-14, 3.651806e-14, 3.650431e-14, 3.6607e-14, 3.655186e-14, 
    3.670841e-14, 3.676545e-14, 3.692634e-14, 3.702477e-14, 3.712488e-14, 
    3.716902e-14, 3.718245e-14, 3.718806e-14 ;

 SMINN_TO_SOIL1N_L2 =
  1.20043e-14, 1.203486e-14, 1.202892e-14, 1.205355e-14, 1.203989e-14, 
    1.205601e-14, 1.20105e-14, 1.203607e-14, 1.201975e-14, 1.200706e-14, 
    1.210125e-14, 1.205465e-14, 1.214962e-14, 1.211995e-14, 1.219443e-14, 
    1.2145e-14, 1.220438e-14, 1.219301e-14, 1.222724e-14, 1.221744e-14, 
    1.226115e-14, 1.223177e-14, 1.22838e-14, 1.225414e-14, 1.225878e-14, 
    1.223079e-14, 1.206404e-14, 1.209545e-14, 1.206218e-14, 1.206666e-14, 
    1.206465e-14, 1.204017e-14, 1.202782e-14, 1.200197e-14, 1.200667e-14, 
    1.202566e-14, 1.206867e-14, 1.205409e-14, 1.209086e-14, 1.209003e-14, 
    1.21309e-14, 1.211248e-14, 1.218108e-14, 1.21616e-14, 1.221785e-14, 
    1.220372e-14, 1.221719e-14, 1.22131e-14, 1.221724e-14, 1.21965e-14, 
    1.220539e-14, 1.218714e-14, 1.211592e-14, 1.213687e-14, 1.207434e-14, 
    1.203666e-14, 1.201162e-14, 1.199384e-14, 1.199635e-14, 1.200115e-14, 
    1.202577e-14, 1.204891e-14, 1.206653e-14, 1.207831e-14, 1.208991e-14, 
    1.212496e-14, 1.214352e-14, 1.218501e-14, 1.217754e-14, 1.21902e-14, 
    1.220231e-14, 1.222261e-14, 1.221927e-14, 1.222821e-14, 1.218987e-14, 
    1.221536e-14, 1.217328e-14, 1.218479e-14, 1.209302e-14, 1.205802e-14, 
    1.20431e-14, 1.203006e-14, 1.199829e-14, 1.202023e-14, 1.201158e-14, 
    1.203217e-14, 1.204523e-14, 1.203877e-14, 1.207863e-14, 1.206314e-14, 
    1.214462e-14, 1.210955e-14, 1.22009e-14, 1.217907e-14, 1.220613e-14, 
    1.219233e-14, 1.221597e-14, 1.219469e-14, 1.223154e-14, 1.223955e-14, 
    1.223407e-14, 1.225511e-14, 1.219351e-14, 1.221718e-14, 1.203859e-14, 
    1.203964e-14, 1.204455e-14, 1.202296e-14, 1.202164e-14, 1.200184e-14, 
    1.201946e-14, 1.202696e-14, 1.204599e-14, 1.205724e-14, 1.206793e-14, 
    1.209141e-14, 1.211761e-14, 1.215422e-14, 1.218049e-14, 1.219808e-14, 
    1.218729e-14, 1.219682e-14, 1.218617e-14, 1.218118e-14, 1.223655e-14, 
    1.220547e-14, 1.225209e-14, 1.224951e-14, 1.222842e-14, 1.22498e-14, 
    1.204038e-14, 1.203432e-14, 1.201324e-14, 1.202974e-14, 1.199969e-14, 
    1.201651e-14, 1.202617e-14, 1.206345e-14, 1.207165e-14, 1.207923e-14, 
    1.209421e-14, 1.211342e-14, 1.214708e-14, 1.217633e-14, 1.220301e-14, 
    1.220106e-14, 1.220175e-14, 1.22077e-14, 1.219295e-14, 1.221012e-14, 
    1.2213e-14, 1.220547e-14, 1.224917e-14, 1.223669e-14, 1.224946e-14, 
    1.224134e-14, 1.203629e-14, 1.204649e-14, 1.204098e-14, 1.205135e-14, 
    1.204404e-14, 1.20765e-14, 1.208622e-14, 1.213168e-14, 1.211304e-14, 
    1.21427e-14, 1.211606e-14, 1.212078e-14, 1.214366e-14, 1.21175e-14, 
    1.217471e-14, 1.213592e-14, 1.220793e-14, 1.216924e-14, 1.221036e-14, 
    1.22029e-14, 1.221525e-14, 1.22263e-14, 1.22402e-14, 1.226582e-14, 
    1.225989e-14, 1.22813e-14, 1.20617e-14, 1.207492e-14, 1.207376e-14, 
    1.208759e-14, 1.209781e-14, 1.211997e-14, 1.215545e-14, 1.214211e-14, 
    1.216659e-14, 1.21715e-14, 1.213431e-14, 1.215715e-14, 1.208377e-14, 
    1.209563e-14, 1.208857e-14, 1.206274e-14, 1.214518e-14, 1.21029e-14, 
    1.218092e-14, 1.215806e-14, 1.222472e-14, 1.219158e-14, 1.225662e-14, 
    1.228435e-14, 1.231046e-14, 1.234089e-14, 1.208214e-14, 1.207316e-14, 
    1.208924e-14, 1.211146e-14, 1.213208e-14, 1.215945e-14, 1.216225e-14, 
    1.216738e-14, 1.218065e-14, 1.21918e-14, 1.216899e-14, 1.21946e-14, 
    1.209836e-14, 1.214884e-14, 1.206976e-14, 1.209359e-14, 1.211015e-14, 
    1.210289e-14, 1.214059e-14, 1.214946e-14, 1.218549e-14, 1.216688e-14, 
    1.227751e-14, 1.222862e-14, 1.236406e-14, 1.232628e-14, 1.207002e-14, 
    1.208211e-14, 1.212413e-14, 1.210415e-14, 1.216128e-14, 1.217532e-14, 
    1.218674e-14, 1.220131e-14, 1.220289e-14, 1.221152e-14, 1.219737e-14, 
    1.221096e-14, 1.215951e-14, 1.218252e-14, 1.211934e-14, 1.213473e-14, 
    1.212765e-14, 1.211989e-14, 1.214385e-14, 1.216935e-14, 1.21699e-14, 
    1.217807e-14, 1.220105e-14, 1.216151e-14, 1.228379e-14, 1.220833e-14, 
    1.209529e-14, 1.211853e-14, 1.212186e-14, 1.211286e-14, 1.217391e-14, 
    1.215181e-14, 1.221131e-14, 1.219524e-14, 1.222156e-14, 1.220849e-14, 
    1.220656e-14, 1.218976e-14, 1.217929e-14, 1.215282e-14, 1.213127e-14, 
    1.211417e-14, 1.211815e-14, 1.213692e-14, 1.217091e-14, 1.220302e-14, 
    1.219599e-14, 1.221956e-14, 1.215714e-14, 1.218333e-14, 1.217321e-14, 
    1.219959e-14, 1.214175e-14, 1.219098e-14, 1.212915e-14, 1.213458e-14, 
    1.215137e-14, 1.21851e-14, 1.219257e-14, 1.220053e-14, 1.219562e-14, 
    1.217177e-14, 1.216787e-14, 1.215096e-14, 1.214629e-14, 1.21334e-14, 
    1.212272e-14, 1.213248e-14, 1.214271e-14, 1.217179e-14, 1.219795e-14, 
    1.222645e-14, 1.223343e-14, 1.226665e-14, 1.223959e-14, 1.228421e-14, 
    1.224626e-14, 1.231192e-14, 1.219385e-14, 1.224516e-14, 1.215214e-14, 
    1.216218e-14, 1.218032e-14, 1.22219e-14, 1.219947e-14, 1.22257e-14, 
    1.216772e-14, 1.213757e-14, 1.212977e-14, 1.211521e-14, 1.213011e-14, 
    1.21289e-14, 1.214315e-14, 1.213857e-14, 1.217275e-14, 1.21544e-14, 
    1.220651e-14, 1.22255e-14, 1.227905e-14, 1.231182e-14, 1.234515e-14, 
    1.235984e-14, 1.236431e-14, 1.236618e-14 ;

 SMINN_TO_SOIL1N_S2 =
  -1.00346e-10, -1.006209e-10, -1.005675e-10, -1.007892e-10, -1.006662e-10, 
    -1.008114e-10, -1.004018e-10, -1.006318e-10, -1.00485e-10, -1.003708e-10, 
    -1.012192e-10, -1.007991e-10, -1.016556e-10, -1.013878e-10, 
    -1.020605e-10, -1.016139e-10, -1.021505e-10, -1.020476e-10, 
    -1.023573e-10, -1.022686e-10, -1.026645e-10, -1.023983e-10, 
    -1.028698e-10, -1.02601e-10, -1.02643e-10, -1.023895e-10, -1.008837e-10, 
    -1.011669e-10, -1.008669e-10, -1.009073e-10, -1.008892e-10, 
    -1.006688e-10, -1.005577e-10, -1.00325e-10, -1.003673e-10, -1.005381e-10, 
    -1.009254e-10, -1.00794e-10, -1.011253e-10, -1.011178e-10, -1.014865e-10, 
    -1.013203e-10, -1.019397e-10, -1.017637e-10, -1.022723e-10, 
    -1.021444e-10, -1.022663e-10, -1.022294e-10, -1.022668e-10, 
    -1.020792e-10, -1.021596e-10, -1.019945e-10, -1.013514e-10, 
    -1.015404e-10, -1.009765e-10, -1.006372e-10, -1.004119e-10, 
    -1.002519e-10, -1.002745e-10, -1.003176e-10, -1.005391e-10, 
    -1.007474e-10, -1.009061e-10, -1.010122e-10, -1.011167e-10, -1.01433e-10, 
    -1.016005e-10, -1.019753e-10, -1.019077e-10, -1.020223e-10, 
    -1.021317e-10, -1.023154e-10, -1.022852e-10, -1.023661e-10, 
    -1.020193e-10, -1.022498e-10, -1.018692e-10, -1.019733e-10, -1.01145e-10, 
    -1.008295e-10, -1.006952e-10, -1.005778e-10, -1.002919e-10, 
    -1.004893e-10, -1.004115e-10, -1.005967e-10, -1.007143e-10, 
    -1.006561e-10, -1.010151e-10, -1.008755e-10, -1.016104e-10, -1.01294e-10, 
    -1.021189e-10, -1.019216e-10, -1.021662e-10, -1.020414e-10, 
    -1.022553e-10, -1.020628e-10, -1.023962e-10, -1.024688e-10, 
    -1.024192e-10, -1.026097e-10, -1.020521e-10, -1.022663e-10, 
    -1.006545e-10, -1.00664e-10, -1.007082e-10, -1.005138e-10, -1.00502e-10, 
    -1.003239e-10, -1.004824e-10, -1.005498e-10, -1.007211e-10, 
    -1.008224e-10, -1.009187e-10, -1.011303e-10, -1.013667e-10, 
    -1.016971e-10, -1.019344e-10, -1.020934e-10, -1.019959e-10, -1.02082e-10, 
    -1.019858e-10, -1.019407e-10, -1.024416e-10, -1.021603e-10, 
    -1.025823e-10, -1.02559e-10, -1.02368e-10, -1.025616e-10, -1.006706e-10, 
    -1.00616e-10, -1.004264e-10, -1.005748e-10, -1.003045e-10, -1.004558e-10, 
    -1.005428e-10, -1.008784e-10, -1.009522e-10, -1.010205e-10, 
    -1.011556e-10, -1.013288e-10, -1.016326e-10, -1.018969e-10, 
    -1.021381e-10, -1.021204e-10, -1.021266e-10, -1.021805e-10, 
    -1.020471e-10, -1.022024e-10, -1.022285e-10, -1.021603e-10, 
    -1.025559e-10, -1.024429e-10, -1.025585e-10, -1.024849e-10, 
    -1.006338e-10, -1.007257e-10, -1.00676e-10, -1.007693e-10, -1.007036e-10, 
    -1.009959e-10, -1.010836e-10, -1.014936e-10, -1.013254e-10, 
    -1.015931e-10, -1.013526e-10, -1.013952e-10, -1.016018e-10, 
    -1.013656e-10, -1.018823e-10, -1.01532e-10, -1.021826e-10, -1.018328e-10, 
    -1.022045e-10, -1.02137e-10, -1.022488e-10, -1.023488e-10, -1.024746e-10, 
    -1.027068e-10, -1.02653e-10, -1.028471e-10, -1.008626e-10, -1.009817e-10, 
    -1.009712e-10, -1.010959e-10, -1.011881e-10, -1.013878e-10, 
    -1.017081e-10, -1.015877e-10, -1.018088e-10, -1.018532e-10, 
    -1.015173e-10, -1.017235e-10, -1.010614e-10, -1.011684e-10, 
    -1.011047e-10, -1.00872e-10, -1.016154e-10, -1.012339e-10, -1.019383e-10, 
    -1.017317e-10, -1.023345e-10, -1.020348e-10, -1.026234e-10, 
    -1.028749e-10, -1.031117e-10, -1.033881e-10, -1.010467e-10, 
    -1.009658e-10, -1.011107e-10, -1.013111e-10, -1.014971e-10, 
    -1.017443e-10, -1.017696e-10, -1.018159e-10, -1.019359e-10, 
    -1.020367e-10, -1.018305e-10, -1.020619e-10, -1.011932e-10, 
    -1.016486e-10, -1.009352e-10, -1.0115e-10, -1.012993e-10, -1.012339e-10, 
    -1.01574e-10, -1.016541e-10, -1.019796e-10, -1.018114e-10, -1.028128e-10, 
    -1.023699e-10, -1.035986e-10, -1.032554e-10, -1.009375e-10, 
    -1.010465e-10, -1.014255e-10, -1.012452e-10, -1.017608e-10, 
    -1.018877e-10, -1.019909e-10, -1.021227e-10, -1.021369e-10, -1.02215e-10, 
    -1.020871e-10, -1.0221e-10, -1.017449e-10, -1.019527e-10, -1.013822e-10, 
    -1.015211e-10, -1.014572e-10, -1.013871e-10, -1.016034e-10, 
    -1.018338e-10, -1.018387e-10, -1.019126e-10, -1.021206e-10, 
    -1.017629e-10, -1.028699e-10, -1.021863e-10, -1.011652e-10, -1.01375e-10, 
    -1.01405e-10, -1.013237e-10, -1.01875e-10, -1.016753e-10, -1.022131e-10, 
    -1.020678e-10, -1.023059e-10, -1.021876e-10, -1.021702e-10, 
    -1.020182e-10, -1.019236e-10, -1.016844e-10, -1.014898e-10, 
    -1.013355e-10, -1.013714e-10, -1.015409e-10, -1.018479e-10, 
    -1.021382e-10, -1.020746e-10, -1.022878e-10, -1.017235e-10, 
    -1.019601e-10, -1.018686e-10, -1.021072e-10, -1.015845e-10, 
    -1.020295e-10, -1.014707e-10, -1.015197e-10, -1.016713e-10, 
    -1.019761e-10, -1.020436e-10, -1.021156e-10, -1.020712e-10, 
    -1.018557e-10, -1.018204e-10, -1.016676e-10, -1.016255e-10, 
    -1.015091e-10, -1.014127e-10, -1.015007e-10, -1.015932e-10, 
    -1.018558e-10, -1.020923e-10, -1.023502e-10, -1.024133e-10, 
    -1.027144e-10, -1.024692e-10, -1.028737e-10, -1.025298e-10, 
    -1.031251e-10, -1.020553e-10, -1.025197e-10, -1.016782e-10, 
    -1.017689e-10, -1.019329e-10, -1.02309e-10, -1.02106e-10, -1.023434e-10, 
    -1.01819e-10, -1.015467e-10, -1.014763e-10, -1.013449e-10, -1.014793e-10, 
    -1.014684e-10, -1.015971e-10, -1.015557e-10, -1.018645e-10, 
    -1.016986e-10, -1.021697e-10, -1.023416e-10, -1.028268e-10, 
    -1.031241e-10, -1.034267e-10, -1.035602e-10, -1.036009e-10, -1.036179e-10 ;

 SMINN_TO_SOIL1N_S3 =
  -2.418412e-12, -2.425036e-12, -2.423749e-12, -2.42909e-12, -2.426127e-12, 
    -2.429624e-12, -2.419756e-12, -2.425298e-12, -2.42176e-12, -2.419009e-12, 
    -2.43945e-12, -2.429328e-12, -2.449965e-12, -2.443512e-12, -2.45972e-12, 
    -2.44896e-12, -2.46189e-12, -2.459411e-12, -2.466873e-12, -2.464735e-12, 
    -2.474275e-12, -2.467859e-12, -2.47922e-12, -2.472743e-12, -2.473756e-12, 
    -2.467647e-12, -2.431367e-12, -2.43819e-12, -2.430962e-12, -2.431935e-12, 
    -2.431499e-12, -2.426188e-12, -2.423511e-12, -2.417906e-12, 
    -2.418924e-12, -2.423041e-12, -2.432373e-12, -2.429206e-12, 
    -2.437188e-12, -2.437008e-12, -2.44589e-12, -2.441886e-12, -2.456811e-12, 
    -2.452571e-12, -2.464825e-12, -2.461743e-12, -2.46468e-12, -2.46379e-12, 
    -2.464691e-12, -2.460172e-12, -2.462108e-12, -2.458132e-12, 
    -2.442636e-12, -2.44719e-12, -2.433603e-12, -2.425427e-12, -2.419998e-12, 
    -2.416145e-12, -2.416689e-12, -2.417728e-12, -2.423065e-12, 
    -2.428083e-12, -2.431906e-12, -2.434463e-12, -2.436982e-12, 
    -2.444603e-12, -2.448638e-12, -2.457668e-12, -2.45604e-12, -2.458799e-12, 
    -2.461437e-12, -2.465863e-12, -2.465134e-12, -2.467084e-12, 
    -2.458727e-12, -2.464281e-12, -2.455112e-12, -2.45762e-12, -2.437663e-12, 
    -2.430061e-12, -2.426825e-12, -2.423996e-12, -2.417108e-12, 
    -2.421865e-12, -2.41999e-12, -2.424451e-12, -2.427285e-12, -2.425883e-12, 
    -2.434533e-12, -2.43117e-12, -2.448877e-12, -2.441252e-12, -2.461129e-12, 
    -2.456374e-12, -2.462269e-12, -2.459261e-12, -2.464414e-12, 
    -2.459777e-12, -2.46781e-12, -2.469558e-12, -2.468363e-12, -2.472954e-12, 
    -2.45952e-12, -2.464679e-12, -2.425844e-12, -2.426073e-12, -2.427138e-12, 
    -2.422455e-12, -2.422169e-12, -2.417878e-12, -2.421697e-12, 
    -2.423322e-12, -2.42745e-12, -2.42989e-12, -2.43221e-12, -2.437309e-12, 
    -2.443003e-12, -2.450964e-12, -2.456682e-12, -2.460515e-12, 
    -2.458165e-12, -2.460239e-12, -2.45792e-12, -2.456834e-12, -2.468903e-12, 
    -2.462126e-12, -2.472294e-12, -2.471732e-12, -2.46713e-12, -2.471795e-12, 
    -2.426233e-12, -2.424918e-12, -2.42035e-12, -2.423925e-12, -2.417411e-12, 
    -2.421057e-12, -2.423153e-12, -2.43124e-12, -2.433017e-12, -2.434664e-12, 
    -2.437917e-12, -2.442091e-12, -2.449411e-12, -2.455778e-12, -2.46159e-12, 
    -2.461165e-12, -2.461315e-12, -2.462612e-12, -2.459397e-12, -2.46314e-12, 
    -2.463768e-12, -2.462126e-12, -2.471656e-12, -2.468934e-12, -2.47172e-12, 
    -2.469947e-12, -2.425346e-12, -2.427559e-12, -2.426363e-12, 
    -2.428612e-12, -2.427027e-12, -2.434071e-12, -2.436183e-12, 
    -2.446061e-12, -2.442008e-12, -2.448459e-12, -2.442664e-12, 
    -2.443691e-12, -2.448668e-12, -2.442978e-12, -2.455426e-12, 
    -2.446986e-12, -2.462663e-12, -2.454235e-12, -2.463191e-12, 
    -2.461565e-12, -2.464257e-12, -2.466667e-12, -2.469699e-12, 
    -2.475292e-12, -2.473997e-12, -2.478674e-12, -2.430858e-12, 
    -2.433728e-12, -2.433476e-12, -2.436479e-12, -2.4387e-12, -2.443514e-12, 
    -2.451231e-12, -2.44833e-12, -2.453657e-12, -2.454726e-12, -2.446633e-12, 
    -2.451602e-12, -2.435649e-12, -2.438226e-12, -2.436692e-12, 
    -2.431084e-12, -2.448997e-12, -2.439806e-12, -2.456777e-12, -2.4518e-12, 
    -2.466323e-12, -2.459101e-12, -2.473284e-12, -2.479343e-12, 
    -2.485047e-12, -2.491708e-12, -2.435295e-12, -2.433345e-12, 
    -2.436837e-12, -2.441666e-12, -2.446147e-12, -2.452103e-12, 
    -2.452713e-12, -2.453828e-12, -2.456718e-12, -2.459147e-12, -2.45418e-12, 
    -2.459755e-12, -2.438823e-12, -2.449795e-12, -2.432607e-12, 
    -2.437783e-12, -2.441381e-12, -2.439804e-12, -2.447998e-12, 
    -2.449929e-12, -2.457773e-12, -2.453719e-12, -2.477847e-12, 
    -2.467175e-12, -2.496781e-12, -2.48851e-12, -2.432663e-12, -2.435288e-12, 
    -2.444421e-12, -2.440076e-12, -2.452501e-12, -2.455558e-12, 
    -2.458043e-12, -2.461219e-12, -2.461562e-12, -2.463444e-12, 
    -2.460361e-12, -2.463322e-12, -2.452116e-12, -2.457124e-12, 
    -2.443378e-12, -2.446724e-12, -2.445185e-12, -2.443496e-12, 
    -2.448708e-12, -2.454258e-12, -2.454378e-12, -2.456157e-12, 
    -2.461168e-12, -2.452551e-12, -2.479222e-12, -2.462753e-12, -2.43815e-12, 
    -2.443203e-12, -2.443927e-12, -2.441969e-12, -2.455251e-12, 
    -2.450439e-12, -2.463398e-12, -2.459897e-12, -2.465634e-12, 
    -2.462783e-12, -2.462364e-12, -2.458702e-12, -2.456422e-12, -2.45066e-12, 
    -2.445971e-12, -2.442253e-12, -2.443118e-12, -2.447202e-12, 
    -2.454598e-12, -2.461593e-12, -2.460061e-12, -2.465198e-12, -2.4516e-12, 
    -2.457302e-12, -2.455098e-12, -2.460845e-12, -2.448252e-12, 
    -2.458973e-12, -2.445511e-12, -2.446692e-12, -2.450344e-12, 
    -2.457688e-12, -2.459314e-12, -2.461049e-12, -2.459979e-12, 
    -2.454786e-12, -2.453935e-12, -2.450255e-12, -2.449239e-12, 
    -2.446435e-12, -2.444112e-12, -2.446234e-12, -2.448462e-12, 
    -2.454788e-12, -2.460488e-12, -2.466701e-12, -2.468222e-12, 
    -2.475476e-12, -2.469569e-12, -2.479314e-12, -2.471027e-12, 
    -2.485371e-12, -2.459596e-12, -2.470785e-12, -2.45051e-12, -2.452696e-12, 
    -2.456647e-12, -2.465709e-12, -2.460818e-12, -2.466538e-12, 
    -2.453902e-12, -2.447342e-12, -2.445646e-12, -2.442479e-12, 
    -2.445719e-12, -2.445455e-12, -2.448554e-12, -2.447559e-12, 
    -2.454998e-12, -2.451003e-12, -2.462353e-12, -2.466493e-12, 
    -2.478184e-12, -2.485347e-12, -2.492638e-12, -2.495856e-12, 
    -2.496835e-12, -2.497244e-12 ;

 SMINN_TO_SOIL2N_L3 =
  3.899645e-15, 3.909572e-15, 3.907644e-15, 3.915643e-15, 3.911208e-15, 
    3.916443e-15, 3.90166e-15, 3.909965e-15, 3.904665e-15, 3.900542e-15, 
    3.931139e-15, 3.916e-15, 3.946852e-15, 3.937215e-15, 3.961407e-15, 
    3.945351e-15, 3.964642e-15, 3.960948e-15, 3.972069e-15, 3.968885e-15, 
    3.983084e-15, 3.973538e-15, 3.990441e-15, 3.980808e-15, 3.982314e-15, 
    3.973222e-15, 3.919052e-15, 3.929255e-15, 3.918446e-15, 3.919902e-15, 
    3.91925e-15, 3.911298e-15, 3.907286e-15, 3.898888e-15, 3.900414e-15, 
    3.906583e-15, 3.920557e-15, 3.915818e-15, 3.927763e-15, 3.927494e-15, 
    3.94077e-15, 3.934786e-15, 3.957072e-15, 3.950745e-15, 3.969018e-15, 
    3.964425e-15, 3.968802e-15, 3.967475e-15, 3.968819e-15, 3.962083e-15, 
    3.964969e-15, 3.959041e-15, 3.935906e-15, 3.942711e-15, 3.922398e-15, 
    3.910156e-15, 3.902024e-15, 3.896247e-15, 3.897063e-15, 3.89862e-15, 
    3.906619e-15, 3.914137e-15, 3.91986e-15, 3.923686e-15, 3.927455e-15, 
    3.938843e-15, 3.944871e-15, 3.958349e-15, 3.955921e-15, 3.960036e-15, 
    3.963969e-15, 3.970564e-15, 3.969479e-15, 3.972383e-15, 3.959929e-15, 
    3.968207e-15, 3.954537e-15, 3.958278e-15, 3.928467e-15, 3.917098e-15, 
    3.91225e-15, 3.908014e-15, 3.897691e-15, 3.904821e-15, 3.902011e-15, 
    3.908697e-15, 3.912942e-15, 3.910843e-15, 3.923791e-15, 3.918759e-15, 
    3.945228e-15, 3.933837e-15, 3.96351e-15, 3.95642e-15, 3.965209e-15, 
    3.960726e-15, 3.968405e-15, 3.961494e-15, 3.973464e-15, 3.976067e-15, 
    3.974288e-15, 3.981123e-15, 3.961111e-15, 3.9688e-15, 3.910784e-15, 
    3.911126e-15, 3.912721e-15, 3.905706e-15, 3.905277e-15, 3.898846e-15, 
    3.904569e-15, 3.907005e-15, 3.913188e-15, 3.916842e-15, 3.920314e-15, 
    3.927944e-15, 3.936455e-15, 3.948345e-15, 3.956879e-15, 3.962594e-15, 
    3.959091e-15, 3.962184e-15, 3.958726e-15, 3.957105e-15, 3.97509e-15, 
    3.964996e-15, 3.98014e-15, 3.979303e-15, 3.972451e-15, 3.979397e-15, 
    3.911366e-15, 3.909397e-15, 3.90255e-15, 3.907908e-15, 3.898146e-15, 
    3.90361e-15, 3.90675e-15, 3.918861e-15, 3.921523e-15, 3.923986e-15, 
    3.928853e-15, 3.935092e-15, 3.946026e-15, 3.95553e-15, 3.964198e-15, 
    3.963564e-15, 3.963787e-15, 3.965721e-15, 3.960928e-15, 3.966507e-15, 
    3.967442e-15, 3.964996e-15, 3.979191e-15, 3.975138e-15, 3.979285e-15, 
    3.976647e-15, 3.910037e-15, 3.913352e-15, 3.911561e-15, 3.914928e-15, 
    3.912555e-15, 3.923098e-15, 3.926256e-15, 3.941023e-15, 3.934969e-15, 
    3.944606e-15, 3.935949e-15, 3.937483e-15, 3.944915e-15, 3.936418e-15, 
    3.955004e-15, 3.942403e-15, 3.965796e-15, 3.953224e-15, 3.966583e-15, 
    3.964161e-15, 3.968172e-15, 3.971761e-15, 3.976277e-15, 3.984599e-15, 
    3.982674e-15, 3.98963e-15, 3.918292e-15, 3.922585e-15, 3.92221e-15, 
    3.926702e-15, 3.930023e-15, 3.937219e-15, 3.948745e-15, 3.944413e-15, 
    3.952366e-15, 3.953961e-15, 3.94188e-15, 3.949297e-15, 3.925459e-15, 
    3.929313e-15, 3.927021e-15, 3.918629e-15, 3.945409e-15, 3.931675e-15, 
    3.95702e-15, 3.949594e-15, 3.971249e-15, 3.960484e-15, 3.981613e-15, 
    3.990622e-15, 3.999102e-15, 4.008988e-15, 3.92493e-15, 3.922014e-15, 
    3.927237e-15, 3.934455e-15, 3.941153e-15, 3.950046e-15, 3.950957e-15, 
    3.952621e-15, 3.956933e-15, 3.960555e-15, 3.953145e-15, 3.961463e-15, 
    3.930202e-15, 3.946601e-15, 3.920909e-15, 3.92865e-15, 3.934031e-15, 
    3.931673e-15, 3.943919e-15, 3.946801e-15, 3.958505e-15, 3.952458e-15, 
    3.988397e-15, 3.972516e-15, 4.016515e-15, 4.004242e-15, 3.920994e-15, 
    3.924922e-15, 3.938573e-15, 3.932081e-15, 3.950641e-15, 3.955202e-15, 
    3.95891e-15, 3.963644e-15, 3.964156e-15, 3.96696e-15, 3.962365e-15, 
    3.966779e-15, 3.950065e-15, 3.957539e-15, 3.937017e-15, 3.942015e-15, 
    3.939717e-15, 3.937193e-15, 3.944978e-15, 3.953261e-15, 3.953442e-15, 
    3.956095e-15, 3.96356e-15, 3.950716e-15, 3.990437e-15, 3.965923e-15, 
    3.929202e-15, 3.936753e-15, 3.937836e-15, 3.934911e-15, 3.954745e-15, 
    3.947563e-15, 3.966892e-15, 3.961673e-15, 3.970223e-15, 3.965976e-15, 
    3.96535e-15, 3.959892e-15, 3.95649e-15, 3.947892e-15, 3.94089e-15, 
    3.935335e-15, 3.936628e-15, 3.942728e-15, 3.953768e-15, 3.964201e-15, 
    3.961916e-15, 3.969574e-15, 3.949296e-15, 3.957803e-15, 3.954515e-15, 
    3.963087e-15, 3.944297e-15, 3.960289e-15, 3.940204e-15, 3.941967e-15, 
    3.94742e-15, 3.958377e-15, 3.960805e-15, 3.96339e-15, 3.961795e-15, 
    3.954049e-15, 3.95278e-15, 3.947289e-15, 3.94577e-15, 3.941584e-15, 
    3.938114e-15, 3.941283e-15, 3.944609e-15, 3.954054e-15, 3.962554e-15, 
    3.971812e-15, 3.974077e-15, 3.984869e-15, 3.97608e-15, 3.990573e-15, 
    3.978246e-15, 3.999577e-15, 3.96122e-15, 3.97789e-15, 3.94767e-15, 
    3.950932e-15, 3.956825e-15, 3.970332e-15, 3.963047e-15, 3.971568e-15, 
    3.952731e-15, 3.942937e-15, 3.940405e-15, 3.935673e-15, 3.940513e-15, 
    3.94012e-15, 3.944749e-15, 3.943262e-15, 3.954367e-15, 3.948404e-15, 
    3.965333e-15, 3.971502e-15, 3.9889e-15, 3.999544e-15, 4.010371e-15, 
    4.015143e-15, 4.016596e-15, 4.017203e-15 ;

 SMINN_TO_SOIL2N_S1 =
  -1.050341e-08, -1.053215e-08, -1.052657e-08, -1.054975e-08, -1.053689e-08, 
    -1.055207e-08, -1.050924e-08, -1.053329e-08, -1.051794e-08, -1.0506e-08, 
    -1.059471e-08, -1.055078e-08, -1.064034e-08, -1.061234e-08, 
    -1.068268e-08, -1.063598e-08, -1.06921e-08, -1.068134e-08, -1.071372e-08, 
    -1.070445e-08, -1.074585e-08, -1.0718e-08, -1.076731e-08, -1.07392e-08, 
    -1.07436e-08, -1.071708e-08, -1.055963e-08, -1.058924e-08, -1.055787e-08, 
    -1.056209e-08, -1.05602e-08, -1.053715e-08, -1.052553e-08, -1.050121e-08, 
    -1.050563e-08, -1.052349e-08, -1.056399e-08, -1.055025e-08, 
    -1.058489e-08, -1.058411e-08, -1.062266e-08, -1.060528e-08, 
    -1.067006e-08, -1.065165e-08, -1.070483e-08, -1.069146e-08, 
    -1.070421e-08, -1.070034e-08, -1.070426e-08, -1.068464e-08, 
    -1.069305e-08, -1.067579e-08, -1.060853e-08, -1.06283e-08, -1.056933e-08, 
    -1.053385e-08, -1.051029e-08, -1.049356e-08, -1.049593e-08, 
    -1.050044e-08, -1.05236e-08, -1.054538e-08, -1.056197e-08, -1.057306e-08, 
    -1.0584e-08, -1.061707e-08, -1.063458e-08, -1.067378e-08, -1.066671e-08, 
    -1.067869e-08, -1.069013e-08, -1.070934e-08, -1.070618e-08, 
    -1.071464e-08, -1.067837e-08, -1.070248e-08, -1.066268e-08, 
    -1.067357e-08, -1.058695e-08, -1.055396e-08, -1.053992e-08, 
    -1.052764e-08, -1.049775e-08, -1.051839e-08, -1.051025e-08, 
    -1.052961e-08, -1.054191e-08, -1.053583e-08, -1.057337e-08, 
    -1.055878e-08, -1.063562e-08, -1.060253e-08, -1.06888e-08, -1.066816e-08, 
    -1.069374e-08, -1.068069e-08, -1.070305e-08, -1.068293e-08, 
    -1.071779e-08, -1.072538e-08, -1.072019e-08, -1.074012e-08, 
    -1.068181e-08, -1.07042e-08, -1.053566e-08, -1.053665e-08, -1.054127e-08, 
    -1.052095e-08, -1.051971e-08, -1.050109e-08, -1.051766e-08, 
    -1.052471e-08, -1.054263e-08, -1.055322e-08, -1.056329e-08, 
    -1.058542e-08, -1.061013e-08, -1.064468e-08, -1.06695e-08, -1.068613e-08, 
    -1.067593e-08, -1.068493e-08, -1.067487e-08, -1.067015e-08, 
    -1.072253e-08, -1.069312e-08, -1.073725e-08, -1.073481e-08, 
    -1.071484e-08, -1.073508e-08, -1.053735e-08, -1.053164e-08, 
    -1.051181e-08, -1.052733e-08, -1.049906e-08, -1.051488e-08, 
    -1.052398e-08, -1.055908e-08, -1.056679e-08, -1.057394e-08, 
    -1.058806e-08, -1.060617e-08, -1.063794e-08, -1.066557e-08, -1.06908e-08, 
    -1.068895e-08, -1.06896e-08, -1.069523e-08, -1.068128e-08, -1.069752e-08, 
    -1.070025e-08, -1.069312e-08, -1.073448e-08, -1.072267e-08, 
    -1.073476e-08, -1.072707e-08, -1.05335e-08, -1.05431e-08, -1.053791e-08, 
    -1.054767e-08, -1.054079e-08, -1.057136e-08, -1.058053e-08, -1.06234e-08, 
    -1.060581e-08, -1.063381e-08, -1.060866e-08, -1.061311e-08, 
    -1.063472e-08, -1.061002e-08, -1.066405e-08, -1.062742e-08, 
    -1.069545e-08, -1.065888e-08, -1.069774e-08, -1.069069e-08, 
    -1.070237e-08, -1.071283e-08, -1.072599e-08, -1.075026e-08, 
    -1.074464e-08, -1.076494e-08, -1.055742e-08, -1.056988e-08, 
    -1.056878e-08, -1.058182e-08, -1.059145e-08, -1.061235e-08, 
    -1.064584e-08, -1.063325e-08, -1.065637e-08, -1.066101e-08, 
    -1.062588e-08, -1.064745e-08, -1.057821e-08, -1.05894e-08, -1.058274e-08, 
    -1.05584e-08, -1.063614e-08, -1.059625e-08, -1.066991e-08, -1.064831e-08, 
    -1.071134e-08, -1.067999e-08, -1.074155e-08, -1.076784e-08, -1.07926e-08, 
    -1.082151e-08, -1.057668e-08, -1.056821e-08, -1.058337e-08, 
    -1.060432e-08, -1.062378e-08, -1.064962e-08, -1.065227e-08, 
    -1.065711e-08, -1.066965e-08, -1.068019e-08, -1.065864e-08, 
    -1.068283e-08, -1.059199e-08, -1.063961e-08, -1.056501e-08, 
    -1.058747e-08, -1.060309e-08, -1.059624e-08, -1.063181e-08, 
    -1.064019e-08, -1.067423e-08, -1.065663e-08, -1.076135e-08, 
    -1.071503e-08, -1.084352e-08, -1.080763e-08, -1.056526e-08, 
    -1.057665e-08, -1.061628e-08, -1.059743e-08, -1.065135e-08, 
    -1.066462e-08, -1.06754e-08, -1.068919e-08, -1.069068e-08, -1.069884e-08, 
    -1.068546e-08, -1.069831e-08, -1.064968e-08, -1.067142e-08, 
    -1.061176e-08, -1.062628e-08, -1.06196e-08, -1.061227e-08, -1.063489e-08, 
    -1.065898e-08, -1.065949e-08, -1.066722e-08, -1.068896e-08, 
    -1.065157e-08, -1.076732e-08, -1.069584e-08, -1.058907e-08, -1.0611e-08, 
    -1.061414e-08, -1.060564e-08, -1.066329e-08, -1.06424e-08, -1.069864e-08, 
    -1.068345e-08, -1.070835e-08, -1.069597e-08, -1.069415e-08, 
    -1.067826e-08, -1.066836e-08, -1.064336e-08, -1.062301e-08, 
    -1.060687e-08, -1.061063e-08, -1.062835e-08, -1.066045e-08, 
    -1.069081e-08, -1.068416e-08, -1.070645e-08, -1.064744e-08, 
    -1.067219e-08, -1.066262e-08, -1.068756e-08, -1.063291e-08, 
    -1.067944e-08, -1.062101e-08, -1.062614e-08, -1.064199e-08, 
    -1.067386e-08, -1.068092e-08, -1.068845e-08, -1.06838e-08, -1.066127e-08, 
    -1.065757e-08, -1.06416e-08, -1.063719e-08, -1.062502e-08, -1.061494e-08, 
    -1.062415e-08, -1.063382e-08, -1.066128e-08, -1.068601e-08, 
    -1.071298e-08, -1.071958e-08, -1.075106e-08, -1.072543e-08, 
    -1.076772e-08, -1.073175e-08, -1.0794e-08, -1.068214e-08, -1.07307e-08, 
    -1.064271e-08, -1.06522e-08, -1.066934e-08, -1.070867e-08, -1.068745e-08, 
    -1.071227e-08, -1.065743e-08, -1.062896e-08, -1.06216e-08, -1.060785e-08, 
    -1.062191e-08, -1.062077e-08, -1.063422e-08, -1.06299e-08, -1.066219e-08, 
    -1.064485e-08, -1.069411e-08, -1.071208e-08, -1.076281e-08, -1.07939e-08, 
    -1.082554e-08, -1.083951e-08, -1.084376e-08, -1.084553e-08 ;

 SMINN_TO_SOIL3N_S1 =
  -1.246224e-10, -1.249636e-10, -1.248973e-10, -1.251724e-10, -1.250198e-10, 
    -1.252e-10, -1.246916e-10, -1.249771e-10, -1.247948e-10, -1.246531e-10, 
    -1.257062e-10, -1.251847e-10, -1.262479e-10, -1.259154e-10, 
    -1.267505e-10, -1.261962e-10, -1.268623e-10, -1.267346e-10, -1.27119e-10, 
    -1.270089e-10, -1.275004e-10, -1.271698e-10, -1.277552e-10, 
    -1.274215e-10, -1.274736e-10, -1.271589e-10, -1.252897e-10, 
    -1.256413e-10, -1.252689e-10, -1.25319e-10, -1.252965e-10, -1.25023e-10, 
    -1.24885e-10, -1.245963e-10, -1.246487e-10, -1.248608e-10, -1.253416e-10, 
    -1.251784e-10, -1.255896e-10, -1.255804e-10, -1.26038e-10, -1.258317e-10, 
    -1.266006e-10, -1.263822e-10, -1.270135e-10, -1.268547e-10, -1.27006e-10, 
    -1.269602e-10, -1.270066e-10, -1.267738e-10, -1.268735e-10, 
    -1.266687e-10, -1.258703e-10, -1.26105e-10, -1.254049e-10, -1.249838e-10, 
    -1.247041e-10, -1.245055e-10, -1.245336e-10, -1.245871e-10, 
    -1.248621e-10, -1.251206e-10, -1.253175e-10, -1.254492e-10, -1.25579e-10, 
    -1.259717e-10, -1.261795e-10, -1.266448e-10, -1.265609e-10, 
    -1.267031e-10, -1.268389e-10, -1.27067e-10, -1.270294e-10, -1.271299e-10, 
    -1.266993e-10, -1.269855e-10, -1.265131e-10, -1.266423e-10, 
    -1.256141e-10, -1.252225e-10, -1.250558e-10, -1.2491e-10, -1.245552e-10, 
    -1.248002e-10, -1.247036e-10, -1.249335e-10, -1.250795e-10, 
    -1.250073e-10, -1.254528e-10, -1.252796e-10, -1.261919e-10, -1.25799e-10, 
    -1.268231e-10, -1.265781e-10, -1.268818e-10, -1.267269e-10, 
    -1.269923e-10, -1.267534e-10, -1.271673e-10, -1.272574e-10, 
    -1.271958e-10, -1.274323e-10, -1.267402e-10, -1.27006e-10, -1.250052e-10, 
    -1.25017e-10, -1.250719e-10, -1.248306e-10, -1.248159e-10, -1.245948e-10, 
    -1.247916e-10, -1.248753e-10, -1.250879e-10, -1.252137e-10, 
    -1.253332e-10, -1.255959e-10, -1.258893e-10, -1.262994e-10, -1.26594e-10, 
    -1.267914e-10, -1.266704e-10, -1.267772e-10, -1.266578e-10, 
    -1.266018e-10, -1.272236e-10, -1.268745e-10, -1.273983e-10, 
    -1.273693e-10, -1.271323e-10, -1.273726e-10, -1.250253e-10, 
    -1.249575e-10, -1.247222e-10, -1.249063e-10, -1.245708e-10, 
    -1.247586e-10, -1.248666e-10, -1.252832e-10, -1.253748e-10, 
    -1.254596e-10, -1.256272e-10, -1.258422e-10, -1.262194e-10, 
    -1.265474e-10, -1.268469e-10, -1.268249e-10, -1.268326e-10, 
    -1.268995e-10, -1.267338e-10, -1.269267e-10, -1.26959e-10, -1.268744e-10, 
    -1.273655e-10, -1.272252e-10, -1.273687e-10, -1.272774e-10, 
    -1.249795e-10, -1.250936e-10, -1.25032e-10, -1.251478e-10, -1.250662e-10, 
    -1.254291e-10, -1.255379e-10, -1.260468e-10, -1.25838e-10, -1.261704e-10, 
    -1.258718e-10, -1.259247e-10, -1.261811e-10, -1.258879e-10, 
    -1.265293e-10, -1.260944e-10, -1.269021e-10, -1.264679e-10, 
    -1.269293e-10, -1.268456e-10, -1.269842e-10, -1.271084e-10, 
    -1.272646e-10, -1.275528e-10, -1.27486e-10, -1.27727e-10, -1.252635e-10, 
    -1.254114e-10, -1.253984e-10, -1.255531e-10, -1.256675e-10, 
    -1.259155e-10, -1.263131e-10, -1.261637e-10, -1.264381e-10, 
    -1.264932e-10, -1.260762e-10, -1.263322e-10, -1.255104e-10, 
    -1.256431e-10, -1.255641e-10, -1.252752e-10, -1.261981e-10, 
    -1.257245e-10, -1.265989e-10, -1.263424e-10, -1.270907e-10, 
    -1.267186e-10, -1.274493e-10, -1.277615e-10, -1.280554e-10, 
    -1.283986e-10, -1.254921e-10, -1.253917e-10, -1.255716e-10, 
    -1.258203e-10, -1.260512e-10, -1.263581e-10, -1.263895e-10, 
    -1.264469e-10, -1.265958e-10, -1.26721e-10, -1.264651e-10, -1.267523e-10, 
    -1.256739e-10, -1.262392e-10, -1.253537e-10, -1.256203e-10, 
    -1.258057e-10, -1.257244e-10, -1.261466e-10, -1.26246e-10, -1.266502e-10, 
    -1.264413e-10, -1.276844e-10, -1.271346e-10, -1.286599e-10, 
    -1.282338e-10, -1.253566e-10, -1.254918e-10, -1.259623e-10, 
    -1.257384e-10, -1.263786e-10, -1.265361e-10, -1.266641e-10, 
    -1.268277e-10, -1.268454e-10, -1.269423e-10, -1.267835e-10, 
    -1.269361e-10, -1.263587e-10, -1.266168e-10, -1.259085e-10, 
    -1.260809e-10, -1.260017e-10, -1.259146e-10, -1.261831e-10, 
    -1.264691e-10, -1.264752e-10, -1.265669e-10, -1.268251e-10, 
    -1.263812e-10, -1.277553e-10, -1.269067e-10, -1.256392e-10, 
    -1.258996e-10, -1.259368e-10, -1.25836e-10, -1.265203e-10, -1.262724e-10, 
    -1.2694e-10, -1.267596e-10, -1.270552e-10, -1.269083e-10, -1.268867e-10, 
    -1.26698e-10, -1.265806e-10, -1.262837e-10, -1.260421e-10, -1.258506e-10, 
    -1.258951e-10, -1.261056e-10, -1.264866e-10, -1.26847e-10, -1.26768e-10, 
    -1.270327e-10, -1.263322e-10, -1.266259e-10, -1.265124e-10, 
    -1.268085e-10, -1.261597e-10, -1.26712e-10, -1.260184e-10, -1.260793e-10, 
    -1.262674e-10, -1.266458e-10, -1.267296e-10, -1.268189e-10, 
    -1.267638e-10, -1.264963e-10, -1.264525e-10, -1.262629e-10, 
    -1.262105e-10, -1.26066e-10, -1.259464e-10, -1.260557e-10, -1.261704e-10, 
    -1.264964e-10, -1.267901e-10, -1.271101e-10, -1.271885e-10, 
    -1.275622e-10, -1.272579e-10, -1.2776e-10, -1.273331e-10, -1.280721e-10, 
    -1.267441e-10, -1.273206e-10, -1.26276e-10, -1.263886e-10, -1.265922e-10, 
    -1.27059e-10, -1.268071e-10, -1.271018e-10, -1.264507e-10, -1.261128e-10, 
    -1.260254e-10, -1.258622e-10, -1.260291e-10, -1.260156e-10, 
    -1.261752e-10, -1.261239e-10, -1.265072e-10, -1.263014e-10, 
    -1.268861e-10, -1.270995e-10, -1.277018e-10, -1.280708e-10, 
    -1.284465e-10, -1.286123e-10, -1.286627e-10, -1.286838e-10 ;

 SMINN_TO_SOIL3N_S2 =
  -1.034011e-11, -1.036843e-11, -1.036293e-11, -1.038577e-11, -1.03731e-11, 
    -1.038806e-11, -1.034585e-11, -1.036956e-11, -1.035443e-11, 
    -1.034266e-11, -1.043008e-11, -1.038679e-11, -1.047505e-11, 
    -1.044745e-11, -1.051677e-11, -1.047075e-11, -1.052605e-11, 
    -1.051545e-11, -1.054736e-11, -1.053822e-11, -1.057902e-11, 
    -1.055158e-11, -1.060017e-11, -1.057247e-11, -1.05768e-11, -1.055067e-11, 
    -1.039551e-11, -1.042469e-11, -1.039378e-11, -1.039794e-11, 
    -1.039607e-11, -1.037336e-11, -1.036191e-11, -1.033794e-11, -1.03423e-11, 
    -1.03599e-11, -1.039981e-11, -1.038627e-11, -1.042041e-11, -1.041963e-11, 
    -1.045762e-11, -1.04405e-11, -1.050433e-11, -1.048619e-11, -1.05386e-11, 
    -1.052542e-11, -1.053798e-11, -1.053417e-11, -1.053803e-11, -1.05187e-11, 
    -1.052698e-11, -1.050998e-11, -1.04437e-11, -1.046318e-11, -1.040507e-11, 
    -1.037011e-11, -1.034689e-11, -1.033041e-11, -1.033274e-11, 
    -1.033718e-11, -1.036001e-11, -1.038147e-11, -1.039782e-11, 
    -1.040875e-11, -1.041952e-11, -1.045212e-11, -1.046937e-11, 
    -1.050799e-11, -1.050103e-11, -1.051283e-11, -1.052411e-11, 
    -1.054304e-11, -1.053993e-11, -1.054826e-11, -1.051252e-11, 
    -1.053628e-11, -1.049706e-11, -1.050779e-11, -1.042244e-11, 
    -1.038992e-11, -1.037609e-11, -1.036399e-11, -1.033453e-11, 
    -1.035487e-11, -1.034685e-11, -1.036593e-11, -1.037805e-11, 
    -1.037206e-11, -1.040905e-11, -1.039467e-11, -1.04704e-11, -1.043779e-11, 
    -1.05228e-11, -1.050246e-11, -1.052767e-11, -1.051481e-11, -1.053684e-11, 
    -1.051701e-11, -1.055137e-11, -1.055884e-11, -1.055373e-11, 
    -1.057337e-11, -1.051591e-11, -1.053798e-11, -1.037189e-11, 
    -1.037287e-11, -1.037742e-11, -1.03574e-11, -1.035617e-11, -1.033782e-11, 
    -1.035415e-11, -1.036111e-11, -1.037876e-11, -1.038919e-11, 
    -1.039911e-11, -1.042093e-11, -1.044528e-11, -1.047932e-11, 
    -1.050378e-11, -1.052017e-11, -1.051012e-11, -1.051899e-11, 
    -1.050907e-11, -1.050442e-11, -1.055604e-11, -1.052706e-11, 
    -1.057055e-11, -1.056814e-11, -1.054846e-11, -1.056841e-11, 
    -1.037355e-11, -1.036793e-11, -1.034839e-11, -1.036368e-11, 
    -1.033583e-11, -1.035142e-11, -1.036038e-11, -1.039497e-11, 
    -1.040257e-11, -1.040961e-11, -1.042352e-11, -1.044137e-11, 
    -1.047268e-11, -1.049991e-11, -1.052477e-11, -1.052295e-11, 
    -1.052359e-11, -1.052914e-11, -1.051539e-11, -1.05314e-11, -1.053408e-11, 
    -1.052706e-11, -1.056782e-11, -1.055617e-11, -1.056809e-11, 
    -1.056051e-11, -1.036976e-11, -1.037922e-11, -1.037411e-11, 
    -1.038373e-11, -1.037695e-11, -1.040707e-11, -1.041611e-11, 
    -1.045835e-11, -1.044102e-11, -1.046861e-11, -1.044383e-11, 
    -1.044822e-11, -1.04695e-11, -1.044517e-11, -1.049841e-11, -1.046231e-11, 
    -1.052935e-11, -1.049331e-11, -1.053161e-11, -1.052466e-11, 
    -1.053617e-11, -1.054648e-11, -1.055945e-11, -1.058337e-11, 
    -1.057783e-11, -1.059783e-11, -1.039334e-11, -1.040561e-11, 
    -1.040453e-11, -1.041737e-11, -1.042687e-11, -1.044746e-11, 
    -1.048046e-11, -1.046806e-11, -1.049084e-11, -1.049541e-11, -1.04608e-11, 
    -1.048205e-11, -1.041382e-11, -1.042485e-11, -1.041829e-11, -1.03943e-11, 
    -1.047091e-11, -1.04316e-11, -1.050418e-11, -1.048289e-11, -1.054501e-11, 
    -1.051412e-11, -1.057478e-11, -1.060069e-11, -1.062509e-11, 
    -1.065358e-11, -1.041231e-11, -1.040397e-11, -1.04189e-11, -1.043956e-11, 
    -1.045872e-11, -1.048419e-11, -1.04868e-11, -1.049157e-11, -1.050393e-11, 
    -1.051432e-11, -1.049308e-11, -1.051692e-11, -1.04274e-11, -1.047432e-11, 
    -1.040081e-11, -1.042295e-11, -1.043834e-11, -1.043159e-11, 
    -1.046664e-11, -1.047489e-11, -1.050844e-11, -1.04911e-11, -1.059429e-11, 
    -1.054865e-11, -1.067527e-11, -1.06399e-11, -1.040106e-11, -1.041228e-11, 
    -1.045134e-11, -1.043276e-11, -1.04859e-11, -1.049897e-11, -1.05096e-11, 
    -1.052318e-11, -1.052465e-11, -1.05327e-11, -1.051951e-11, -1.053218e-11, 
    -1.048425e-11, -1.050567e-11, -1.044688e-11, -1.046119e-11, 
    -1.045461e-11, -1.044738e-11, -1.046967e-11, -1.049341e-11, 
    -1.049392e-11, -1.050153e-11, -1.052296e-11, -1.048611e-11, 
    -1.060018e-11, -1.052974e-11, -1.042452e-11, -1.044613e-11, 
    -1.044922e-11, -1.044085e-11, -1.049766e-11, -1.047708e-11, -1.05325e-11, 
    -1.051753e-11, -1.054206e-11, -1.052987e-11, -1.052807e-11, 
    -1.051241e-11, -1.050266e-11, -1.047802e-11, -1.045797e-11, 
    -1.044207e-11, -1.044577e-11, -1.046323e-11, -1.049486e-11, 
    -1.052478e-11, -1.051823e-11, -1.05402e-11, -1.048204e-11, -1.050643e-11, 
    -1.0497e-11, -1.052158e-11, -1.046772e-11, -1.051357e-11, -1.0456e-11, 
    -1.046105e-11, -1.047667e-11, -1.050808e-11, -1.051504e-11, 
    -1.052245e-11, -1.051788e-11, -1.049567e-11, -1.049203e-11, 
    -1.047629e-11, -1.047194e-11, -1.045995e-11, -1.045002e-11, 
    -1.045909e-11, -1.046862e-11, -1.049568e-11, -1.052005e-11, 
    -1.054662e-11, -1.055313e-11, -1.058415e-11, -1.055889e-11, 
    -1.060057e-11, -1.056513e-11, -1.062647e-11, -1.051624e-11, 
    -1.056409e-11, -1.047738e-11, -1.048673e-11, -1.050363e-11, 
    -1.054238e-11, -1.052147e-11, -1.054593e-11, -1.049189e-11, 
    -1.046383e-11, -1.045658e-11, -1.044303e-11, -1.045689e-11, 
    -1.045576e-11, -1.046902e-11, -1.046476e-11, -1.049658e-11, 
    -1.047949e-11, -1.052803e-11, -1.054574e-11, -1.059573e-11, 
    -1.062637e-11, -1.065755e-11, -1.067131e-11, -1.06755e-11, -1.067725e-11 ;

 SMIN_NH4 =
  0.0005315545, 0.00053295, 0.0005326787, 0.0005338039, 0.0005331797, 
    0.0005339163, 0.0005318372, 0.0005330049, 0.0005322595, 0.0005316797, 
    0.000535986, 0.0005338537, 0.0005382006, 0.0005368413, 0.000540255, 
    0.0005379888, 0.0005407118, 0.0005401897, 0.0005417611, 0.0005413109, 
    0.0005433196, 0.0005419686, 0.0005443607, 0.000542997, 0.0005432102, 
    0.0005419237, 0.0005342835, 0.000535721, 0.0005341981, 0.0005344031, 
    0.0005343111, 0.0005331924, 0.0005326283, 0.0005314474, 0.0005316617, 
    0.0005325291, 0.000534495, 0.0005338278, 0.0005355091, 0.0005354712, 
    0.0005373421, 0.0005364986, 0.0005396422, 0.0005387489, 0.0005413296, 
    0.0005406807, 0.000541299, 0.0005411115, 0.0005413013, 0.0005403496, 
    0.0005407573, 0.0005399198, 0.0005366572, 0.0005376165, 0.0005347544, 
    0.0005330321, 0.0005318882, 0.0005310762, 0.0005311908, 0.0005314097, 
    0.0005325341, 0.0005335911, 0.0005343964, 0.000534935, 0.0005354656, 
    0.000537071, 0.0005379207, 0.0005398226, 0.0005394795, 0.0005400606, 
    0.000540616, 0.000541548, 0.0005413946, 0.0005418051, 0.0005400451, 
    0.0005412148, 0.0005392836, 0.0005398119, 0.0005356097, 0.000534008, 
    0.0005333265, 0.0005327303, 0.0005312791, 0.0005322812, 0.0005318861, 
    0.0005328259, 0.0005334229, 0.0005331276, 0.0005349496, 0.0005342413, 
    0.000537971, 0.0005363649, 0.0005405513, 0.0005395499, 0.0005407911, 
    0.0005401578, 0.0005412428, 0.0005402662, 0.0005419578, 0.000542326, 
    0.0005420743, 0.000543041, 0.0005402117, 0.0005412984, 0.0005331197, 
    0.0005331678, 0.0005333921, 0.0005324056, 0.0005323452, 0.0005314411, 
    0.0005322455, 0.000532588, 0.0005334574, 0.0005339715, 0.0005344601, 
    0.0005355345, 0.0005367338, 0.0005384104, 0.0005396147, 0.0005404216, 
    0.0005399268, 0.0005403636, 0.0005398752, 0.0005396463, 0.0005421878, 
    0.0005407608, 0.0005429017, 0.0005427834, 0.0005418144, 0.0005427966, 
    0.0005332015, 0.0005329243, 0.0005319619, 0.000532715, 0.0005313426, 
    0.0005321107, 0.0005325523, 0.0005342559, 0.0005346302, 0.0005349771, 
    0.0005356623, 0.0005365413, 0.0005380831, 0.0005394242, 0.0005406481, 
    0.0005405584, 0.0005405899, 0.0005408631, 0.000540186, 0.0005409742, 
    0.0005411064, 0.0005407606, 0.0005427673, 0.0005421941, 0.0005427806, 
    0.0005424073, 0.0005330144, 0.0005334805, 0.0005332285, 0.0005337023, 
    0.0005333684, 0.0005348523, 0.000535297, 0.0005373778, 0.0005365241, 
    0.0005378829, 0.000536662, 0.0005368784, 0.0005379267, 0.0005367279, 
    0.0005393499, 0.0005375721, 0.0005408737, 0.0005390988, 0.0005409848, 
    0.0005406424, 0.0005412091, 0.0005417166, 0.0005423551, 0.0005435327, 
    0.00054326, 0.0005442448, 0.0005341756, 0.00053478, 0.0005347269, 
    0.0005353595, 0.0005358272, 0.0005368412, 0.0005384666, 0.0005378554, 
    0.0005389773, 0.0005392025, 0.0005374978, 0.0005385444, 0.0005351841, 
    0.000535727, 0.0005354038, 0.0005342223, 0.0005379956, 0.0005360594, 
    0.0005396339, 0.0005385856, 0.0005416441, 0.0005401232, 0.0005431098, 
    0.0005443856, 0.0005455865, 0.0005469888, 0.00053511, 0.0005346992, 
    0.0005354346, 0.0005364519, 0.0005373957, 0.0005386501, 0.0005387785, 
    0.0005390133, 0.0005396218, 0.0005401333, 0.0005390873, 0.0005402614, 
    0.0005358526, 0.0005381636, 0.0005345431, 0.0005356334, 0.0005363912, 
    0.0005360589, 0.0005377848, 0.0005381914, 0.0005398433, 0.0005389896, 
    0.0005440706, 0.0005418233, 0.0005480565, 0.0005463155, 0.0005345556, 
    0.0005351084, 0.0005370321, 0.0005361169, 0.0005387338, 0.0005393776, 
    0.000539901, 0.0005405698, 0.000540642, 0.0005410382, 0.0005403887, 
    0.0005410125, 0.0005386522, 0.0005397071, 0.0005368118, 0.0005375165, 
    0.0005371923, 0.0005368365, 0.0005379342, 0.0005391031, 0.0005391283, 
    0.0005395029, 0.0005405582, 0.0005387434, 0.0005443599, 0.0005408918, 
    0.0005357112, 0.0005367756, 0.0005369278, 0.0005365154, 0.0005393129, 
    0.0005382995, 0.0005410286, 0.0005402911, 0.0005414992, 0.0005408989, 
    0.0005408104, 0.0005400393, 0.0005395589, 0.0005383455, 0.0005373578, 
    0.0005365746, 0.0005367566, 0.000537617, 0.0005391745, 0.0005406477, 
    0.000540325, 0.0005414067, 0.000538543, 0.0005397439, 0.0005392796, 
    0.0005404899, 0.0005378389, 0.0005400968, 0.0005372614, 0.00053751, 
    0.0005382792, 0.0005398261, 0.0005401684, 0.0005405336, 0.0005403081, 
    0.0005392145, 0.0005390353, 0.0005382602, 0.000538046, 0.0005374554, 
    0.0005369661, 0.000537413, 0.0005378821, 0.0005392146, 0.0005404149, 
    0.0005417232, 0.0005420434, 0.0005435708, 0.0005423271, 0.0005443789, 
    0.0005426341, 0.0005456542, 0.0005402278, 0.0005425842, 0.0005383143, 
    0.0005387745, 0.0005396066, 0.0005415149, 0.0005404848, 0.0005416895, 
    0.0005390283, 0.0005376466, 0.0005372892, 0.0005366221, 0.0005373044, 
    0.0005372489, 0.0005379017, 0.0005376918, 0.0005392587, 0.0005384171, 
    0.0005408074, 0.0005416794, 0.0005441409, 0.000545649, 0.0005471839, 
    0.0005478612, 0.0005480674, 0.0005481535 ;

 SMIN_NH4_vr =
  0.002921869, 0.002926673, 0.002925733, 0.002929604, 0.002927454, 
    0.002929982, 0.002922828, 0.002926841, 0.002924276, 0.002922276, 
    0.002937075, 0.002929752, 0.002944677, 0.002940009, 0.002951712, 
    0.002943942, 0.002953274, 0.002951483, 0.002956863, 0.002955317, 
    0.002962184, 0.002957566, 0.002965739, 0.002961077, 0.002961802, 
    0.002957398, 0.002931251, 0.002936187, 0.002930952, 0.002931657, 
    0.002931337, 0.002927484, 0.002925541, 0.002921474, 0.002922208, 
    0.002925193, 0.002931951, 0.002929654, 0.002935429, 0.0029353, 
    0.002941717, 0.002938822, 0.002949603, 0.002946536, 0.002955378, 
    0.002953151, 0.002955267, 0.002954621, 0.002955267, 0.002952007, 
    0.002953397, 0.002950529, 0.002939401, 0.002942689, 0.002932858, 
    0.002926928, 0.002922991, 0.002920196, 0.002920585, 0.002921338, 
    0.002925204, 0.002928837, 0.002931606, 0.002933452, 0.002935272, 
    0.002940782, 0.002943696, 0.002950213, 0.002949038, 0.002951024, 
    0.002952926, 0.002956113, 0.002955587, 0.002956987, 0.002950956, 
    0.002954962, 0.002948341, 0.002950152, 0.00293579, 0.002930287, 
    0.002927938, 0.002925885, 0.002920886, 0.002924336, 0.002922972, 
    0.002926203, 0.002928256, 0.002927236, 0.002933499, 0.00293106, 
    0.002943864, 0.002938352, 0.002952708, 0.002949272, 0.002953522, 
    0.002951353, 0.002955062, 0.002951718, 0.002957504, 0.002958764, 
    0.002957897, 0.002961205, 0.002951514, 0.002955235, 0.002927225, 
    0.002927391, 0.002928159, 0.002924759, 0.002924551, 0.002921434, 
    0.0029242, 0.002925379, 0.002928367, 0.00293013, 0.002931806, 
    0.002935498, 0.002939613, 0.002945362, 0.002949491, 0.002952252, 
    0.002950555, 0.002952047, 0.002950372, 0.002949584, 0.002958283, 
    0.002953398, 0.002960721, 0.002960316, 0.002956996, 0.002960353, 
    0.002927501, 0.002926544, 0.002923229, 0.002925818, 0.002921089, 
    0.002923734, 0.002925249, 0.002931104, 0.002932389, 0.002933581, 
    0.002935932, 0.002938947, 0.002944236, 0.002948831, 0.002953025, 
    0.002952713, 0.002952819, 0.00295375, 0.002951429, 0.002954125, 
    0.002954573, 0.00295339, 0.002960253, 0.002958292, 0.002960295, 
    0.002959014, 0.00292685, 0.002928449, 0.002927578, 0.002929208, 
    0.002928053, 0.002933155, 0.002934679, 0.00294182, 0.002938887, 
    0.002943551, 0.002939355, 0.002940098, 0.002943689, 0.002939574, 
    0.002948566, 0.002942463, 0.002953783, 0.002947693, 0.002954158, 
    0.002952981, 0.002954918, 0.002956656, 0.002958834, 0.002962862, 
    0.002961924, 0.002965291, 0.002930836, 0.002932908, 0.002932726, 
    0.002934895, 0.002936497, 0.002939981, 0.002945554, 0.002943453, 
    0.002947298, 0.00294807, 0.002942217, 0.002945807, 0.002934267, 
    0.002936126, 0.002935017, 0.002930951, 0.002943908, 0.002937257, 
    0.002949522, 0.002945923, 0.002956399, 0.002951189, 0.002961408, 
    0.002965768, 0.002969869, 0.002974648, 0.00293404, 0.002932624, 
    0.002935147, 0.00293864, 0.002941875, 0.002946179, 0.002946616, 
    0.002947417, 0.002949499, 0.002951253, 0.002947662, 0.002951683, 
    0.002936552, 0.002944484, 0.002932048, 0.002935794, 0.002938391, 
    0.002937251, 0.002943174, 0.002944564, 0.002950222, 0.002947298, 
    0.002964682, 0.002956997, 0.002978286, 0.002972346, 0.002932127, 
    0.002934023, 0.002940624, 0.002937483, 0.002946458, 0.002948666, 
    0.002950454, 0.002952745, 0.002952987, 0.002954344, 0.002952114, 
    0.002954251, 0.002946155, 0.002949773, 0.002939838, 0.002942251, 
    0.002941138, 0.002939912, 0.002943675, 0.002947683, 0.002947767, 
    0.002949046, 0.002952655, 0.002946437, 0.002965656, 0.002953788, 
    0.00293609, 0.002939739, 0.002940259, 0.002938845, 0.002948436, 
    0.002944961, 0.002954311, 0.002951781, 0.002955914, 0.00295386, 
    0.00295355, 0.002950909, 0.002949256, 0.002945096, 0.0029417, 
    0.002939013, 0.002939632, 0.002942584, 0.00294792, 0.00295297, 
    0.002951859, 0.002955561, 0.002945744, 0.002949861, 0.002948263, 
    0.002952412, 0.002943384, 0.002951121, 0.0029414, 0.002942248, 
    0.002944883, 0.002950185, 0.002951354, 0.002952605, 0.002951828, 
    0.002948079, 0.002947461, 0.002944799, 0.00294406, 0.002942035, 
    0.002940349, 0.002941883, 0.002943486, 0.002948057, 0.002952166, 
    0.002956642, 0.002957737, 0.002962953, 0.002958699, 0.002965707, 
    0.002959739, 0.002970059, 0.002951564, 0.002959632, 0.002945004, 
    0.002946578, 0.002949428, 0.00295596, 0.002952431, 0.002956555, 
    0.002947435, 0.00294269, 0.002941462, 0.002939172, 0.002941508, 
    0.002941318, 0.002943554, 0.00294283, 0.002948199, 0.002945315, 
    0.0029535, 0.002956486, 0.002964902, 0.002970048, 0.002975288, 
    0.002977593, 0.002978295, 0.002978585,
  0.001884459, 0.001889418, 0.001888455, 0.00189245, 0.001890235, 0.00189285, 
    0.001885466, 0.001889614, 0.001886967, 0.001884907, 0.001900191, 
    0.001892629, 0.001908041, 0.001903227, 0.001915312, 0.001907291, 
    0.001916928, 0.001915083, 0.001920638, 0.001919047, 0.00192614, 
    0.001921372, 0.001929815, 0.001925003, 0.001925756, 0.001921214, 
    0.001894154, 0.00189925, 0.001893851, 0.001894578, 0.001894252, 
    0.00189028, 0.001888276, 0.001884081, 0.001884843, 0.001887925, 
    0.001894905, 0.001892538, 0.001898505, 0.001898371, 0.001905003, 
    0.001902014, 0.001913146, 0.001909986, 0.001919114, 0.00191682, 
    0.001919006, 0.001918343, 0.001919014, 0.00191565, 0.001917091, 
    0.00191413, 0.001902573, 0.001905972, 0.001895825, 0.001889709, 
    0.001885647, 0.001882761, 0.001883169, 0.001883947, 0.001887943, 
    0.001891698, 0.001894557, 0.001896469, 0.001898351, 0.00190404, 
    0.001907051, 0.001913784, 0.001912571, 0.001914627, 0.001916592, 
    0.001919886, 0.001919344, 0.001920795, 0.001914574, 0.001918709, 
    0.00191188, 0.001913749, 0.001898856, 0.001893177, 0.001890756, 
    0.00188864, 0.001883483, 0.001887044, 0.001885641, 0.001888981, 
    0.001891101, 0.001890053, 0.001896521, 0.001894007, 0.00190723, 
    0.00190154, 0.001916362, 0.001912821, 0.001917211, 0.001914972, 
    0.001918808, 0.001915356, 0.001921335, 0.001922635, 0.001921746, 
    0.001925161, 0.001915164, 0.001919005, 0.001890023, 0.001890194, 
    0.001890991, 0.001887486, 0.001887272, 0.00188406, 0.001886919, 
    0.001888136, 0.001891225, 0.00189305, 0.001894784, 0.001898596, 
    0.001902847, 0.001908787, 0.00191305, 0.001915905, 0.001914155, 
    0.0019157, 0.001913973, 0.001913163, 0.001922147, 0.001917104, 
    0.00192467, 0.001924252, 0.001920829, 0.001924299, 0.001890314, 
    0.00188933, 0.00188591, 0.001888587, 0.00188371, 0.00188644, 0.001888008, 
    0.001894058, 0.001895388, 0.001896619, 0.00189905, 0.001902167, 
    0.001907629, 0.001912376, 0.001916706, 0.001916389, 0.001916501, 
    0.001917467, 0.001915072, 0.00191786, 0.001918327, 0.001917105, 
    0.001924196, 0.001922171, 0.001924243, 0.001922925, 0.001889651, 
    0.001891306, 0.001890411, 0.001892093, 0.001890908, 0.001896175, 
    0.001897752, 0.001905129, 0.001902105, 0.001906919, 0.001902595, 
    0.001903361, 0.001907073, 0.001902829, 0.001912113, 0.001905819, 
    0.001917504, 0.001911224, 0.001917897, 0.001916687, 0.001918691, 
    0.001920484, 0.00192274, 0.001926897, 0.001925935, 0.001929411, 
    0.001893774, 0.001895919, 0.001895731, 0.001897976, 0.001899634, 
    0.001903229, 0.001908987, 0.001906823, 0.001910796, 0.001911592, 
    0.001905557, 0.001909263, 0.001897354, 0.001899279, 0.001898134, 
    0.001893942, 0.00190732, 0.001900459, 0.00191312, 0.001909411, 
    0.001920228, 0.001914851, 0.001925405, 0.001929906, 0.001934142, 
    0.001939081, 0.00189709, 0.001895633, 0.001898243, 0.001901848, 
    0.001905194, 0.001909637, 0.001910092, 0.001910923, 0.001913077, 
    0.001914886, 0.001911184, 0.00191534, 0.001899723, 0.001907915, 
    0.001895081, 0.001898948, 0.001901636, 0.001900458, 0.001906576, 
    0.001908016, 0.001913862, 0.001910842, 0.001928794, 0.001920861, 
    0.001942841, 0.00193671, 0.001895124, 0.001897086, 0.001903906, 
    0.001900662, 0.001909934, 0.001912212, 0.001914065, 0.001916429, 
    0.001916685, 0.001918086, 0.00191579, 0.001917996, 0.001909646, 
    0.00191338, 0.001903128, 0.001905625, 0.001904477, 0.001903216, 
    0.001907105, 0.001911242, 0.001911333, 0.001912658, 0.001916387, 
    0.001909971, 0.001929813, 0.001917567, 0.001899224, 0.001902996, 
    0.001903537, 0.001902076, 0.001911984, 0.001908396, 0.001918052, 
    0.001915445, 0.001919716, 0.001917594, 0.001917282, 0.001914555, 
    0.001912856, 0.00190856, 0.001905063, 0.001902288, 0.001902934, 
    0.001905981, 0.001911496, 0.001916707, 0.001915566, 0.001919392, 
    0.001909262, 0.001913512, 0.001911869, 0.001916151, 0.001906765, 
    0.001914753, 0.00190472, 0.001905601, 0.001908325, 0.001913798, 
    0.001915011, 0.001916302, 0.001915506, 0.001911636, 0.001911003, 
    0.001908259, 0.001907501, 0.001905409, 0.001903676, 0.001905259, 
    0.001906921, 0.001911639, 0.001915885, 0.00192051, 0.001921641, 
    0.001927032, 0.001922641, 0.001929881, 0.001923723, 0.001934379, 
    0.001915218, 0.001923545, 0.00190845, 0.001910079, 0.001913023, 
    0.00191977, 0.001916131, 0.001920387, 0.001910978, 0.001906085, 
    0.001904821, 0.001902456, 0.001904875, 0.001904678, 0.001906991, 
    0.001906248, 0.001911795, 0.001908816, 0.001917273, 0.001920354, 
    0.001929046, 0.001934363, 0.001939772, 0.001942156, 0.001942882, 
    0.001943185,
  0.001890241, 0.001895266, 0.00189429, 0.001898339, 0.001896093, 
    0.001898744, 0.001891261, 0.001895464, 0.001892782, 0.001890694, 
    0.001906187, 0.00189852, 0.001914145, 0.001909263, 0.00192152, 
    0.001913385, 0.001923159, 0.001921287, 0.001926923, 0.001925309, 
    0.001932508, 0.001927667, 0.001936238, 0.001931353, 0.001932117, 
    0.001927507, 0.001900065, 0.001905232, 0.001899758, 0.001900495, 
    0.001900165, 0.001896139, 0.001894109, 0.001889858, 0.00189063, 
    0.001893753, 0.001900827, 0.001898427, 0.001904475, 0.001904339, 
    0.001911063, 0.001908032, 0.001919322, 0.001916116, 0.001925376, 
    0.001923049, 0.001925267, 0.001924595, 0.001925275, 0.001921862, 
    0.001923325, 0.00192032, 0.0019086, 0.001912047, 0.001901759, 
    0.001895562, 0.001891445, 0.001888521, 0.001888934, 0.001889722, 
    0.001893771, 0.001897576, 0.001900474, 0.001902411, 0.001904319, 
    0.001910088, 0.001913141, 0.00191997, 0.001918739, 0.001920824, 
    0.001922817, 0.00192616, 0.00192561, 0.001927082, 0.00192077, 
    0.001924965, 0.001918038, 0.001919933, 0.001904833, 0.001899075, 
    0.001896622, 0.001894477, 0.001889252, 0.001892861, 0.001891438, 
    0.001894822, 0.001896971, 0.001895909, 0.001902464, 0.001899916, 
    0.001913322, 0.001907552, 0.001922585, 0.001918992, 0.001923446, 
    0.001921174, 0.001925066, 0.001921563, 0.00192763, 0.00192895, 
    0.001928048, 0.001931512, 0.001921369, 0.001925266, 0.001895879, 
    0.001896052, 0.00189686, 0.001893308, 0.001893091, 0.001889836, 
    0.001892733, 0.001893966, 0.001897096, 0.001898946, 0.001900704, 
    0.001904567, 0.001908878, 0.001914901, 0.001919225, 0.001922121, 
    0.001920345, 0.001921913, 0.00192016, 0.001919339, 0.001928455, 
    0.001923338, 0.001931014, 0.00193059, 0.001927117, 0.001930638, 
    0.001896174, 0.001895176, 0.001891711, 0.001894423, 0.001889482, 
    0.001892248, 0.001893837, 0.001899968, 0.001901316, 0.001902563, 
    0.001905027, 0.001908187, 0.001913726, 0.001918541, 0.001922933, 
    0.001922612, 0.001922725, 0.001923705, 0.001921276, 0.001924104, 
    0.001924578, 0.001923338, 0.001930533, 0.001928479, 0.001930581, 
    0.001929244, 0.001895501, 0.001897179, 0.001896272, 0.001897977, 
    0.001896776, 0.001902114, 0.001903713, 0.001911192, 0.001908125, 
    0.001913007, 0.001908621, 0.001909399, 0.001913164, 0.001908859, 
    0.001918275, 0.001911891, 0.001923743, 0.001917374, 0.001924142, 
    0.001922914, 0.001924947, 0.001926767, 0.001929056, 0.001933276, 
    0.001932299, 0.001935827, 0.00189968, 0.001901854, 0.001901663, 
    0.001903938, 0.00190562, 0.001909265, 0.001915103, 0.001912909, 
    0.001916938, 0.001917746, 0.001911625, 0.001915383, 0.001903309, 
    0.001905261, 0.0019041, 0.001899851, 0.001913413, 0.001906457, 
    0.001919296, 0.001915533, 0.001926507, 0.001921052, 0.001931761, 
    0.00193633, 0.00194063, 0.001945646, 0.001903041, 0.001901564, 
    0.001904209, 0.001907865, 0.001911258, 0.001915763, 0.001916224, 
    0.001917067, 0.001919252, 0.001921087, 0.001917333, 0.001921547, 
    0.001905712, 0.001914017, 0.001901005, 0.001904925, 0.00190765, 
    0.001906456, 0.001912658, 0.001914118, 0.001920048, 0.001916984, 
    0.001935202, 0.00192715, 0.001949465, 0.001943239, 0.001901048, 
    0.001903036, 0.001909951, 0.001906662, 0.001916064, 0.001918375, 
    0.001920254, 0.001922653, 0.001922912, 0.001924333, 0.001922004, 
    0.001924242, 0.001915772, 0.001919559, 0.001909162, 0.001911694, 
    0.00191053, 0.001909252, 0.001913195, 0.001917392, 0.001917483, 
    0.001918827, 0.001922612, 0.001916102, 0.001936238, 0.001923809, 
    0.001905204, 0.001909029, 0.001909577, 0.001908095, 0.001918143, 
    0.001914504, 0.001924299, 0.001921654, 0.001925987, 0.001923834, 
    0.001923517, 0.001920751, 0.001919028, 0.001914671, 0.001911124, 
    0.00190831, 0.001908965, 0.001912055, 0.001917648, 0.001922935, 
    0.001921777, 0.001925658, 0.001915382, 0.001919693, 0.001918027, 
    0.00192237, 0.00191285, 0.001920954, 0.001910776, 0.00191167, 
    0.001914432, 0.001919984, 0.001921214, 0.001922524, 0.001921716, 
    0.001917791, 0.001917148, 0.001914365, 0.001913596, 0.001911475, 
    0.001909718, 0.001911323, 0.001913008, 0.001917793, 0.0019221, 
    0.001926793, 0.001927941, 0.001933413, 0.001928957, 0.001936307, 
    0.001930056, 0.001940873, 0.001921425, 0.001929875, 0.001914558, 
    0.001916211, 0.001919197, 0.001926043, 0.00192235, 0.001926669, 
    0.001917123, 0.001912161, 0.001910878, 0.001908481, 0.001910933, 
    0.001910734, 0.001913079, 0.001912326, 0.001917952, 0.00191493, 
    0.001923509, 0.001926636, 0.001935457, 0.001940855, 0.001946347, 
    0.001948769, 0.001949506, 0.001949814,
  0.001831959, 0.001836913, 0.00183595, 0.001839945, 0.001837729, 
    0.001840344, 0.001832964, 0.00183711, 0.001834463, 0.001832405, 
    0.001847691, 0.001840123, 0.001855548, 0.001850726, 0.001862836, 
    0.001854797, 0.001864456, 0.001862605, 0.001868177, 0.001866581, 
    0.001873703, 0.001868913, 0.001877394, 0.00187256, 0.001873316, 
    0.001868755, 0.001841647, 0.001846749, 0.001841344, 0.001842072, 
    0.001841746, 0.001837775, 0.001835773, 0.00183158, 0.001832342, 
    0.001835421, 0.001842399, 0.001840031, 0.001845999, 0.001845864, 
    0.001852503, 0.001849511, 0.001860663, 0.001857495, 0.001866647, 
    0.001864346, 0.001866539, 0.001865874, 0.001866548, 0.001863173, 
    0.001864619, 0.001861649, 0.001850071, 0.001853475, 0.001843319, 
    0.001837206, 0.001833146, 0.001830262, 0.00183067, 0.001831447, 
    0.001835439, 0.001839192, 0.00184205, 0.001843962, 0.001845845, 
    0.001851542, 0.001854557, 0.001861303, 0.001860086, 0.001862148, 
    0.001864117, 0.001867422, 0.001866879, 0.001868334, 0.001862094, 
    0.001866242, 0.001859393, 0.001861267, 0.001846355, 0.00184067, 
    0.001838252, 0.001836135, 0.001830983, 0.001834541, 0.001833139, 
    0.001836476, 0.001838595, 0.001837547, 0.001844014, 0.0018415, 
    0.001854735, 0.001849037, 0.001863888, 0.001860336, 0.001864739, 
    0.001862493, 0.001866341, 0.001862878, 0.001868876, 0.001870182, 
    0.00186929, 0.001872717, 0.001862685, 0.001866539, 0.001837517, 
    0.001837688, 0.001838485, 0.001834983, 0.001834769, 0.001831559, 
    0.001834416, 0.001835631, 0.001838718, 0.001840543, 0.001842277, 
    0.00184609, 0.001850346, 0.001856295, 0.001860566, 0.001863429, 
    0.001861674, 0.001863223, 0.001861491, 0.001860679, 0.001869693, 
    0.001864632, 0.001872224, 0.001871804, 0.001868369, 0.001871852, 
    0.001837808, 0.001836825, 0.001833408, 0.001836082, 0.00183121, 
    0.001833937, 0.001835505, 0.001841552, 0.001842881, 0.001844112, 
    0.001846544, 0.001849664, 0.001855134, 0.001859891, 0.001864232, 
    0.001863914, 0.001864026, 0.001864995, 0.001862594, 0.001865389, 
    0.001865858, 0.001864632, 0.001871748, 0.001869716, 0.001871795, 
    0.001870472, 0.001837144, 0.0018388, 0.001837905, 0.001839587, 
    0.001838402, 0.001843669, 0.001845248, 0.001852631, 0.001849602, 
    0.001854423, 0.001850092, 0.00185086, 0.00185458, 0.001850327, 
    0.001859628, 0.001853322, 0.001865033, 0.001858738, 0.001865427, 
    0.001864213, 0.001866223, 0.001868023, 0.001870287, 0.001874462, 
    0.001873496, 0.001876986, 0.001841267, 0.001843413, 0.001843224, 
    0.001845469, 0.001847129, 0.001850727, 0.001856494, 0.001854326, 
    0.001858306, 0.001859105, 0.001853058, 0.001856771, 0.001844849, 
    0.001846775, 0.001845628, 0.001841436, 0.001854825, 0.001847956, 
    0.001860637, 0.001856919, 0.001867766, 0.001862373, 0.001872963, 
    0.001877486, 0.001881742, 0.001886712, 0.001844584, 0.001843126, 
    0.001845736, 0.001849346, 0.001852695, 0.001857145, 0.001857601, 
    0.001858434, 0.001860593, 0.001862407, 0.001858697, 0.001862862, 
    0.001847222, 0.001855421, 0.001842575, 0.001846444, 0.001849134, 
    0.001847954, 0.001854078, 0.001855521, 0.001861381, 0.001858352, 
    0.00187637, 0.001868403, 0.001890495, 0.001884326, 0.001842617, 
    0.001844579, 0.001851405, 0.001848158, 0.001857443, 0.001859726, 
    0.001861583, 0.001863955, 0.001864211, 0.001865616, 0.001863314, 
    0.001865525, 0.001857155, 0.001860896, 0.001850626, 0.001853126, 
    0.001851976, 0.001850714, 0.001854609, 0.001858755, 0.001858845, 
    0.001860174, 0.001863917, 0.00185748, 0.001877396, 0.001865101, 
    0.001846718, 0.001850496, 0.001851036, 0.001849573, 0.001859497, 
    0.001855902, 0.001865582, 0.001862967, 0.001867251, 0.001865123, 
    0.00186481, 0.001862075, 0.001860371, 0.001856067, 0.001852564, 
    0.001849785, 0.001850431, 0.001853483, 0.001859009, 0.001864234, 
    0.00186309, 0.001866926, 0.00185677, 0.001861029, 0.001859383, 
    0.001863675, 0.001854268, 0.001862278, 0.00185222, 0.001853102, 
    0.001855831, 0.001861318, 0.001862532, 0.001863828, 0.001863028, 
    0.00185915, 0.001858514, 0.001855765, 0.001855005, 0.00185291, 
    0.001851175, 0.00185276, 0.001854425, 0.001859151, 0.001863409, 
    0.001868048, 0.001869184, 0.0018746, 0.00187019, 0.001877465, 
    0.001871279, 0.001881985, 0.001862743, 0.001871098, 0.001855955, 
    0.001857588, 0.00186054, 0.001867308, 0.001863655, 0.001867927, 
    0.001858489, 0.001853588, 0.001852321, 0.001849954, 0.001852375, 
    0.001852178, 0.001854494, 0.00185375, 0.001859308, 0.001856323, 
    0.001864802, 0.001867894, 0.00187662, 0.001881966, 0.001887405, 
    0.001889805, 0.001890535, 0.001890841,
  0.001659593, 0.001664243, 0.001663339, 0.001667091, 0.00166501, 
    0.001667466, 0.001660536, 0.001664428, 0.001661943, 0.001660012, 
    0.001674374, 0.001667258, 0.001681769, 0.001677228, 0.001688639, 
    0.001681063, 0.001690167, 0.00168842, 0.001693678, 0.001692172, 
    0.001698899, 0.001694373, 0.001702388, 0.001697818, 0.001698533, 
    0.001694224, 0.00166869, 0.001673488, 0.001668406, 0.00166909, 
    0.001668783, 0.001665053, 0.001663173, 0.001659238, 0.001659952, 
    0.001662843, 0.001669397, 0.001667172, 0.001672781, 0.001672655, 
    0.001678902, 0.001676085, 0.001686589, 0.001683603, 0.001692234, 
    0.001690063, 0.001692132, 0.001691505, 0.001692141, 0.001688956, 
    0.001690321, 0.001687519, 0.001676612, 0.001679817, 0.001670262, 
    0.001664519, 0.001660706, 0.001658001, 0.001658384, 0.001659113, 
    0.00166286, 0.001666383, 0.001669069, 0.001670866, 0.001672636, 
    0.001677998, 0.001680836, 0.001687193, 0.001686046, 0.00168799, 
    0.001689847, 0.001692966, 0.001692453, 0.001693827, 0.001687938, 
    0.001691852, 0.001685392, 0.001687158, 0.001673118, 0.001667772, 
    0.001665501, 0.001663513, 0.001658678, 0.001662017, 0.0016607, 
    0.001663832, 0.001665822, 0.001664838, 0.001670915, 0.001668552, 
    0.001681004, 0.001675639, 0.00168963, 0.001686281, 0.001690433, 
    0.001688314, 0.001691945, 0.001688677, 0.001694339, 0.001695572, 
    0.001694729, 0.001697966, 0.001688496, 0.001692132, 0.00166481, 
    0.001664971, 0.001665719, 0.001662431, 0.00166223, 0.001659218, 
    0.001661898, 0.00166304, 0.001665938, 0.001667652, 0.001669282, 
    0.001672867, 0.001676871, 0.001682473, 0.001686498, 0.001689197, 
    0.001687542, 0.001689003, 0.00168737, 0.001686604, 0.00169511, 
    0.001690333, 0.001697501, 0.001697104, 0.00169386, 0.001697149, 
    0.001665084, 0.00166416, 0.001660953, 0.001663463, 0.00165889, 
    0.001661449, 0.001662921, 0.001668601, 0.00166985, 0.001671007, 
    0.001673294, 0.001676229, 0.001681379, 0.001685862, 0.001689955, 
    0.001689655, 0.001689761, 0.001690676, 0.00168841, 0.001691047, 
    0.00169149, 0.001690333, 0.001697051, 0.001695131, 0.001697096, 
    0.001695846, 0.00166446, 0.001666015, 0.001665175, 0.001666754, 
    0.001665642, 0.001670591, 0.001672075, 0.001679023, 0.001676171, 
    0.00168071, 0.001676632, 0.001677355, 0.001680858, 0.001676852, 
    0.001685615, 0.001679674, 0.001690711, 0.001684776, 0.001691083, 
    0.001689938, 0.001691834, 0.001693533, 0.001695671, 0.001699616, 
    0.001698702, 0.001702002, 0.001668333, 0.00167035, 0.001670172, 
    0.001672283, 0.001673845, 0.00167723, 0.00168266, 0.001680618, 
    0.001684368, 0.001685121, 0.001679424, 0.001682921, 0.0016717, 
    0.001673512, 0.001672433, 0.001668492, 0.001681088, 0.001674623, 
    0.001686565, 0.00168306, 0.001693291, 0.001688202, 0.001698199, 
    0.001702476, 0.001706502, 0.001711208, 0.001671451, 0.00167008, 
    0.001672534, 0.00167593, 0.001679082, 0.001683274, 0.001683703, 
    0.001684488, 0.001686523, 0.001688234, 0.001684737, 0.001688663, 
    0.001673933, 0.00168165, 0.001669562, 0.001673201, 0.00167573, 
    0.001674621, 0.001680384, 0.001681743, 0.001687266, 0.001684411, 
    0.00170142, 0.001693892, 0.001714793, 0.001708949, 0.001669601, 
    0.001671446, 0.001677868, 0.001674812, 0.001683554, 0.001685706, 
    0.001687456, 0.001689694, 0.001689936, 0.001691262, 0.001689089, 
    0.001691176, 0.001683283, 0.001686809, 0.001677134, 0.001679488, 
    0.001678405, 0.001677217, 0.001680884, 0.001684792, 0.001684875, 
    0.001686128, 0.001689661, 0.001683589, 0.001702392, 0.001690777, 
    0.001673458, 0.001677012, 0.00167752, 0.001676143, 0.00168549, 
    0.001682103, 0.001691229, 0.001688762, 0.001692805, 0.001690796, 
    0.0016905, 0.00168792, 0.001686314, 0.001682258, 0.001678959, 
    0.001676343, 0.001676951, 0.001679825, 0.001685031, 0.001689958, 
    0.001688878, 0.001692497, 0.00168292, 0.001686935, 0.001685383, 
    0.00168943, 0.001680564, 0.001688114, 0.001678634, 0.001679465, 
    0.001682036, 0.001687207, 0.001688352, 0.001689574, 0.00168882, 
    0.001685163, 0.001684564, 0.001681973, 0.001681258, 0.001679284, 
    0.00167765, 0.001679143, 0.001680711, 0.001685164, 0.001689179, 
    0.001693557, 0.001694629, 0.001699747, 0.001695581, 0.001702457, 
    0.001696611, 0.001706733, 0.001688552, 0.001696439, 0.001682153, 
    0.001683691, 0.001686474, 0.001692859, 0.001689411, 0.001693443, 
    0.00168454, 0.001679924, 0.001678729, 0.001676502, 0.00167878, 
    0.001678595, 0.001680776, 0.001680075, 0.001685312, 0.001682499, 
    0.001690493, 0.001693411, 0.001701656, 0.001706714, 0.001711864, 
    0.001714138, 0.001714831, 0.00171512,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3 =
  1.823172e-06, 1.833022e-06, 1.831105e-06, 1.839062e-06, 1.834647e-06, 
    1.839859e-06, 1.825167e-06, 1.833412e-06, 1.828147e-06, 1.824058e-06, 
    1.854546e-06, 1.839417e-06, 1.870326e-06, 1.860632e-06, 1.885027e-06, 
    1.868815e-06, 1.888304e-06, 1.88456e-06, 1.895842e-06, 1.892607e-06, 
    1.907068e-06, 1.897336e-06, 1.914586e-06, 1.904742e-06, 1.90628e-06, 
    1.897014e-06, 1.842459e-06, 1.85266e-06, 1.841855e-06, 1.843308e-06, 
    1.842656e-06, 1.834737e-06, 1.830751e-06, 1.82242e-06, 1.823931e-06, 
    1.830051e-06, 1.84396e-06, 1.839234e-06, 1.851158e-06, 1.850888e-06, 
    1.864202e-06, 1.858194e-06, 1.880637e-06, 1.874246e-06, 1.892741e-06, 
    1.888082e-06, 1.892522e-06, 1.891175e-06, 1.892539e-06, 1.885708e-06, 
    1.888633e-06, 1.882627e-06, 1.85932e-06, 1.866156e-06, 1.845798e-06, 
    1.833604e-06, 1.825528e-06, 1.819805e-06, 1.820614e-06, 1.822155e-06, 
    1.830087e-06, 1.837559e-06, 1.843263e-06, 1.847082e-06, 1.850849e-06, 
    1.86227e-06, 1.86833e-06, 1.881929e-06, 1.879473e-06, 1.883636e-06, 
    1.887619e-06, 1.894312e-06, 1.89321e-06, 1.896161e-06, 1.883526e-06, 
    1.891918e-06, 1.878073e-06, 1.881855e-06, 1.851871e-06, 1.840509e-06, 
    1.835686e-06, 1.831472e-06, 1.821235e-06, 1.828301e-06, 1.825514e-06, 
    1.832149e-06, 1.83637e-06, 1.834281e-06, 1.847186e-06, 1.842164e-06, 
    1.868689e-06, 1.857243e-06, 1.887154e-06, 1.879977e-06, 1.888876e-06, 
    1.884333e-06, 1.892119e-06, 1.885111e-06, 1.89726e-06, 1.89991e-06, 
    1.898098e-06, 1.905061e-06, 1.884721e-06, 1.89252e-06, 1.834224e-06, 
    1.834564e-06, 1.836151e-06, 1.829179e-06, 1.828753e-06, 1.822378e-06, 
    1.82805e-06, 1.830468e-06, 1.836614e-06, 1.840253e-06, 1.843715e-06, 
    1.851339e-06, 1.859869e-06, 1.871828e-06, 1.880441e-06, 1.886225e-06, 
    1.882678e-06, 1.885809e-06, 1.882308e-06, 1.880668e-06, 1.898916e-06, 
    1.88866e-06, 1.904058e-06, 1.903205e-06, 1.89623e-06, 1.903301e-06, 
    1.834803e-06, 1.832844e-06, 1.826048e-06, 1.831365e-06, 1.821684e-06, 
    1.827099e-06, 1.830216e-06, 1.842268e-06, 1.844921e-06, 1.847382e-06, 
    1.852248e-06, 1.8585e-06, 1.869491e-06, 1.879078e-06, 1.88785e-06, 
    1.887206e-06, 1.887433e-06, 1.889394e-06, 1.884536e-06, 1.890192e-06, 
    1.891141e-06, 1.888658e-06, 1.90309e-06, 1.898962e-06, 1.903186e-06, 
    1.900498e-06, 1.83348e-06, 1.836777e-06, 1.834995e-06, 1.838347e-06, 
    1.835985e-06, 1.846496e-06, 1.849653e-06, 1.864458e-06, 1.858376e-06, 
    1.868061e-06, 1.859359e-06, 1.860899e-06, 1.868375e-06, 1.859829e-06, 
    1.878547e-06, 1.865846e-06, 1.88947e-06, 1.876751e-06, 1.890268e-06, 
    1.887811e-06, 1.89188e-06, 1.895527e-06, 1.900121e-06, 1.90861e-06, 
    1.906643e-06, 1.913752e-06, 1.841698e-06, 1.845984e-06, 1.845607e-06, 
    1.850097e-06, 1.85342e-06, 1.860634e-06, 1.872229e-06, 1.867865e-06, 
    1.875881e-06, 1.877492e-06, 1.865315e-06, 1.872786e-06, 1.848853e-06, 
    1.852709e-06, 1.850414e-06, 1.842033e-06, 1.868868e-06, 1.855074e-06, 
    1.880582e-06, 1.873083e-06, 1.895007e-06, 1.884088e-06, 1.90556e-06, 
    1.91477e-06, 1.923461e-06, 1.933635e-06, 1.848325e-06, 1.845411e-06, 
    1.850631e-06, 1.857863e-06, 1.864586e-06, 1.873541e-06, 1.874459e-06, 
    1.876138e-06, 1.880494e-06, 1.884159e-06, 1.876668e-06, 1.885078e-06, 
    1.853603e-06, 1.870068e-06, 1.844307e-06, 1.852046e-06, 1.857434e-06, 
    1.85507e-06, 1.867365e-06, 1.870267e-06, 1.882083e-06, 1.875972e-06, 
    1.912494e-06, 1.896296e-06, 1.9414e-06, 1.928747e-06, 1.844393e-06, 
    1.848315e-06, 1.861995e-06, 1.85548e-06, 1.87414e-06, 1.878745e-06, 
    1.882493e-06, 1.887289e-06, 1.887807e-06, 1.890651e-06, 1.885991e-06, 
    1.890467e-06, 1.873559e-06, 1.881106e-06, 1.860428e-06, 1.865451e-06, 
    1.863139e-06, 1.860605e-06, 1.868431e-06, 1.876784e-06, 1.876964e-06, 
    1.879646e-06, 1.88721e-06, 1.874213e-06, 1.914586e-06, 1.889604e-06, 
    1.852596e-06, 1.860168e-06, 1.861252e-06, 1.858316e-06, 1.878283e-06, 
    1.871037e-06, 1.890582e-06, 1.885291e-06, 1.893964e-06, 1.889652e-06, 
    1.889017e-06, 1.883486e-06, 1.880046e-06, 1.871367e-06, 1.86432e-06, 
    1.85874e-06, 1.860037e-06, 1.866168e-06, 1.877296e-06, 1.887851e-06, 
    1.885537e-06, 1.893302e-06, 1.872781e-06, 1.881373e-06, 1.878049e-06, 
    1.88672e-06, 1.867748e-06, 1.883897e-06, 1.86363e-06, 1.865403e-06, 
    1.870893e-06, 1.881957e-06, 1.884411e-06, 1.88703e-06, 1.885414e-06, 
    1.87758e-06, 1.876298e-06, 1.870759e-06, 1.86923e-06, 1.865016e-06, 
    1.861529e-06, 1.864714e-06, 1.868061e-06, 1.877583e-06, 1.886182e-06, 
    1.895577e-06, 1.897881e-06, 1.908888e-06, 1.899923e-06, 1.914724e-06, 
    1.902134e-06, 1.923954e-06, 1.884837e-06, 1.90177e-06, 1.871143e-06, 
    1.874432e-06, 1.880386e-06, 1.894077e-06, 1.886682e-06, 1.895332e-06, 
    1.876248e-06, 1.866379e-06, 1.863831e-06, 1.859079e-06, 1.86394e-06, 
    1.863544e-06, 1.8682e-06, 1.866703e-06, 1.877899e-06, 1.871881e-06, 
    1.888999e-06, 1.895263e-06, 1.913004e-06, 1.923916e-06, 1.935055e-06, 
    1.939981e-06, 1.941482e-06, 1.942109e-06 ;

 SMIN_NO3_LEACHED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_RUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_vr =
  8.069541e-06, 8.10375e-06, 8.097082e-06, 8.124684e-06, 8.109367e-06, 
    8.127424e-06, 8.076438e-06, 8.105044e-06, 8.086773e-06, 8.072558e-06, 
    8.17821e-06, 8.12585e-06, 8.23274e-06, 8.199266e-06, 8.283384e-06, 
    8.227498e-06, 8.294656e-06, 8.281766e-06, 8.320574e-06, 8.309439e-06, 
    8.359071e-06, 8.325685e-06, 8.38484e-06, 8.35109e-06, 8.356351e-06, 
    8.32454e-06, 8.136457e-06, 8.171744e-06, 8.134347e-06, 8.139379e-06, 
    8.137115e-06, 8.109641e-06, 8.095795e-06, 8.066861e-06, 8.072102e-06, 
    8.093353e-06, 8.141581e-06, 8.125197e-06, 8.166491e-06, 8.165561e-06, 
    8.211567e-06, 8.190809e-06, 8.268247e-06, 8.246211e-06, 8.309895e-06, 
    8.293853e-06, 8.309122e-06, 8.304479e-06, 8.309157e-06, 8.285656e-06, 
    8.295704e-06, 8.275036e-06, 8.194793e-06, 8.218396e-06, 8.147993e-06, 
    8.105688e-06, 8.077654e-06, 8.057771e-06, 8.060563e-06, 8.06592e-06, 
    8.093461e-06, 8.119384e-06, 8.139154e-06, 8.15237e-06, 8.165402e-06, 
    8.204865e-06, 8.225792e-06, 8.272675e-06, 8.264218e-06, 8.278536e-06, 
    8.29225e-06, 8.315255e-06, 8.311465e-06, 8.321593e-06, 8.278124e-06, 
    8.306998e-06, 8.259327e-06, 8.272355e-06, 8.168975e-06, 8.129654e-06, 
    8.112906e-06, 8.098285e-06, 8.062718e-06, 8.087267e-06, 8.077576e-06, 
    8.100609e-06, 8.115249e-06, 8.107995e-06, 8.152722e-06, 8.135311e-06, 
    8.22702e-06, 8.187489e-06, 8.290661e-06, 8.265935e-06, 8.296563e-06, 
    8.280931e-06, 8.3077e-06, 8.283593e-06, 8.325355e-06, 8.334453e-06, 
    8.328217e-06, 8.352128e-06, 8.282203e-06, 8.309031e-06, 8.10784e-06, 
    8.109022e-06, 8.114517e-06, 8.090303e-06, 8.088823e-06, 8.066664e-06, 
    8.086363e-06, 8.094757e-06, 8.11608e-06, 8.128682e-06, 8.14067e-06, 
    8.167068e-06, 8.196548e-06, 8.237829e-06, 8.267527e-06, 8.287432e-06, 
    8.275218e-06, 8.285984e-06, 8.273928e-06, 8.268269e-06, 8.331016e-06, 
    8.295762e-06, 8.348663e-06, 8.345737e-06, 8.321766e-06, 8.346043e-06, 
    8.109834e-06, 8.103027e-06, 8.079424e-06, 8.097879e-06, 8.064237e-06, 
    8.083052e-06, 8.09386e-06, 8.13565e-06, 8.144843e-06, 8.153364e-06, 
    8.170198e-06, 8.191807e-06, 8.229758e-06, 8.262807e-06, 8.293016e-06, 
    8.290789e-06, 8.291564e-06, 8.298297e-06, 8.281577e-06, 8.301025e-06, 
    8.304276e-06, 8.295742e-06, 8.34532e-06, 8.331148e-06, 8.345641e-06, 
    8.336399e-06, 8.105228e-06, 8.116651e-06, 8.110459e-06, 8.122082e-06, 
    8.113871e-06, 8.150298e-06, 8.161213e-06, 8.212392e-06, 8.191377e-06, 
    8.224826e-06, 8.194761e-06, 8.200083e-06, 8.225865e-06, 8.196367e-06, 
    8.260945e-06, 8.217115e-06, 8.29855e-06, 8.254716e-06, 8.301279e-06, 
    8.292815e-06, 8.306803e-06, 8.319339e-06, 8.335105e-06, 8.36423e-06, 
    8.357468e-06, 8.381847e-06, 8.133703e-06, 8.14853e-06, 8.147231e-06, 
    8.162762e-06, 8.174248e-06, 8.199198e-06, 8.239215e-06, 8.224149e-06, 
    8.25179e-06, 8.257342e-06, 8.21532e-06, 8.241095e-06, 8.158388e-06, 
    8.171712e-06, 8.163775e-06, 8.134738e-06, 8.227531e-06, 8.179859e-06, 
    8.267913e-06, 8.242053e-06, 8.317525e-06, 8.279959e-06, 8.353748e-06, 
    8.385311e-06, 8.415076e-06, 8.449822e-06, 8.156635e-06, 8.146534e-06, 
    8.164598e-06, 8.1896e-06, 8.212824e-06, 8.243729e-06, 8.246887e-06, 
    8.252663e-06, 8.267664e-06, 8.280288e-06, 8.254463e-06, 8.283429e-06, 
    8.174774e-06, 8.231673e-06, 8.1426e-06, 8.169383e-06, 8.188012e-06, 
    8.179844e-06, 8.222321e-06, 8.232324e-06, 8.273037e-06, 8.251988e-06, 
    8.377484e-06, 8.321908e-06, 8.476326e-06, 8.43311e-06, 8.142998e-06, 
    8.156569e-06, 8.203861e-06, 8.18135e-06, 8.245775e-06, 8.261649e-06, 
    8.274547e-06, 8.29105e-06, 8.292821e-06, 8.302604e-06, 8.286557e-06, 
    8.301959e-06, 8.243703e-06, 8.269722e-06, 8.198373e-06, 8.215704e-06, 
    8.207724e-06, 8.198956e-06, 8.225972e-06, 8.25477e-06, 8.255392e-06, 
    8.264615e-06, 8.290614e-06, 8.245879e-06, 8.384597e-06, 8.298829e-06, 
    8.171379e-06, 8.197533e-06, 8.201282e-06, 8.191139e-06, 8.260032e-06, 
    8.23505e-06, 8.302368e-06, 8.284151e-06, 8.313975e-06, 8.299147e-06, 
    8.296946e-06, 8.277914e-06, 8.266044e-06, 8.236124e-06, 8.211781e-06, 
    8.192513e-06, 8.196977e-06, 8.218149e-06, 8.256512e-06, 8.29287e-06, 
    8.28489e-06, 8.3116e-06, 8.240924e-06, 8.270533e-06, 8.259062e-06, 
    8.288935e-06, 8.223709e-06, 8.279344e-06, 8.209486e-06, 8.215596e-06, 
    8.23453e-06, 8.272658e-06, 8.281107e-06, 8.290118e-06, 8.284544e-06, 
    8.257553e-06, 8.25313e-06, 8.234018e-06, 8.228725e-06, 8.214188e-06, 
    8.202127e-06, 8.213126e-06, 8.224657e-06, 8.257505e-06, 8.287107e-06, 
    8.319409e-06, 8.327325e-06, 8.365062e-06, 8.3343e-06, 8.385029e-06, 
    8.341844e-06, 8.416625e-06, 8.282572e-06, 8.340786e-06, 8.235399e-06, 
    8.24673e-06, 8.267233e-06, 8.31433e-06, 8.288898e-06, 8.31864e-06, 
    8.252952e-06, 8.218884e-06, 8.210089e-06, 8.193669e-06, 8.210447e-06, 
    8.209084e-06, 8.22515e-06, 8.21997e-06, 8.258572e-06, 8.237829e-06, 
    8.296774e-06, 8.318309e-06, 8.379187e-06, 8.416529e-06, 8.454613e-06, 
    8.471414e-06, 8.476531e-06, 8.478661e-06,
  5.554614e-06, 5.583951e-06, 5.578247e-06, 5.601928e-06, 5.588793e-06, 
    5.604301e-06, 5.560563e-06, 5.585112e-06, 5.56944e-06, 5.55726e-06, 
    5.647951e-06, 5.602987e-06, 5.694814e-06, 5.666051e-06, 5.738395e-06, 
    5.690329e-06, 5.748103e-06, 5.73702e-06, 5.770426e-06, 5.760851e-06, 
    5.80361e-06, 5.774847e-06, 5.825828e-06, 5.796744e-06, 5.801287e-06, 
    5.773896e-06, 5.612039e-06, 5.642343e-06, 5.610242e-06, 5.614561e-06, 
    5.612625e-06, 5.58906e-06, 5.577187e-06, 5.552381e-06, 5.556885e-06, 
    5.575109e-06, 5.616504e-06, 5.60245e-06, 5.63791e-06, 5.637109e-06, 
    5.676652e-06, 5.658812e-06, 5.725397e-06, 5.706454e-06, 5.761251e-06, 
    5.747455e-06, 5.7606e-06, 5.756615e-06, 5.760652e-06, 5.740423e-06, 
    5.749087e-06, 5.7313e-06, 5.66215e-06, 5.682445e-06, 5.62197e-06, 
    5.585677e-06, 5.561637e-06, 5.544588e-06, 5.546997e-06, 5.551589e-06, 
    5.575216e-06, 5.597466e-06, 5.614437e-06, 5.625795e-06, 5.636994e-06, 
    5.6709e-06, 5.688895e-06, 5.729224e-06, 5.72195e-06, 5.734281e-06, 
    5.746083e-06, 5.765898e-06, 5.762637e-06, 5.771369e-06, 5.733963e-06, 
    5.758812e-06, 5.717806e-06, 5.729012e-06, 5.639999e-06, 5.606242e-06, 
    5.591877e-06, 5.579342e-06, 5.548849e-06, 5.569899e-06, 5.561597e-06, 
    5.581363e-06, 5.593926e-06, 5.587713e-06, 5.626105e-06, 5.611169e-06, 
    5.689962e-06, 5.655986e-06, 5.744706e-06, 5.723444e-06, 5.749807e-06, 
    5.736353e-06, 5.759408e-06, 5.738657e-06, 5.774623e-06, 5.782458e-06, 
    5.777103e-06, 5.797695e-06, 5.737506e-06, 5.760596e-06, 5.587537e-06, 
    5.58855e-06, 5.593275e-06, 5.572515e-06, 5.571248e-06, 5.552256e-06, 
    5.569158e-06, 5.576356e-06, 5.594658e-06, 5.605484e-06, 5.615784e-06, 
    5.638448e-06, 5.663784e-06, 5.699278e-06, 5.724821e-06, 5.741958e-06, 
    5.731451e-06, 5.740727e-06, 5.730356e-06, 5.725499e-06, 5.779519e-06, 
    5.749166e-06, 5.794732e-06, 5.792209e-06, 5.771575e-06, 5.792494e-06, 
    5.589262e-06, 5.583432e-06, 5.563192e-06, 5.57903e-06, 5.55019e-06, 
    5.566323e-06, 5.575603e-06, 5.611472e-06, 5.619372e-06, 5.626687e-06, 
    5.641151e-06, 5.659725e-06, 5.692347e-06, 5.720778e-06, 5.746772e-06, 
    5.744867e-06, 5.745537e-06, 5.751344e-06, 5.736958e-06, 5.753707e-06, 
    5.756515e-06, 5.749167e-06, 5.791871e-06, 5.779663e-06, 5.792156e-06, 
    5.784207e-06, 5.585328e-06, 5.595141e-06, 5.589838e-06, 5.59981e-06, 
    5.592781e-06, 5.624046e-06, 5.63343e-06, 5.677407e-06, 5.659357e-06, 
    5.688103e-06, 5.662278e-06, 5.66685e-06, 5.689024e-06, 5.663676e-06, 
    5.719201e-06, 5.681526e-06, 5.751569e-06, 5.713872e-06, 5.753933e-06, 
    5.746659e-06, 5.758708e-06, 5.7695e-06, 5.783093e-06, 5.808183e-06, 
    5.802372e-06, 5.823378e-06, 5.609784e-06, 5.622525e-06, 5.62141e-06, 
    5.634758e-06, 5.644633e-06, 5.666064e-06, 5.700473e-06, 5.687529e-06, 
    5.711306e-06, 5.71608e-06, 5.679964e-06, 5.702124e-06, 5.631063e-06, 
    5.642519e-06, 5.635703e-06, 5.610784e-06, 5.690501e-06, 5.649546e-06, 
    5.725242e-06, 5.70301e-06, 5.76796e-06, 5.735626e-06, 5.799172e-06, 
    5.826374e-06, 5.852041e-06, 5.882031e-06, 5.629491e-06, 5.620828e-06, 
    5.636348e-06, 5.657826e-06, 5.677797e-06, 5.704364e-06, 5.707088e-06, 
    5.712067e-06, 5.72498e-06, 5.735839e-06, 5.713635e-06, 5.738563e-06, 
    5.645162e-06, 5.694063e-06, 5.617548e-06, 5.640547e-06, 5.656562e-06, 
    5.649543e-06, 5.686052e-06, 5.694664e-06, 5.729691e-06, 5.711581e-06, 
    5.81965e-06, 5.77177e-06, 5.904918e-06, 5.867625e-06, 5.617801e-06, 
    5.629464e-06, 5.6701e-06, 5.650756e-06, 5.706143e-06, 5.719795e-06, 
    5.730907e-06, 5.745107e-06, 5.746646e-06, 5.755066e-06, 5.741269e-06, 
    5.754523e-06, 5.704421e-06, 5.726797e-06, 5.665461e-06, 5.680368e-06, 
    5.673512e-06, 5.665987e-06, 5.689217e-06, 5.713982e-06, 5.714524e-06, 
    5.722469e-06, 5.744852e-06, 5.706368e-06, 5.825814e-06, 5.751948e-06, 
    5.64219e-06, 5.664673e-06, 5.667901e-06, 5.659184e-06, 5.718426e-06, 
    5.69694e-06, 5.754862e-06, 5.739194e-06, 5.764874e-06, 5.752109e-06, 
    5.750231e-06, 5.73385e-06, 5.723655e-06, 5.697922e-06, 5.677011e-06, 
    5.66045e-06, 5.664301e-06, 5.682497e-06, 5.715501e-06, 5.74678e-06, 
    5.739922e-06, 5.762922e-06, 5.702122e-06, 5.727589e-06, 5.717738e-06, 
    5.743435e-06, 5.687183e-06, 5.735038e-06, 5.674964e-06, 5.680226e-06, 
    5.696514e-06, 5.729309e-06, 5.73659e-06, 5.744344e-06, 5.739561e-06, 
    5.716342e-06, 5.712545e-06, 5.69612e-06, 5.691581e-06, 5.679081e-06, 
    5.668732e-06, 5.678185e-06, 5.688114e-06, 5.716357e-06, 5.741835e-06, 
    5.769652e-06, 5.77647e-06, 5.808995e-06, 5.782497e-06, 5.826224e-06, 
    5.789017e-06, 5.853477e-06, 5.737833e-06, 5.787948e-06, 5.697259e-06, 
    5.707013e-06, 5.724655e-06, 5.7652e-06, 5.743314e-06, 5.768917e-06, 
    5.712398e-06, 5.683119e-06, 5.675565e-06, 5.661454e-06, 5.675888e-06, 
    5.674714e-06, 5.688533e-06, 5.684092e-06, 5.717295e-06, 5.699454e-06, 
    5.75018e-06, 5.768718e-06, 5.821171e-06, 5.85338e-06, 5.886233e-06, 
    5.900746e-06, 5.905166e-06, 5.907013e-06,
  6.001858e-06, 6.033908e-06, 6.027676e-06, 6.053554e-06, 6.039197e-06, 
    6.056146e-06, 6.008355e-06, 6.035178e-06, 6.018053e-06, 6.004746e-06, 
    6.103865e-06, 6.05471e-06, 6.155101e-06, 6.123645e-06, 6.202774e-06, 
    6.150198e-06, 6.213394e-06, 6.201265e-06, 6.237818e-06, 6.22734e-06, 
    6.274147e-06, 6.242656e-06, 6.29847e-06, 6.266628e-06, 6.271602e-06, 
    6.241617e-06, 6.064601e-06, 6.097736e-06, 6.062637e-06, 6.067358e-06, 
    6.065241e-06, 6.03949e-06, 6.026521e-06, 5.999416e-06, 6.004336e-06, 
    6.024248e-06, 6.069482e-06, 6.054121e-06, 6.092877e-06, 6.092001e-06, 
    6.135236e-06, 6.115729e-06, 6.188549e-06, 6.167827e-06, 6.227777e-06, 
    6.212682e-06, 6.227066e-06, 6.222705e-06, 6.227123e-06, 6.204989e-06, 
    6.214469e-06, 6.195006e-06, 6.119379e-06, 6.141572e-06, 6.075455e-06, 
    6.0358e-06, 6.009529e-06, 5.990903e-06, 5.993536e-06, 5.998552e-06, 
    6.024365e-06, 6.048675e-06, 6.06722e-06, 6.079634e-06, 6.091875e-06, 
    6.128954e-06, 6.148628e-06, 6.192738e-06, 6.184778e-06, 6.198271e-06, 
    6.211181e-06, 6.232864e-06, 6.229295e-06, 6.238852e-06, 6.197921e-06, 
    6.225112e-06, 6.180243e-06, 6.192504e-06, 6.095174e-06, 6.058265e-06, 
    6.042573e-06, 6.028872e-06, 5.995559e-06, 6.018556e-06, 6.009486e-06, 
    6.031078e-06, 6.044806e-06, 6.038017e-06, 6.079973e-06, 6.063649e-06, 
    6.149794e-06, 6.112641e-06, 6.209675e-06, 6.186412e-06, 6.215256e-06, 
    6.200534e-06, 6.225763e-06, 6.203056e-06, 6.242413e-06, 6.250989e-06, 
    6.245127e-06, 6.267666e-06, 6.201797e-06, 6.227063e-06, 6.037825e-06, 
    6.038932e-06, 6.044093e-06, 6.021414e-06, 6.020029e-06, 5.99928e-06, 
    6.017744e-06, 6.02561e-06, 6.045605e-06, 6.057437e-06, 6.068693e-06, 
    6.093467e-06, 6.121168e-06, 6.159981e-06, 6.187919e-06, 6.206667e-06, 
    6.195171e-06, 6.20532e-06, 6.193974e-06, 6.188659e-06, 6.247773e-06, 
    6.214555e-06, 6.264423e-06, 6.261661e-06, 6.239079e-06, 6.261972e-06, 
    6.03971e-06, 6.033339e-06, 6.011227e-06, 6.028529e-06, 5.997023e-06, 
    6.014648e-06, 6.024788e-06, 6.063984e-06, 6.072614e-06, 6.08061e-06, 
    6.096421e-06, 6.116727e-06, 6.152401e-06, 6.183497e-06, 6.211933e-06, 
    6.209849e-06, 6.210583e-06, 6.216937e-06, 6.201196e-06, 6.219523e-06, 
    6.222597e-06, 6.214555e-06, 6.261291e-06, 6.247928e-06, 6.261602e-06, 
    6.252902e-06, 6.03541e-06, 6.046134e-06, 6.040338e-06, 6.051237e-06, 
    6.043556e-06, 6.077727e-06, 6.087985e-06, 6.136066e-06, 6.116325e-06, 
    6.147759e-06, 6.119518e-06, 6.124519e-06, 6.148773e-06, 6.121046e-06, 
    6.181775e-06, 6.140571e-06, 6.217184e-06, 6.175949e-06, 6.219771e-06, 
    6.211811e-06, 6.224995e-06, 6.236806e-06, 6.251682e-06, 6.27915e-06, 
    6.272788e-06, 6.295785e-06, 6.062136e-06, 6.076063e-06, 6.074842e-06, 
    6.089432e-06, 6.100228e-06, 6.123657e-06, 6.161286e-06, 6.147129e-06, 
    6.173134e-06, 6.178356e-06, 6.138856e-06, 6.163094e-06, 6.085394e-06, 
    6.09792e-06, 6.090465e-06, 6.063231e-06, 6.150382e-06, 6.105602e-06, 
    6.18838e-06, 6.164061e-06, 6.235121e-06, 6.199743e-06, 6.269285e-06, 
    6.299072e-06, 6.327173e-06, 6.36003e-06, 6.083675e-06, 6.074206e-06, 
    6.091169e-06, 6.114654e-06, 6.136488e-06, 6.165542e-06, 6.168521e-06, 
    6.173968e-06, 6.188092e-06, 6.199973e-06, 6.175685e-06, 6.202952e-06, 
    6.100815e-06, 6.154277e-06, 6.070622e-06, 6.095765e-06, 6.113271e-06, 
    6.105596e-06, 6.145513e-06, 6.154931e-06, 6.193248e-06, 6.173434e-06, 
    6.29171e-06, 6.239294e-06, 6.385103e-06, 6.344247e-06, 6.070897e-06, 
    6.083645e-06, 6.128073e-06, 6.106922e-06, 6.167487e-06, 6.182421e-06, 
    6.194576e-06, 6.210114e-06, 6.211797e-06, 6.22101e-06, 6.205913e-06, 
    6.220416e-06, 6.165605e-06, 6.19008e-06, 6.122997e-06, 6.139299e-06, 
    6.1318e-06, 6.123572e-06, 6.148975e-06, 6.176066e-06, 6.176655e-06, 
    6.185348e-06, 6.20985e-06, 6.167733e-06, 6.298468e-06, 6.217611e-06, 
    6.097556e-06, 6.122141e-06, 6.125667e-06, 6.116135e-06, 6.180923e-06, 
    6.157422e-06, 6.220787e-06, 6.203643e-06, 6.231743e-06, 6.217774e-06, 
    6.215719e-06, 6.197796e-06, 6.186644e-06, 6.158497e-06, 6.135629e-06, 
    6.117518e-06, 6.121729e-06, 6.141628e-06, 6.177726e-06, 6.211944e-06, 
    6.204443e-06, 6.229606e-06, 6.163089e-06, 6.190948e-06, 6.180173e-06, 
    6.208284e-06, 6.146751e-06, 6.199109e-06, 6.133388e-06, 6.139143e-06, 
    6.156956e-06, 6.192833e-06, 6.200793e-06, 6.209279e-06, 6.204044e-06, 
    6.178645e-06, 6.174491e-06, 6.156525e-06, 6.151563e-06, 6.137891e-06, 
    6.126574e-06, 6.136911e-06, 6.14777e-06, 6.17866e-06, 6.206534e-06, 
    6.236973e-06, 6.244433e-06, 6.280047e-06, 6.251038e-06, 6.298917e-06, 
    6.258185e-06, 6.328758e-06, 6.202162e-06, 6.257006e-06, 6.15777e-06, 
    6.168439e-06, 6.187741e-06, 6.232104e-06, 6.208152e-06, 6.236172e-06, 
    6.174329e-06, 6.14231e-06, 6.134046e-06, 6.118617e-06, 6.134399e-06, 
    6.133115e-06, 6.148226e-06, 6.14337e-06, 6.179686e-06, 6.160171e-06, 
    6.215665e-06, 6.235953e-06, 6.29337e-06, 6.328644e-06, 6.364628e-06, 
    6.380529e-06, 6.385372e-06, 6.387396e-06,
  6.365673e-06, 6.400292e-06, 6.393558e-06, 6.421522e-06, 6.406005e-06, 
    6.424325e-06, 6.372687e-06, 6.401667e-06, 6.383162e-06, 6.368789e-06, 
    6.47593e-06, 6.422772e-06, 6.531359e-06, 6.497314e-06, 6.582981e-06, 
    6.526055e-06, 6.594486e-06, 6.581342e-06, 6.620947e-06, 6.609591e-06, 
    6.660345e-06, 6.626191e-06, 6.686724e-06, 6.652185e-06, 6.657581e-06, 
    6.625065e-06, 6.43346e-06, 6.469301e-06, 6.431338e-06, 6.436444e-06, 
    6.434153e-06, 6.406324e-06, 6.392316e-06, 6.363033e-06, 6.368346e-06, 
    6.389857e-06, 6.43874e-06, 6.422132e-06, 6.46403e-06, 6.463083e-06, 
    6.509854e-06, 6.488749e-06, 6.567569e-06, 6.545129e-06, 6.610065e-06, 
    6.593709e-06, 6.609296e-06, 6.604569e-06, 6.609358e-06, 6.585377e-06, 
    6.595646e-06, 6.574562e-06, 6.492698e-06, 6.516712e-06, 6.445196e-06, 
    6.402343e-06, 6.373956e-06, 6.353841e-06, 6.356683e-06, 6.362102e-06, 
    6.389983e-06, 6.416246e-06, 6.43629e-06, 6.449711e-06, 6.462947e-06, 
    6.503067e-06, 6.524353e-06, 6.572108e-06, 6.563484e-06, 6.578101e-06, 
    6.592084e-06, 6.61558e-06, 6.611711e-06, 6.62207e-06, 6.577719e-06, 
    6.60718e-06, 6.558572e-06, 6.571851e-06, 6.466531e-06, 6.426612e-06, 
    6.409661e-06, 6.394851e-06, 6.358869e-06, 6.383707e-06, 6.373911e-06, 
    6.397232e-06, 6.412066e-06, 6.404729e-06, 6.450078e-06, 6.432431e-06, 
    6.525615e-06, 6.48541e-06, 6.590451e-06, 6.565254e-06, 6.596497e-06, 
    6.580548e-06, 6.607885e-06, 6.58328e-06, 6.625929e-06, 6.635229e-06, 
    6.628873e-06, 6.653307e-06, 6.581917e-06, 6.609294e-06, 6.404522e-06, 
    6.405719e-06, 6.411295e-06, 6.386795e-06, 6.385298e-06, 6.362887e-06, 
    6.382828e-06, 6.391327e-06, 6.412928e-06, 6.425716e-06, 6.437884e-06, 
    6.464669e-06, 6.494636e-06, 6.536639e-06, 6.566886e-06, 6.587192e-06, 
    6.574739e-06, 6.585733e-06, 6.573443e-06, 6.567686e-06, 6.631742e-06, 
    6.595742e-06, 6.649791e-06, 6.646796e-06, 6.622317e-06, 6.647133e-06, 
    6.406559e-06, 6.399674e-06, 6.37579e-06, 6.394478e-06, 6.360448e-06, 
    6.379486e-06, 6.390442e-06, 6.432796e-06, 6.442122e-06, 6.450768e-06, 
    6.467863e-06, 6.489828e-06, 6.528433e-06, 6.562099e-06, 6.592898e-06, 
    6.590639e-06, 6.591434e-06, 6.59832e-06, 6.581267e-06, 6.601122e-06, 
    6.604455e-06, 6.595739e-06, 6.646394e-06, 6.631907e-06, 6.646732e-06, 
    6.637298e-06, 6.401912e-06, 6.413501e-06, 6.407237e-06, 6.419016e-06, 
    6.410716e-06, 6.447654e-06, 6.458747e-06, 6.510757e-06, 6.489395e-06, 
    6.52341e-06, 6.492848e-06, 6.498258e-06, 6.524514e-06, 6.494499e-06, 
    6.560238e-06, 6.515634e-06, 6.598587e-06, 6.553933e-06, 6.60139e-06, 
    6.592764e-06, 6.60705e-06, 6.619853e-06, 6.635977e-06, 6.665765e-06, 
    6.658863e-06, 6.683808e-06, 6.430794e-06, 6.445853e-06, 6.44453e-06, 
    6.460305e-06, 6.471982e-06, 6.497324e-06, 6.53805e-06, 6.522724e-06, 
    6.550874e-06, 6.55653e-06, 6.513769e-06, 6.540008e-06, 6.455942e-06, 
    6.469491e-06, 6.461425e-06, 6.431981e-06, 6.52625e-06, 6.477799e-06, 
    6.567386e-06, 6.541053e-06, 6.618026e-06, 6.579698e-06, 6.655064e-06, 
    6.687381e-06, 6.717869e-06, 6.753552e-06, 6.454081e-06, 6.443842e-06, 
    6.462184e-06, 6.48759e-06, 6.511209e-06, 6.542657e-06, 6.54588e-06, 
    6.551779e-06, 6.567072e-06, 6.57994e-06, 6.553642e-06, 6.583168e-06, 
    6.47263e-06, 6.530463e-06, 6.43997e-06, 6.467161e-06, 6.486092e-06, 
    6.477788e-06, 6.520974e-06, 6.531168e-06, 6.57266e-06, 6.5512e-06, 
    6.679396e-06, 6.622554e-06, 6.780782e-06, 6.736411e-06, 6.440265e-06, 
    6.454047e-06, 6.502105e-06, 6.479222e-06, 6.54476e-06, 6.560932e-06, 
    6.574094e-06, 6.590929e-06, 6.59275e-06, 6.602734e-06, 6.586376e-06, 
    6.602088e-06, 6.542724e-06, 6.569226e-06, 6.496609e-06, 6.514251e-06, 
    6.506134e-06, 6.497232e-06, 6.524721e-06, 6.554054e-06, 6.554686e-06, 
    6.564103e-06, 6.59066e-06, 6.545027e-06, 6.686738e-06, 6.599068e-06, 
    6.46909e-06, 6.495691e-06, 6.499499e-06, 6.489186e-06, 6.55931e-06, 
    6.533866e-06, 6.602491e-06, 6.583917e-06, 6.614363e-06, 6.599226e-06, 
    6.597e-06, 6.577583e-06, 6.565504e-06, 6.535031e-06, 6.510279e-06, 
    6.490682e-06, 6.495238e-06, 6.516772e-06, 6.555852e-06, 6.592912e-06, 
    6.584787e-06, 6.612047e-06, 6.54e-06, 6.570169e-06, 6.5585e-06, 
    6.588944e-06, 6.522316e-06, 6.579022e-06, 6.507852e-06, 6.51408e-06, 
    6.533362e-06, 6.572214e-06, 6.58083e-06, 6.590025e-06, 6.584351e-06, 
    6.556846e-06, 6.552346e-06, 6.532894e-06, 6.527524e-06, 6.512724e-06, 
    6.500479e-06, 6.511666e-06, 6.523421e-06, 6.556859e-06, 6.587051e-06, 
    6.620034e-06, 6.628118e-06, 6.666747e-06, 6.635288e-06, 6.687227e-06, 
    6.64305e-06, 6.719604e-06, 6.582322e-06, 6.64176e-06, 6.534241e-06, 
    6.545791e-06, 6.566699e-06, 6.614762e-06, 6.588802e-06, 6.619169e-06, 
    6.55217e-06, 6.517514e-06, 6.508565e-06, 6.491872e-06, 6.508947e-06, 
    6.507557e-06, 6.523911e-06, 6.518654e-06, 6.557971e-06, 6.53684e-06, 
    6.596943e-06, 6.618931e-06, 6.681191e-06, 6.719471e-06, 6.758537e-06, 
    6.775811e-06, 6.781072e-06, 6.783273e-06,
  6.298839e-06, 6.334344e-06, 6.327433e-06, 6.356134e-06, 6.340204e-06, 
    6.35901e-06, 6.306028e-06, 6.335755e-06, 6.316769e-06, 6.302031e-06, 
    6.412042e-06, 6.357417e-06, 6.469063e-06, 6.43402e-06, 6.522257e-06, 
    6.463604e-06, 6.534121e-06, 6.520561e-06, 6.561421e-06, 6.549701e-06, 
    6.602123e-06, 6.566835e-06, 6.629391e-06, 6.593686e-06, 6.599264e-06, 
    6.565673e-06, 6.368388e-06, 6.405226e-06, 6.366209e-06, 6.371454e-06, 
    6.3691e-06, 6.340533e-06, 6.326164e-06, 6.29613e-06, 6.301576e-06, 
    6.323638e-06, 6.373813e-06, 6.356756e-06, 6.399793e-06, 6.39882e-06, 
    6.446922e-06, 6.425209e-06, 6.506363e-06, 6.483239e-06, 6.550189e-06, 
    6.533316e-06, 6.549396e-06, 6.544518e-06, 6.54946e-06, 6.524722e-06, 
    6.535314e-06, 6.51357e-06, 6.429272e-06, 6.453982e-06, 6.380443e-06, 
    6.336455e-06, 6.30733e-06, 6.286709e-06, 6.289622e-06, 6.295177e-06, 
    6.323768e-06, 6.350714e-06, 6.371293e-06, 6.385079e-06, 6.39868e-06, 
    6.439947e-06, 6.46185e-06, 6.511045e-06, 6.502151e-06, 6.517222e-06, 
    6.531638e-06, 6.555882e-06, 6.551888e-06, 6.562582e-06, 6.516824e-06, 
    6.547215e-06, 6.497088e-06, 6.510777e-06, 6.402381e-06, 6.361355e-06, 
    6.343963e-06, 6.328761e-06, 6.291863e-06, 6.317331e-06, 6.307284e-06, 
    6.3312e-06, 6.346424e-06, 6.338892e-06, 6.385456e-06, 6.367331e-06, 
    6.463149e-06, 6.421778e-06, 6.529955e-06, 6.503976e-06, 6.536191e-06, 
    6.519741e-06, 6.547942e-06, 6.522559e-06, 6.566565e-06, 6.57617e-06, 
    6.569605e-06, 6.594842e-06, 6.521153e-06, 6.549396e-06, 6.338681e-06, 
    6.339909e-06, 6.345631e-06, 6.320498e-06, 6.318961e-06, 6.295981e-06, 
    6.316427e-06, 6.325145e-06, 6.347307e-06, 6.360436e-06, 6.372931e-06, 
    6.400452e-06, 6.431268e-06, 6.474498e-06, 6.505658e-06, 6.526593e-06, 
    6.513751e-06, 6.525088e-06, 6.512416e-06, 6.506481e-06, 6.57257e-06, 
    6.535414e-06, 6.591209e-06, 6.588115e-06, 6.562837e-06, 6.588463e-06, 
    6.340772e-06, 6.333706e-06, 6.30921e-06, 6.328376e-06, 6.293481e-06, 
    6.313e-06, 6.324239e-06, 6.367709e-06, 6.377283e-06, 6.386167e-06, 
    6.403734e-06, 6.426319e-06, 6.466048e-06, 6.500727e-06, 6.532477e-06, 
    6.530147e-06, 6.530968e-06, 6.538072e-06, 6.520483e-06, 6.540962e-06, 
    6.544403e-06, 6.535409e-06, 6.5877e-06, 6.572737e-06, 6.588049e-06, 
    6.578304e-06, 6.336002e-06, 6.347896e-06, 6.341467e-06, 6.353559e-06, 
    6.345039e-06, 6.382972e-06, 6.39437e-06, 6.447855e-06, 6.425874e-06, 
    6.460877e-06, 6.429425e-06, 6.434992e-06, 6.462021e-06, 6.431123e-06, 
    6.498812e-06, 6.452877e-06, 6.538348e-06, 6.492319e-06, 6.541239e-06, 
    6.53234e-06, 6.547077e-06, 6.560293e-06, 6.57694e-06, 6.60772e-06, 
    6.600585e-06, 6.626373e-06, 6.36565e-06, 6.381119e-06, 6.379757e-06, 
    6.395966e-06, 6.407969e-06, 6.434028e-06, 6.475949e-06, 6.460167e-06, 
    6.489157e-06, 6.494986e-06, 6.45095e-06, 6.477967e-06, 6.391484e-06, 
    6.405412e-06, 6.397117e-06, 6.36687e-06, 6.463802e-06, 6.413953e-06, 
    6.506174e-06, 6.479042e-06, 6.558407e-06, 6.518869e-06, 6.59666e-06, 
    6.630076e-06, 6.661614e-06, 6.698581e-06, 6.389571e-06, 6.379049e-06, 
    6.397896e-06, 6.424021e-06, 6.448316e-06, 6.480694e-06, 6.484012e-06, 
    6.490091e-06, 6.505848e-06, 6.519115e-06, 6.492013e-06, 6.522443e-06, 
    6.408646e-06, 6.468139e-06, 6.375075e-06, 6.403018e-06, 6.42248e-06, 
    6.413938e-06, 6.458365e-06, 6.468861e-06, 6.511613e-06, 6.489493e-06, 
    6.621819e-06, 6.563087e-06, 6.726806e-06, 6.68082e-06, 6.375376e-06, 
    6.389535e-06, 6.438951e-06, 6.415412e-06, 6.482859e-06, 6.499522e-06, 
    6.513087e-06, 6.530449e-06, 6.532325e-06, 6.542627e-06, 6.525751e-06, 
    6.541959e-06, 6.480764e-06, 6.50807e-06, 6.433292e-06, 6.451447e-06, 
    6.443091e-06, 6.433933e-06, 6.462223e-06, 6.492439e-06, 6.493085e-06, 
    6.502792e-06, 6.530189e-06, 6.483134e-06, 6.629422e-06, 6.538859e-06, 
    6.404995e-06, 6.432354e-06, 6.436267e-06, 6.425657e-06, 6.497851e-06, 
    6.47164e-06, 6.542375e-06, 6.523215e-06, 6.554626e-06, 6.539006e-06, 
    6.53671e-06, 6.516685e-06, 6.504234e-06, 6.472841e-06, 6.44736e-06, 
    6.427195e-06, 6.431882e-06, 6.454043e-06, 6.49429e-06, 6.532495e-06, 
    6.524116e-06, 6.552235e-06, 6.477956e-06, 6.509044e-06, 6.497019e-06, 
    6.528401e-06, 6.459748e-06, 6.518184e-06, 6.444859e-06, 6.451269e-06, 
    6.47112e-06, 6.511155e-06, 6.520032e-06, 6.529517e-06, 6.523663e-06, 
    6.495314e-06, 6.490675e-06, 6.470637e-06, 6.465111e-06, 6.449873e-06, 
    6.437273e-06, 6.448785e-06, 6.460887e-06, 6.495325e-06, 6.52645e-06, 
    6.56048e-06, 6.568825e-06, 6.608744e-06, 6.576238e-06, 6.629929e-06, 
    6.584267e-06, 6.663426e-06, 6.52158e-06, 6.582925e-06, 6.472024e-06, 
    6.48392e-06, 6.505469e-06, 6.555044e-06, 6.528253e-06, 6.559591e-06, 
    6.490494e-06, 6.454808e-06, 6.445593e-06, 6.42842e-06, 6.445986e-06, 
    6.444556e-06, 6.461388e-06, 6.455976e-06, 6.496471e-06, 6.474701e-06, 
    6.536653e-06, 6.559344e-06, 6.623668e-06, 6.663279e-06, 6.70374e-06, 
    6.721649e-06, 6.727105e-06, 6.729387e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOINTABS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWDP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWLIQ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_DEPTH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SINKS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SOURCES =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1C =
  5.777232, 5.777217, 5.77722, 5.777209, 5.777215, 5.777207, 5.777229, 
    5.777217, 5.777225, 5.777231, 5.777186, 5.777208, 5.777163, 5.777177, 
    5.777141, 5.777165, 5.777136, 5.777142, 5.777125, 5.77713, 5.777109, 
    5.777123, 5.777098, 5.777112, 5.77711, 5.777123, 5.777204, 5.777189, 
    5.777205, 5.777202, 5.777203, 5.777215, 5.777221, 5.777233, 5.777231, 
    5.777222, 5.777201, 5.777208, 5.777191, 5.777191, 5.777172, 5.77718, 
    5.777147, 5.777157, 5.77713, 5.777136, 5.77713, 5.777132, 5.77713, 
    5.77714, 5.777136, 5.777144, 5.777179, 5.777169, 5.777199, 5.777217, 
    5.777229, 5.777237, 5.777236, 5.777234, 5.777222, 5.777211, 5.777203, 
    5.777197, 5.777191, 5.777174, 5.777165, 5.777145, 5.777149, 5.777143, 
    5.777137, 5.777127, 5.777129, 5.777125, 5.777143, 5.777131, 5.777151, 
    5.777146, 5.77719, 5.777206, 5.777214, 5.77722, 5.777235, 5.777225, 
    5.777229, 5.777219, 5.777213, 5.777215, 5.777196, 5.777204, 5.777165, 
    5.777182, 5.777138, 5.777148, 5.777135, 5.777142, 5.777131, 5.777141, 
    5.777123, 5.777119, 5.777122, 5.777112, 5.777142, 5.77713, 5.777216, 
    5.777215, 5.777213, 5.777223, 5.777224, 5.777234, 5.777225, 5.777221, 
    5.777212, 5.777207, 5.777202, 5.777191, 5.777178, 5.77716, 5.777148, 
    5.777139, 5.777144, 5.77714, 5.777145, 5.777147, 5.777121, 5.777136, 
    5.777113, 5.777114, 5.777125, 5.777114, 5.777215, 5.777218, 5.777228, 
    5.77722, 5.777235, 5.777226, 5.777222, 5.777204, 5.7772, 5.777196, 
    5.777189, 5.77718, 5.777164, 5.77715, 5.777137, 5.777138, 5.777137, 
    5.777134, 5.777142, 5.777133, 5.777132, 5.777136, 5.777115, 5.777121, 
    5.777114, 5.777119, 5.777217, 5.777212, 5.777215, 5.77721, 5.777213, 
    5.777198, 5.777193, 5.777171, 5.77718, 5.777166, 5.777179, 5.777176, 
    5.777165, 5.777178, 5.777151, 5.777169, 5.777134, 5.777153, 5.777133, 
    5.777137, 5.777131, 5.777126, 5.777119, 5.777107, 5.77711, 5.777099, 
    5.777205, 5.777198, 5.777199, 5.777192, 5.777187, 5.777177, 5.77716, 
    5.777166, 5.777154, 5.777152, 5.77717, 5.777159, 5.777194, 5.777188, 
    5.777192, 5.777204, 5.777164, 5.777185, 5.777147, 5.777159, 5.777126, 
    5.777143, 5.777111, 5.777098, 5.777085, 5.777071, 5.777195, 5.777199, 
    5.777192, 5.777181, 5.777171, 5.777158, 5.777156, 5.777154, 5.777148, 
    5.777143, 5.777153, 5.777141, 5.777187, 5.777163, 5.777201, 5.777189, 
    5.777182, 5.777185, 5.777167, 5.777163, 5.777145, 5.777154, 5.777101, 
    5.777124, 5.777059, 5.777078, 5.777201, 5.777195, 5.777175, 5.777184, 
    5.777157, 5.77715, 5.777145, 5.777138, 5.777137, 5.777133, 5.77714, 
    5.777133, 5.777158, 5.777147, 5.777177, 5.77717, 5.777173, 5.777177, 
    5.777165, 5.777153, 5.777153, 5.777149, 5.777138, 5.777157, 5.777098, 
    5.777134, 5.777189, 5.777177, 5.777176, 5.77718, 5.777151, 5.777162, 
    5.777133, 5.777141, 5.777128, 5.777134, 5.777135, 5.777143, 5.777148, 
    5.777161, 5.777171, 5.77718, 5.777178, 5.777169, 5.777153, 5.777137, 
    5.77714, 5.777129, 5.777159, 5.777146, 5.777151, 5.777139, 5.777166, 
    5.777143, 5.777173, 5.77717, 5.777162, 5.777145, 5.777142, 5.777138, 
    5.777141, 5.777152, 5.777154, 5.777162, 5.777164, 5.77717, 5.777175, 
    5.777171, 5.777166, 5.777152, 5.777139, 5.777126, 5.777122, 5.777106, 
    5.777119, 5.777098, 5.777116, 5.777084, 5.777141, 5.777117, 5.777161, 
    5.777156, 5.777148, 5.777128, 5.777139, 5.777126, 5.777154, 5.777168, 
    5.777172, 5.777179, 5.777172, 5.777173, 5.777166, 5.777168, 5.777152, 
    5.77716, 5.777135, 5.777126, 5.7771, 5.777084, 5.777069, 5.777061, 
    5.777059, 5.777058 ;

 SOIL1C_TO_SOIL2C =
  3.814669e-08, 3.825103e-08, 3.823075e-08, 3.831488e-08, 3.826822e-08, 
    3.83233e-08, 3.816785e-08, 3.825516e-08, 3.819943e-08, 3.815609e-08, 
    3.847808e-08, 3.831864e-08, 3.864371e-08, 3.854206e-08, 3.879737e-08, 
    3.862788e-08, 3.883154e-08, 3.87925e-08, 3.891003e-08, 3.887637e-08, 
    3.902662e-08, 3.892557e-08, 3.910451e-08, 3.90025e-08, 3.901845e-08, 
    3.892223e-08, 3.835075e-08, 3.845823e-08, 3.834437e-08, 3.83597e-08, 
    3.835283e-08, 3.826918e-08, 3.822701e-08, 3.813872e-08, 3.815475e-08, 
    3.82196e-08, 3.83666e-08, 3.831672e-08, 3.844245e-08, 3.843961e-08, 
    3.857953e-08, 3.851645e-08, 3.875155e-08, 3.868475e-08, 3.887777e-08, 
    3.882923e-08, 3.887549e-08, 3.886147e-08, 3.887567e-08, 3.880449e-08, 
    3.883499e-08, 3.877235e-08, 3.852826e-08, 3.860001e-08, 3.838597e-08, 
    3.82572e-08, 3.817168e-08, 3.811097e-08, 3.811955e-08, 3.813591e-08, 
    3.821998e-08, 3.829902e-08, 3.835925e-08, 3.839952e-08, 3.843921e-08, 
    3.855925e-08, 3.862281e-08, 3.876505e-08, 3.87394e-08, 3.878286e-08, 
    3.882441e-08, 3.889412e-08, 3.888265e-08, 3.891336e-08, 3.878173e-08, 
    3.886921e-08, 3.872479e-08, 3.876429e-08, 3.844993e-08, 3.833018e-08, 
    3.827922e-08, 3.823465e-08, 3.812615e-08, 3.820107e-08, 3.817154e-08, 
    3.824182e-08, 3.828645e-08, 3.826438e-08, 3.840062e-08, 3.834766e-08, 
    3.862657e-08, 3.850646e-08, 3.881956e-08, 3.874467e-08, 3.883751e-08, 
    3.879014e-08, 3.88713e-08, 3.879826e-08, 3.892479e-08, 3.895233e-08, 
    3.893351e-08, 3.900582e-08, 3.879421e-08, 3.887548e-08, 3.826376e-08, 
    3.826736e-08, 3.828413e-08, 3.821038e-08, 3.820587e-08, 3.813828e-08, 
    3.819843e-08, 3.822403e-08, 3.828905e-08, 3.832749e-08, 3.836403e-08, 
    3.844437e-08, 3.853405e-08, 3.865945e-08, 3.874952e-08, 3.880988e-08, 
    3.877287e-08, 3.880555e-08, 3.876902e-08, 3.87519e-08, 3.894201e-08, 
    3.883527e-08, 3.899542e-08, 3.898656e-08, 3.891408e-08, 3.898756e-08, 
    3.826989e-08, 3.824917e-08, 3.817721e-08, 3.823352e-08, 3.813092e-08, 
    3.818835e-08, 3.822137e-08, 3.834876e-08, 3.837675e-08, 3.840269e-08, 
    3.845393e-08, 3.851968e-08, 3.863498e-08, 3.873528e-08, 3.882683e-08, 
    3.882012e-08, 3.882248e-08, 3.884292e-08, 3.879228e-08, 3.885124e-08, 
    3.886113e-08, 3.883526e-08, 3.898537e-08, 3.89425e-08, 3.898637e-08, 
    3.895846e-08, 3.825591e-08, 3.829077e-08, 3.827193e-08, 3.830735e-08, 
    3.828239e-08, 3.839335e-08, 3.842661e-08, 3.858222e-08, 3.851838e-08, 
    3.862e-08, 3.852871e-08, 3.854489e-08, 3.862329e-08, 3.853365e-08, 
    3.872974e-08, 3.859679e-08, 3.884372e-08, 3.871097e-08, 3.885203e-08, 
    3.882643e-08, 3.886883e-08, 3.890678e-08, 3.895455e-08, 3.904264e-08, 
    3.902224e-08, 3.909591e-08, 3.834274e-08, 3.838795e-08, 3.838398e-08, 
    3.843129e-08, 3.846627e-08, 3.854209e-08, 3.866366e-08, 3.861795e-08, 
    3.870187e-08, 3.871871e-08, 3.859122e-08, 3.866949e-08, 3.841821e-08, 
    3.845881e-08, 3.843464e-08, 3.834631e-08, 3.862847e-08, 3.848368e-08, 
    3.875101e-08, 3.867261e-08, 3.890137e-08, 3.878761e-08, 3.901101e-08, 
    3.910644e-08, 3.919629e-08, 3.93012e-08, 3.841263e-08, 3.838192e-08, 
    3.843692e-08, 3.851298e-08, 3.858358e-08, 3.867739e-08, 3.868699e-08, 
    3.870456e-08, 3.875008e-08, 3.878834e-08, 3.871011e-08, 3.879792e-08, 
    3.84682e-08, 3.864104e-08, 3.83703e-08, 3.845183e-08, 3.85085e-08, 
    3.848365e-08, 3.861273e-08, 3.864314e-08, 3.876669e-08, 3.870284e-08, 
    3.908288e-08, 3.891479e-08, 3.938109e-08, 3.925083e-08, 3.837118e-08, 
    3.841253e-08, 3.855638e-08, 3.848794e-08, 3.868366e-08, 3.873181e-08, 
    3.877096e-08, 3.882098e-08, 3.882639e-08, 3.885602e-08, 3.880746e-08, 
    3.885411e-08, 3.867759e-08, 3.875648e-08, 3.853996e-08, 3.859266e-08, 
    3.856842e-08, 3.854182e-08, 3.862391e-08, 3.871133e-08, 3.871322e-08, 
    3.874124e-08, 3.882017e-08, 3.868445e-08, 3.910454e-08, 3.884513e-08, 
    3.845761e-08, 3.853721e-08, 3.85486e-08, 3.851776e-08, 3.872698e-08, 
    3.865118e-08, 3.88553e-08, 3.880015e-08, 3.889051e-08, 3.884561e-08, 
    3.8839e-08, 3.878133e-08, 3.874541e-08, 3.865466e-08, 3.85808e-08, 
    3.852223e-08, 3.853586e-08, 3.860019e-08, 3.871668e-08, 3.882687e-08, 
    3.880273e-08, 3.888365e-08, 3.866947e-08, 3.875929e-08, 3.872457e-08, 
    3.881509e-08, 3.861674e-08, 3.87856e-08, 3.857355e-08, 3.859215e-08, 
    3.864968e-08, 3.876536e-08, 3.879098e-08, 3.881829e-08, 3.880144e-08, 
    3.871964e-08, 3.870625e-08, 3.864828e-08, 3.863227e-08, 3.858811e-08, 
    3.855153e-08, 3.858494e-08, 3.862003e-08, 3.871968e-08, 3.880946e-08, 
    3.890732e-08, 3.893128e-08, 3.904553e-08, 3.89525e-08, 3.910598e-08, 
    3.897546e-08, 3.920139e-08, 3.879541e-08, 3.897166e-08, 3.86523e-08, 
    3.868672e-08, 3.874896e-08, 3.889169e-08, 3.881466e-08, 3.890475e-08, 
    3.870572e-08, 3.86024e-08, 3.857568e-08, 3.852579e-08, 3.857682e-08, 
    3.857267e-08, 3.862149e-08, 3.860581e-08, 3.872299e-08, 3.866005e-08, 
    3.883883e-08, 3.890405e-08, 3.908818e-08, 3.9201e-08, 3.931584e-08, 
    3.936652e-08, 3.938194e-08, 3.938839e-08 ;

 SOIL1C_TO_SOIL3C =
  4.523851e-10, 4.536231e-10, 4.533825e-10, 4.543807e-10, 4.538271e-10, 
    4.544806e-10, 4.526362e-10, 4.536721e-10, 4.530109e-10, 4.524967e-10, 
    4.56317e-10, 4.544253e-10, 4.582821e-10, 4.570761e-10, 4.601054e-10, 
    4.580944e-10, 4.605108e-10, 4.600476e-10, 4.614421e-10, 4.610427e-10, 
    4.628255e-10, 4.616265e-10, 4.637497e-10, 4.625393e-10, 4.627286e-10, 
    4.615869e-10, 4.548062e-10, 4.560815e-10, 4.547306e-10, 4.549125e-10, 
    4.548309e-10, 4.538384e-10, 4.533381e-10, 4.522906e-10, 4.524808e-10, 
    4.532502e-10, 4.549943e-10, 4.544025e-10, 4.558942e-10, 4.558606e-10, 
    4.575207e-10, 4.567723e-10, 4.595617e-10, 4.587692e-10, 4.610594e-10, 
    4.604835e-10, 4.610323e-10, 4.608659e-10, 4.610344e-10, 4.601898e-10, 
    4.605517e-10, 4.598085e-10, 4.569124e-10, 4.577636e-10, 4.552242e-10, 
    4.536963e-10, 4.526816e-10, 4.519613e-10, 4.520631e-10, 4.522572e-10, 
    4.532547e-10, 4.541925e-10, 4.549071e-10, 4.553849e-10, 4.558557e-10, 
    4.5728e-10, 4.580342e-10, 4.597219e-10, 4.594176e-10, 4.599333e-10, 
    4.604262e-10, 4.612533e-10, 4.611173e-10, 4.614816e-10, 4.599198e-10, 
    4.609578e-10, 4.592441e-10, 4.597129e-10, 4.55983e-10, 4.545622e-10, 
    4.539575e-10, 4.534287e-10, 4.521414e-10, 4.530304e-10, 4.526799e-10, 
    4.535138e-10, 4.540434e-10, 4.537815e-10, 4.55398e-10, 4.547696e-10, 
    4.580789e-10, 4.566537e-10, 4.603687e-10, 4.5948e-10, 4.605817e-10, 
    4.600196e-10, 4.609826e-10, 4.601159e-10, 4.616172e-10, 4.61944e-10, 
    4.617207e-10, 4.625787e-10, 4.600679e-10, 4.610322e-10, 4.537741e-10, 
    4.538168e-10, 4.540159e-10, 4.531408e-10, 4.530872e-10, 4.522853e-10, 
    4.529989e-10, 4.533028e-10, 4.540741e-10, 4.545302e-10, 4.549638e-10, 
    4.559169e-10, 4.569811e-10, 4.584689e-10, 4.595377e-10, 4.602538e-10, 
    4.598147e-10, 4.602024e-10, 4.59769e-10, 4.595659e-10, 4.618215e-10, 
    4.605551e-10, 4.624553e-10, 4.623502e-10, 4.614903e-10, 4.62362e-10, 
    4.538468e-10, 4.53601e-10, 4.527472e-10, 4.534154e-10, 4.52198e-10, 
    4.528794e-10, 4.532711e-10, 4.547825e-10, 4.551147e-10, 4.554225e-10, 
    4.560305e-10, 4.568105e-10, 4.581786e-10, 4.593687e-10, 4.604549e-10, 
    4.603753e-10, 4.604033e-10, 4.606459e-10, 4.60045e-10, 4.607445e-10, 
    4.608619e-10, 4.60555e-10, 4.623361e-10, 4.618274e-10, 4.62348e-10, 
    4.620167e-10, 4.536809e-10, 4.540946e-10, 4.538711e-10, 4.542913e-10, 
    4.539952e-10, 4.553117e-10, 4.557063e-10, 4.575526e-10, 4.567952e-10, 
    4.580008e-10, 4.569177e-10, 4.571096e-10, 4.580399e-10, 4.569763e-10, 
    4.593029e-10, 4.577254e-10, 4.606553e-10, 4.590802e-10, 4.60754e-10, 
    4.604502e-10, 4.609532e-10, 4.614036e-10, 4.619703e-10, 4.630156e-10, 
    4.627736e-10, 4.636477e-10, 4.547112e-10, 4.552476e-10, 4.552005e-10, 
    4.557618e-10, 4.561768e-10, 4.570765e-10, 4.585188e-10, 4.579765e-10, 
    4.589722e-10, 4.59172e-10, 4.576594e-10, 4.585881e-10, 4.556066e-10, 
    4.560883e-10, 4.558016e-10, 4.547535e-10, 4.581013e-10, 4.563835e-10, 
    4.595553e-10, 4.586251e-10, 4.613394e-10, 4.599896e-10, 4.626403e-10, 
    4.637727e-10, 4.648388e-10, 4.660836e-10, 4.555404e-10, 4.55176e-10, 
    4.558286e-10, 4.567311e-10, 4.575687e-10, 4.586818e-10, 4.587957e-10, 
    4.590042e-10, 4.595442e-10, 4.599982e-10, 4.590699e-10, 4.60112e-10, 
    4.561998e-10, 4.582505e-10, 4.550381e-10, 4.560055e-10, 4.566779e-10, 
    4.563831e-10, 4.579146e-10, 4.582754e-10, 4.597414e-10, 4.589837e-10, 
    4.634931e-10, 4.614986e-10, 4.670316e-10, 4.65486e-10, 4.550486e-10, 
    4.555392e-10, 4.57246e-10, 4.56434e-10, 4.587561e-10, 4.593275e-10, 
    4.59792e-10, 4.603855e-10, 4.604497e-10, 4.608013e-10, 4.602251e-10, 
    4.607786e-10, 4.586841e-10, 4.596202e-10, 4.570511e-10, 4.576765e-10, 
    4.573888e-10, 4.570732e-10, 4.580473e-10, 4.590845e-10, 4.591069e-10, 
    4.594394e-10, 4.603759e-10, 4.587656e-10, 4.637501e-10, 4.606721e-10, 
    4.560741e-10, 4.570185e-10, 4.571536e-10, 4.567878e-10, 4.592702e-10, 
    4.583709e-10, 4.607928e-10, 4.601384e-10, 4.612106e-10, 4.606778e-10, 
    4.605994e-10, 4.599151e-10, 4.594889e-10, 4.584121e-10, 4.575358e-10, 
    4.568409e-10, 4.570025e-10, 4.577658e-10, 4.59148e-10, 4.604554e-10, 
    4.60169e-10, 4.611291e-10, 4.585878e-10, 4.596535e-10, 4.592416e-10, 
    4.603156e-10, 4.579621e-10, 4.599657e-10, 4.574497e-10, 4.576704e-10, 
    4.58353e-10, 4.597256e-10, 4.600295e-10, 4.603536e-10, 4.601537e-10, 
    4.591832e-10, 4.590242e-10, 4.583365e-10, 4.581465e-10, 4.576224e-10, 
    4.571884e-10, 4.575849e-10, 4.580012e-10, 4.591836e-10, 4.602489e-10, 
    4.6141e-10, 4.616942e-10, 4.630499e-10, 4.619461e-10, 4.637672e-10, 
    4.622186e-10, 4.648993e-10, 4.600821e-10, 4.621734e-10, 4.583841e-10, 
    4.587926e-10, 4.59531e-10, 4.612246e-10, 4.603106e-10, 4.613796e-10, 
    4.59018e-10, 4.57792e-10, 4.57475e-10, 4.568831e-10, 4.574885e-10, 
    4.574393e-10, 4.580186e-10, 4.578324e-10, 4.592229e-10, 4.584761e-10, 
    4.605974e-10, 4.613712e-10, 4.63556e-10, 4.648947e-10, 4.662574e-10, 
    4.668587e-10, 4.670417e-10, 4.671182e-10 ;

 SOIL1C_vr =
  19.98041, 19.98036, 19.98037, 19.98033, 19.98035, 19.98032, 19.9804, 
    19.98036, 19.98038, 19.98041, 19.98025, 19.98033, 19.98017, 19.98022, 
    19.9801, 19.98018, 19.98008, 19.9801, 19.98004, 19.98006, 19.97999, 
    19.98004, 19.97995, 19.98, 19.97999, 19.98004, 19.98031, 19.98026, 
    19.98031, 19.98031, 19.98031, 19.98035, 19.98037, 19.98041, 19.98041, 
    19.98038, 19.9803, 19.98033, 19.98027, 19.98027, 19.9802, 19.98023, 
    19.98012, 19.98015, 19.98006, 19.98008, 19.98006, 19.98007, 19.98006, 
    19.98009, 19.98008, 19.98011, 19.98023, 19.98019, 19.9803, 19.98036, 
    19.9804, 19.98043, 19.98042, 19.98042, 19.98037, 19.98034, 19.98031, 
    19.98029, 19.98027, 19.98021, 19.98018, 19.98011, 19.98013, 19.9801, 
    19.98008, 19.98005, 19.98005, 19.98004, 19.9801, 19.98006, 19.98013, 
    19.98011, 19.98026, 19.98032, 19.98035, 19.98037, 19.98042, 19.98038, 
    19.9804, 19.98036, 19.98034, 19.98035, 19.98029, 19.98031, 19.98018, 
    19.98024, 19.98009, 19.98012, 19.98008, 19.9801, 19.98006, 19.9801, 
    19.98004, 19.98002, 19.98003, 19.98, 19.9801, 19.98006, 19.98035, 
    19.98035, 19.98034, 19.98038, 19.98038, 19.98041, 19.98038, 19.98037, 
    19.98034, 19.98032, 19.9803, 19.98027, 19.98022, 19.98016, 19.98012, 
    19.98009, 19.98011, 19.98009, 19.98011, 19.98012, 19.98003, 19.98008, 
    19.98, 19.98001, 19.98004, 19.98001, 19.98035, 19.98036, 19.98039, 
    19.98037, 19.98042, 19.98039, 19.98037, 19.98031, 19.9803, 19.98029, 
    19.98026, 19.98023, 19.98018, 19.98013, 19.98008, 19.98009, 19.98009, 
    19.98007, 19.9801, 19.98007, 19.98007, 19.98008, 19.98001, 19.98003, 
    19.98001, 19.98002, 19.98036, 19.98034, 19.98035, 19.98033, 19.98034, 
    19.98029, 19.98027, 19.9802, 19.98023, 19.98018, 19.98023, 19.98022, 
    19.98018, 19.98022, 19.98013, 19.98019, 19.98007, 19.98014, 19.98007, 
    19.98008, 19.98006, 19.98004, 19.98002, 19.97998, 19.97999, 19.97995, 
    19.98031, 19.98029, 19.9803, 19.98027, 19.98026, 19.98022, 19.98016, 
    19.98018, 19.98014, 19.98013, 19.9802, 19.98016, 19.98028, 19.98026, 
    19.98027, 19.98031, 19.98018, 19.98025, 19.98012, 19.98016, 19.98005, 
    19.9801, 19.97999, 19.97995, 19.97991, 19.97986, 19.98028, 19.9803, 
    19.98027, 19.98023, 19.9802, 19.98015, 19.98015, 19.98014, 19.98012, 
    19.9801, 19.98014, 19.9801, 19.98026, 19.98017, 19.9803, 19.98026, 
    19.98024, 19.98025, 19.98018, 19.98017, 19.98011, 19.98014, 19.97996, 
    19.98004, 19.97982, 19.97988, 19.9803, 19.98028, 19.98021, 19.98025, 
    19.98015, 19.98013, 19.98011, 19.98009, 19.98008, 19.98007, 19.98009, 
    19.98007, 19.98015, 19.98012, 19.98022, 19.98019, 19.98021, 19.98022, 
    19.98018, 19.98014, 19.98014, 19.98012, 19.98009, 19.98015, 19.97995, 
    19.98007, 19.98026, 19.98022, 19.98022, 19.98023, 19.98013, 19.98017, 
    19.98007, 19.98009, 19.98005, 19.98007, 19.98008, 19.9801, 19.98012, 
    19.98017, 19.9802, 19.98023, 19.98022, 19.98019, 19.98013, 19.98008, 
    19.98009, 19.98005, 19.98016, 19.98012, 19.98013, 19.98009, 19.98018, 
    19.9801, 19.9802, 19.9802, 19.98017, 19.98011, 19.9801, 19.98009, 
    19.98009, 19.98013, 19.98014, 19.98017, 19.98018, 19.9802, 19.98022, 
    19.9802, 19.98018, 19.98013, 19.98009, 19.98004, 19.98003, 19.97998, 
    19.98002, 19.97995, 19.98001, 19.9799, 19.9801, 19.98001, 19.98017, 
    19.98015, 19.98012, 19.98005, 19.98009, 19.98005, 19.98014, 19.98019, 
    19.9802, 19.98023, 19.9802, 19.9802, 19.98018, 19.98019, 19.98013, 
    19.98016, 19.98008, 19.98005, 19.97996, 19.9799, 19.97985, 19.97982, 
    19.97982, 19.97981,
  19.98022, 19.98017, 19.98018, 19.98014, 19.98016, 19.98013, 19.98021, 
    19.98017, 19.9802, 19.98022, 19.98006, 19.98014, 19.97997, 19.98002, 
    19.9799, 19.97998, 19.97988, 19.9799, 19.97984, 19.97986, 19.97978, 
    19.97983, 19.97974, 19.9798, 19.97979, 19.97984, 19.98012, 19.98007, 
    19.98012, 19.98012, 19.98012, 19.98016, 19.98018, 19.98023, 19.98022, 
    19.98019, 19.98011, 19.98014, 19.98007, 19.98008, 19.98001, 19.98004, 
    19.97992, 19.97995, 19.97986, 19.97988, 19.97986, 19.97987, 19.97986, 
    19.97989, 19.97988, 19.97991, 19.98003, 19.98, 19.9801, 19.98017, 
    19.98021, 19.98024, 19.98024, 19.98023, 19.98019, 19.98015, 19.98012, 
    19.9801, 19.98008, 19.98002, 19.97998, 19.97991, 19.97993, 19.9799, 
    19.97988, 19.97985, 19.97985, 19.97984, 19.97991, 19.97986, 19.97993, 
    19.97991, 19.98007, 19.98013, 19.98016, 19.98018, 19.98023, 19.9802, 
    19.98021, 19.98018, 19.98015, 19.98016, 19.98009, 19.98012, 19.97998, 
    19.98004, 19.97989, 19.97992, 19.97988, 19.9799, 19.97986, 19.9799, 
    19.97983, 19.97982, 19.97983, 19.97979, 19.9799, 19.97986, 19.98016, 
    19.98016, 19.98015, 19.98019, 19.98019, 19.98023, 19.9802, 19.98018, 
    19.98015, 19.98013, 19.98011, 19.98007, 19.98003, 19.97997, 19.97992, 
    19.97989, 19.97991, 19.97989, 19.97991, 19.97992, 19.97983, 19.97988, 
    19.9798, 19.9798, 19.97984, 19.9798, 19.98016, 19.98017, 19.98021, 
    19.98018, 19.98023, 19.9802, 19.98018, 19.98012, 19.98011, 19.98009, 
    19.98007, 19.98004, 19.97998, 19.97993, 19.97988, 19.97989, 19.97989, 
    19.97988, 19.9799, 19.97987, 19.97987, 19.97988, 19.9798, 19.97983, 
    19.9798, 19.97982, 19.98017, 19.98015, 19.98016, 19.98014, 19.98015, 
    19.9801, 19.98008, 19.98001, 19.98004, 19.97999, 19.98003, 19.98002, 
    19.97998, 19.98003, 19.97993, 19.98, 19.97987, 19.97994, 19.97987, 
    19.97988, 19.97986, 19.97984, 19.97982, 19.97978, 19.97979, 19.97975, 
    19.98012, 19.9801, 19.9801, 19.98008, 19.98006, 19.98002, 19.97996, 
    19.97999, 19.97994, 19.97994, 19.98, 19.97996, 19.98009, 19.98007, 
    19.98008, 19.98012, 19.97998, 19.98005, 19.97992, 19.97996, 19.97985, 
    19.9799, 19.97979, 19.97974, 19.9797, 19.97965, 19.98009, 19.9801, 
    19.98008, 19.98004, 19.98, 19.97996, 19.97995, 19.97994, 19.97992, 
    19.9799, 19.97994, 19.9799, 19.98006, 19.97997, 19.98011, 19.98007, 
    19.98004, 19.98005, 19.97999, 19.97997, 19.97991, 19.97994, 19.97976, 
    19.97984, 19.97961, 19.97967, 19.98011, 19.98009, 19.98002, 19.98005, 
    19.97995, 19.97993, 19.97991, 19.97989, 19.97988, 19.97987, 19.97989, 
    19.97987, 19.97996, 19.97992, 19.98003, 19.98, 19.98001, 19.98002, 
    19.97998, 19.97994, 19.97994, 19.97993, 19.97989, 19.97995, 19.97974, 
    19.97987, 19.98007, 19.98003, 19.98002, 19.98004, 19.97993, 19.97997, 
    19.97987, 19.9799, 19.97985, 19.97987, 19.97988, 19.97991, 19.97992, 
    19.97997, 19.98001, 19.98003, 19.98003, 19.98, 19.97994, 19.97988, 
    19.97989, 19.97985, 19.97996, 19.97992, 19.97993, 19.97989, 19.97999, 
    19.9799, 19.98001, 19.98, 19.97997, 19.97991, 19.9799, 19.97989, 
    19.97989, 19.97994, 19.97994, 19.97997, 19.97998, 19.98, 19.98002, 19.98, 
    19.97999, 19.97994, 19.97989, 19.97984, 19.97983, 19.97977, 19.97982, 
    19.97974, 19.97981, 19.9797, 19.9799, 19.97981, 19.97997, 19.97995, 
    19.97992, 19.97985, 19.97989, 19.97985, 19.97994, 19.97999, 19.98001, 
    19.98003, 19.98001, 19.98001, 19.97998, 19.97999, 19.97993, 19.97997, 
    19.97988, 19.97985, 19.97975, 19.9797, 19.97964, 19.97961, 19.97961, 
    19.9796,
  19.98016, 19.9801, 19.98011, 19.98007, 19.98009, 19.98007, 19.98015, 
    19.9801, 19.98013, 19.98015, 19.97999, 19.98007, 19.97991, 19.97996, 
    19.97983, 19.97991, 19.97981, 19.97983, 19.97977, 19.97979, 19.97971, 
    19.97976, 19.97967, 19.97972, 19.97972, 19.97976, 19.98005, 19.98, 
    19.98006, 19.98005, 19.98005, 19.98009, 19.98012, 19.98016, 19.98015, 
    19.98012, 19.98005, 19.98007, 19.98001, 19.98001, 19.97994, 19.97997, 
    19.97985, 19.97989, 19.97979, 19.97981, 19.97979, 19.9798, 19.97979, 
    19.97982, 19.97981, 19.97984, 19.97996, 19.97993, 19.98004, 19.9801, 
    19.98014, 19.98018, 19.98017, 19.98016, 19.98012, 19.98008, 19.98005, 
    19.98003, 19.98001, 19.97995, 19.97992, 19.97984, 19.97986, 19.97984, 
    19.97981, 19.97978, 19.97978, 19.97977, 19.97984, 19.97979, 19.97986, 
    19.97985, 19.98, 19.98006, 19.98009, 19.98011, 19.98017, 19.98013, 
    19.98014, 19.98011, 19.98009, 19.9801, 19.98003, 19.98005, 19.97991, 
    19.97997, 19.97982, 19.97985, 19.97981, 19.97983, 19.97979, 19.97983, 
    19.97976, 19.97975, 19.97976, 19.97972, 19.97983, 19.97979, 19.9801, 
    19.9801, 19.98009, 19.98013, 19.98013, 19.98016, 19.98013, 19.98012, 
    19.98009, 19.98007, 19.98005, 19.98001, 19.97996, 19.9799, 19.97985, 
    19.97982, 19.97984, 19.97982, 19.97984, 19.97985, 19.97976, 19.97981, 
    19.97973, 19.97973, 19.97977, 19.97973, 19.98009, 19.9801, 19.98014, 
    19.98011, 19.98017, 19.98014, 19.98012, 19.98005, 19.98004, 19.98003, 
    19.98, 19.97997, 19.97991, 19.97986, 19.97981, 19.97982, 19.97981, 
    19.9798, 19.97983, 19.9798, 19.9798, 19.97981, 19.97973, 19.97975, 
    19.97973, 19.97975, 19.9801, 19.98008, 19.98009, 19.98008, 19.98009, 
    19.98003, 19.98001, 19.97994, 19.97997, 19.97992, 19.97996, 19.97996, 
    19.97992, 19.97996, 19.97986, 19.97993, 19.9798, 19.97987, 19.9798, 
    19.97981, 19.97979, 19.97977, 19.97975, 19.9797, 19.97971, 19.97968, 
    19.98006, 19.98004, 19.98004, 19.98001, 19.98, 19.97996, 19.97989, 
    19.97992, 19.97988, 19.97987, 19.97993, 19.97989, 19.98002, 19.98, 
    19.98001, 19.98006, 19.97991, 19.97999, 19.97985, 19.97989, 19.97977, 
    19.97983, 19.97972, 19.97967, 19.97963, 19.97957, 19.98002, 19.98004, 
    19.98001, 19.97997, 19.97994, 19.97989, 19.97988, 19.97988, 19.97985, 
    19.97983, 19.97987, 19.97983, 19.97999, 19.97991, 19.98004, 19.98, 
    19.97997, 19.97999, 19.97992, 19.97991, 19.97984, 19.97988, 19.97968, 
    19.97977, 19.97953, 19.9796, 19.98004, 19.98002, 19.97995, 19.97998, 
    19.97989, 19.97986, 19.97984, 19.97982, 19.97981, 19.9798, 19.97982, 
    19.9798, 19.97989, 19.97985, 19.97996, 19.97993, 19.97994, 19.97996, 
    19.97992, 19.97987, 19.97987, 19.97986, 19.97982, 19.97989, 19.97967, 
    19.9798, 19.98, 19.97996, 19.97995, 19.97997, 19.97986, 19.9799, 19.9798, 
    19.97983, 19.97978, 19.9798, 19.97981, 19.97984, 19.97985, 19.9799, 
    19.97994, 19.97997, 19.97996, 19.97993, 19.97987, 19.97981, 19.97982, 
    19.97978, 19.97989, 19.97985, 19.97986, 19.97982, 19.97992, 19.97983, 
    19.97994, 19.97993, 19.9799, 19.97984, 19.97983, 19.97982, 19.97983, 
    19.97987, 19.97987, 19.9799, 19.97991, 19.97993, 19.97995, 19.97993, 
    19.97992, 19.97987, 19.97982, 19.97977, 19.97976, 19.9797, 19.97975, 
    19.97967, 19.97974, 19.97962, 19.97983, 19.97974, 19.9799, 19.97988, 
    19.97985, 19.97978, 19.97982, 19.97977, 19.97987, 19.97993, 19.97994, 
    19.97997, 19.97994, 19.97994, 19.97992, 19.97993, 19.97987, 19.9799, 
    19.97981, 19.97977, 19.97968, 19.97962, 19.97957, 19.97954, 19.97953, 
    19.97953,
  19.98076, 19.98071, 19.98072, 19.98068, 19.9807, 19.98067, 19.98075, 
    19.98071, 19.98074, 19.98076, 19.9806, 19.98068, 19.98051, 19.98057, 
    19.98044, 19.98052, 19.98042, 19.98044, 19.98038, 19.9804, 19.98032, 
    19.98037, 19.98028, 19.98034, 19.98033, 19.98038, 19.98066, 19.98061, 
    19.98067, 19.98066, 19.98066, 19.9807, 19.98072, 19.98077, 19.98076, 
    19.98073, 19.98065, 19.98068, 19.98062, 19.98062, 19.98055, 19.98058, 
    19.98046, 19.98049, 19.9804, 19.98042, 19.9804, 19.98041, 19.9804, 
    19.98043, 19.98042, 19.98045, 19.98057, 19.98054, 19.98064, 19.98071, 
    19.98075, 19.98078, 19.98078, 19.98077, 19.98073, 19.98069, 19.98066, 
    19.98064, 19.98062, 19.98056, 19.98053, 19.98045, 19.98047, 19.98045, 
    19.98042, 19.98039, 19.98039, 19.98038, 19.98045, 19.9804, 19.98047, 
    19.98045, 19.98061, 19.98067, 19.9807, 19.98072, 19.98077, 19.98074, 
    19.98075, 19.98071, 19.98069, 19.98071, 19.98064, 19.98066, 19.98052, 
    19.98058, 19.98043, 19.98046, 19.98042, 19.98044, 19.9804, 19.98044, 
    19.98037, 19.98036, 19.98037, 19.98033, 19.98044, 19.9804, 19.98071, 
    19.9807, 19.98069, 19.98073, 19.98073, 19.98077, 19.98074, 19.98072, 
    19.98069, 19.98067, 19.98065, 19.98061, 19.98057, 19.98051, 19.98046, 
    19.98043, 19.98045, 19.98043, 19.98045, 19.98046, 19.98037, 19.98042, 
    19.98034, 19.98034, 19.98038, 19.98034, 19.9807, 19.98071, 19.98075, 
    19.98072, 19.98077, 19.98074, 19.98073, 19.98066, 19.98065, 19.98063, 
    19.98061, 19.98058, 19.98052, 19.98047, 19.98042, 19.98043, 19.98042, 
    19.98042, 19.98044, 19.98041, 19.98041, 19.98042, 19.98034, 19.98037, 
    19.98034, 19.98036, 19.98071, 19.98069, 19.9807, 19.98068, 19.9807, 
    19.98064, 19.98062, 19.98055, 19.98058, 19.98053, 19.98057, 19.98056, 
    19.98052, 19.98057, 19.98047, 19.98054, 19.98042, 19.98048, 19.98041, 
    19.98042, 19.9804, 19.98038, 19.98036, 19.98032, 19.98033, 19.98029, 
    19.98067, 19.98064, 19.98064, 19.98062, 19.9806, 19.98057, 19.9805, 
    19.98053, 19.98049, 19.98048, 19.98054, 19.9805, 19.98063, 19.98061, 
    19.98062, 19.98066, 19.98052, 19.98059, 19.98046, 19.9805, 19.98039, 
    19.98044, 19.98033, 19.98028, 19.98024, 19.98019, 19.98063, 19.98065, 
    19.98062, 19.98058, 19.98055, 19.9805, 19.98049, 19.98048, 19.98046, 
    19.98044, 19.98048, 19.98044, 19.9806, 19.98052, 19.98065, 19.98061, 
    19.98058, 19.98059, 19.98053, 19.98051, 19.98045, 19.98049, 19.9803, 
    19.98038, 19.98015, 19.98021, 19.98065, 19.98063, 19.98056, 19.98059, 
    19.9805, 19.98047, 19.98045, 19.98043, 19.98042, 19.98041, 19.98043, 
    19.98041, 19.9805, 19.98046, 19.98057, 19.98054, 19.98055, 19.98057, 
    19.98052, 19.98048, 19.98048, 19.98046, 19.98043, 19.98049, 19.98028, 
    19.98041, 19.98061, 19.98057, 19.98056, 19.98058, 19.98047, 19.98051, 
    19.98041, 19.98044, 19.98039, 19.98041, 19.98042, 19.98045, 19.98046, 
    19.98051, 19.98055, 19.98058, 19.98057, 19.98054, 19.98048, 19.98042, 
    19.98043, 19.98039, 19.9805, 19.98046, 19.98047, 19.98043, 19.98053, 
    19.98044, 19.98055, 19.98054, 19.98051, 19.98045, 19.98044, 19.98043, 
    19.98044, 19.98048, 19.98048, 19.98051, 19.98052, 19.98054, 19.98056, 
    19.98054, 19.98053, 19.98048, 19.98043, 19.98038, 19.98037, 19.98031, 
    19.98036, 19.98028, 19.98035, 19.98024, 19.98044, 19.98035, 19.98051, 
    19.98049, 19.98046, 19.98039, 19.98043, 19.98038, 19.98048, 19.98054, 
    19.98055, 19.98057, 19.98055, 19.98055, 19.98053, 19.98053, 19.98047, 
    19.98051, 19.98042, 19.98038, 19.98029, 19.98024, 19.98018, 19.98015, 
    19.98015, 19.98014,
  19.98279, 19.98274, 19.98275, 19.98272, 19.98274, 19.98271, 19.98278, 
    19.98274, 19.98277, 19.98279, 19.98264, 19.98271, 19.98256, 19.98261, 
    19.98249, 19.98257, 19.98248, 19.98249, 19.98244, 19.98245, 19.98238, 
    19.98243, 19.98235, 19.9824, 19.98239, 19.98243, 19.9827, 19.98265, 
    19.9827, 19.98269, 19.9827, 19.98274, 19.98276, 19.9828, 19.98279, 
    19.98276, 19.98269, 19.98271, 19.98266, 19.98266, 19.98259, 19.98262, 
    19.98251, 19.98254, 19.98245, 19.98248, 19.98245, 19.98246, 19.98245, 
    19.98249, 19.98247, 19.9825, 19.98262, 19.98258, 19.98268, 19.98274, 
    19.98278, 19.98281, 19.98281, 19.9828, 19.98276, 19.98272, 19.98269, 
    19.98268, 19.98266, 19.9826, 19.98257, 19.98251, 19.98252, 19.9825, 
    19.98248, 19.98244, 19.98245, 19.98244, 19.9825, 19.98246, 19.98252, 
    19.98251, 19.98265, 19.98271, 19.98273, 19.98275, 19.9828, 19.98277, 
    19.98278, 19.98275, 19.98273, 19.98274, 19.98268, 19.9827, 19.98257, 
    19.98263, 19.98248, 19.98252, 19.98247, 19.98249, 19.98246, 19.98249, 
    19.98243, 19.98242, 19.98243, 19.98239, 19.98249, 19.98245, 19.98274, 
    19.98274, 19.98273, 19.98276, 19.98277, 19.9828, 19.98277, 19.98276, 
    19.98273, 19.98271, 19.98269, 19.98265, 19.98261, 19.98256, 19.98251, 
    19.98248, 19.9825, 19.98249, 19.9825, 19.98251, 19.98242, 19.98247, 
    19.9824, 19.9824, 19.98244, 19.9824, 19.98274, 19.98275, 19.98278, 
    19.98275, 19.9828, 19.98277, 19.98276, 19.9827, 19.98269, 19.98267, 
    19.98265, 19.98262, 19.98257, 19.98252, 19.98248, 19.98248, 19.98248, 
    19.98247, 19.98249, 19.98247, 19.98246, 19.98247, 19.9824, 19.98242, 
    19.9824, 19.98242, 19.98274, 19.98273, 19.98273, 19.98272, 19.98273, 
    19.98268, 19.98266, 19.98259, 19.98262, 19.98257, 19.98262, 19.98261, 
    19.98257, 19.98261, 19.98252, 19.98258, 19.98247, 19.98253, 19.98247, 
    19.98248, 19.98246, 19.98244, 19.98242, 19.98238, 19.98239, 19.98235, 
    19.9827, 19.98268, 19.98268, 19.98266, 19.98265, 19.98261, 19.98255, 
    19.98257, 19.98253, 19.98253, 19.98259, 19.98255, 19.98267, 19.98265, 
    19.98266, 19.9827, 19.98257, 19.98264, 19.98251, 19.98255, 19.98244, 
    19.98249, 19.98239, 19.98235, 19.9823, 19.98226, 19.98267, 19.98268, 
    19.98266, 19.98262, 19.98259, 19.98255, 19.98254, 19.98253, 19.98251, 
    19.98249, 19.98253, 19.98249, 19.98264, 19.98256, 19.98269, 19.98265, 
    19.98262, 19.98264, 19.98258, 19.98256, 19.9825, 19.98253, 19.98236, 
    19.98244, 19.98222, 19.98228, 19.98269, 19.98267, 19.9826, 19.98263, 
    19.98254, 19.98252, 19.9825, 19.98248, 19.98248, 19.98246, 19.98249, 
    19.98246, 19.98255, 19.98251, 19.98261, 19.98259, 19.9826, 19.98261, 
    19.98257, 19.98253, 19.98253, 19.98252, 19.98248, 19.98254, 19.98235, 
    19.98247, 19.98265, 19.98261, 19.98261, 19.98262, 19.98252, 19.98256, 
    19.98246, 19.98249, 19.98245, 19.98247, 19.98247, 19.9825, 19.98252, 
    19.98256, 19.98259, 19.98262, 19.98261, 19.98258, 19.98253, 19.98248, 
    19.98249, 19.98245, 19.98255, 19.98251, 19.98252, 19.98248, 19.98257, 
    19.9825, 19.9826, 19.98259, 19.98256, 19.98251, 19.98249, 19.98248, 
    19.98249, 19.98253, 19.98253, 19.98256, 19.98257, 19.98259, 19.9826, 
    19.98259, 19.98257, 19.98253, 19.98248, 19.98244, 19.98243, 19.98237, 
    19.98242, 19.98235, 19.98241, 19.9823, 19.98249, 19.98241, 19.98256, 
    19.98254, 19.98251, 19.98245, 19.98248, 19.98244, 19.98253, 19.98258, 
    19.98259, 19.98262, 19.98259, 19.9826, 19.98257, 19.98258, 19.98252, 
    19.98255, 19.98247, 19.98244, 19.98236, 19.9823, 19.98225, 19.98223, 
    19.98222, 19.98221,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N =
  0.722154, 0.7221522, 0.7221525, 0.7221511, 0.7221519, 0.7221509, 0.7221537, 
    0.7221521, 0.7221531, 0.7221538, 0.7221482, 0.722151, 0.7221453, 
    0.7221471, 0.7221426, 0.7221456, 0.722142, 0.7221427, 0.7221407, 
    0.7221413, 0.7221386, 0.7221404, 0.7221373, 0.7221391, 0.7221388, 
    0.7221404, 0.7221504, 0.7221486, 0.7221506, 0.7221503, 0.7221504, 
    0.7221519, 0.7221526, 0.7221541, 0.7221539, 0.7221528, 0.7221501, 
    0.722151, 0.7221488, 0.7221489, 0.7221465, 0.7221475, 0.7221434, 
    0.7221446, 0.7221412, 0.722142, 0.7221413, 0.7221415, 0.7221413, 
    0.7221425, 0.722142, 0.7221431, 0.7221473, 0.7221461, 0.7221498, 
    0.7221521, 0.7221536, 0.7221547, 0.7221545, 0.7221542, 0.7221528, 
    0.7221513, 0.7221503, 0.7221496, 0.7221489, 0.7221468, 0.7221457, 
    0.7221432, 0.7221437, 0.7221429, 0.7221422, 0.7221409, 0.7221411, 
    0.7221406, 0.7221429, 0.7221414, 0.7221439, 0.7221432, 0.7221487, 
    0.7221508, 0.7221517, 0.7221525, 0.7221544, 0.7221531, 0.7221536, 
    0.7221524, 0.7221516, 0.7221519, 0.7221496, 0.7221505, 0.7221456, 
    0.7221477, 0.7221422, 0.7221435, 0.7221419, 0.7221428, 0.7221413, 
    0.7221426, 0.7221404, 0.7221399, 0.7221403, 0.722139, 0.7221427, 
    0.7221413, 0.722152, 0.7221519, 0.7221516, 0.7221529, 0.722153, 
    0.7221542, 0.7221531, 0.7221527, 0.7221515, 0.7221509, 0.7221502, 
    0.7221488, 0.7221472, 0.722145, 0.7221435, 0.7221424, 0.7221431, 
    0.7221425, 0.7221431, 0.7221434, 0.7221401, 0.722142, 0.7221392, 
    0.7221393, 0.7221406, 0.7221393, 0.7221519, 0.7221522, 0.7221535, 
    0.7221525, 0.7221543, 0.7221533, 0.7221527, 0.7221505, 0.72215, 
    0.7221496, 0.7221487, 0.7221475, 0.7221455, 0.7221437, 0.7221421, 
    0.7221422, 0.7221422, 0.7221418, 0.7221427, 0.7221417, 0.7221415, 
    0.722142, 0.7221394, 0.7221401, 0.7221393, 0.7221398, 0.7221521, 
    0.7221515, 0.7221518, 0.7221512, 0.7221516, 0.7221497, 0.7221491, 
    0.7221464, 0.7221475, 0.7221457, 0.7221473, 0.722147, 0.7221457, 
    0.7221472, 0.7221438, 0.7221462, 0.7221418, 0.7221441, 0.7221417, 
    0.7221421, 0.7221414, 0.7221407, 0.7221399, 0.7221383, 0.7221387, 
    0.7221374, 0.7221506, 0.7221498, 0.7221498, 0.722149, 0.7221484, 
    0.7221471, 0.722145, 0.7221458, 0.7221443, 0.722144, 0.7221462, 
    0.7221448, 0.7221493, 0.7221485, 0.722149, 0.7221505, 0.7221456, 
    0.7221481, 0.7221434, 0.7221448, 0.7221408, 0.7221428, 0.7221389, 
    0.7221372, 0.7221357, 0.7221338, 0.7221494, 0.7221499, 0.722149, 
    0.7221476, 0.7221464, 0.7221447, 0.7221445, 0.7221442, 0.7221435, 
    0.7221428, 0.7221441, 0.7221426, 0.7221484, 0.7221454, 0.7221501, 
    0.7221487, 0.7221477, 0.7221481, 0.7221459, 0.7221453, 0.7221432, 
    0.7221443, 0.7221376, 0.7221406, 0.7221324, 0.7221347, 0.7221501, 
    0.7221494, 0.7221469, 0.7221481, 0.7221446, 0.7221438, 0.7221431, 
    0.7221422, 0.7221421, 0.7221416, 0.7221425, 0.7221416, 0.7221447, 
    0.7221434, 0.7221471, 0.7221462, 0.7221466, 0.7221471, 0.7221457, 
    0.7221441, 0.7221441, 0.7221436, 0.7221422, 0.7221446, 0.7221373, 
    0.7221418, 0.7221486, 0.7221472, 0.722147, 0.7221475, 0.7221439, 
    0.7221452, 0.7221416, 0.7221426, 0.722141, 0.7221418, 0.7221419, 
    0.7221429, 0.7221435, 0.7221451, 0.7221464, 0.7221475, 0.7221472, 
    0.7221461, 0.7221441, 0.7221421, 0.7221425, 0.7221411, 0.7221448, 
    0.7221433, 0.7221439, 0.7221423, 0.7221458, 0.7221428, 0.7221466, 
    0.7221462, 0.7221452, 0.7221432, 0.7221428, 0.7221423, 0.7221426, 
    0.722144, 0.7221442, 0.7221453, 0.7221455, 0.7221463, 0.7221469, 
    0.7221463, 0.7221457, 0.722144, 0.7221424, 0.7221407, 0.7221403, 
    0.7221383, 0.7221399, 0.7221372, 0.7221395, 0.7221355, 0.7221426, 
    0.7221396, 0.7221451, 0.7221445, 0.7221435, 0.722141, 0.7221423, 
    0.7221407, 0.7221442, 0.722146, 0.7221465, 0.7221474, 0.7221465, 
    0.7221466, 0.7221457, 0.722146, 0.7221439, 0.722145, 0.7221419, 
    0.7221408, 0.7221375, 0.7221355, 0.7221336, 0.7221327, 0.7221324, 
    0.7221323 ;

 SOIL1N_TNDNCY_VERT_TRANS =
  0, -5.139921e-21, 3.083953e-20, 1.541976e-20, -5.139921e-21, 1.027984e-20, 
    2.569961e-20, 1.027984e-20, 5.139921e-21, 0, -2.055969e-20, 
    -3.083953e-20, 2.006177e-36, 5.139921e-21, -5.139921e-21, 0, 
    -1.027984e-20, 5.139921e-21, -1.541976e-20, 3.083953e-20, 1.541976e-20, 
    -3.083953e-20, 1.541976e-20, 5.139921e-21, 2.006177e-36, -1.027984e-20, 
    0, -3.597945e-20, 5.139921e-21, 0, -3.083953e-20, 2.055969e-20, 
    5.139921e-21, -2.569961e-20, -5.139921e-21, 5.139921e-21, -2.055969e-20, 
    -3.083953e-20, 5.139921e-21, -1.027984e-20, 1.027984e-20, 3.083953e-20, 
    1.541976e-20, 4.111937e-20, -3.083953e-20, -1.027984e-20, 3.083953e-20, 
    -5.139921e-21, 1.027984e-20, -1.027984e-20, -5.139921e-21, -1.027984e-20, 
    -2.569961e-20, 5.139921e-21, 5.139921e-21, 2.055969e-20, -3.083953e-20, 
    1.541976e-20, 2.569961e-20, 2.055969e-20, -4.111937e-20, 3.083953e-20, 
    1.027984e-20, 0, -5.139921e-21, 1.027984e-20, 5.139921e-21, 1.541976e-20, 
    1.541976e-20, -5.139921e-21, 1.541976e-20, -4.625929e-20, 0, 
    -1.027984e-20, -1.541976e-20, -2.055969e-20, -2.569961e-20, 5.139921e-21, 
    -1.027984e-20, 5.139921e-21, 2.055969e-20, 2.006177e-36, -5.139921e-21, 
    -1.541976e-20, -3.597945e-20, -1.027984e-20, 5.139921e-21, 3.083953e-20, 
    -5.139921e-21, -1.027984e-20, -2.569961e-20, 1.027984e-20, 0, 
    -2.055969e-20, 2.055969e-20, -5.139921e-21, 4.111937e-20, 1.541976e-20, 
    0, -5.139921e-21, -5.139921e-21, 3.083953e-20, 1.541976e-20, 
    -2.569961e-20, 3.083953e-20, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    -3.083953e-20, -5.139921e-21, 5.139921e-21, -1.027984e-20, 5.139921e-21, 
    1.541976e-20, 5.139921e-21, 1.541976e-20, 5.139921e-21, -5.139921e-21, 
    2.055969e-20, -1.541976e-20, -5.139921e-21, 3.083953e-20, 0, 
    1.027984e-20, -2.055969e-20, 2.569961e-20, -3.083953e-20, 1.541976e-20, 
    -2.055969e-20, -5.139921e-21, 2.569961e-20, 1.541976e-20, 2.569961e-20, 
    1.027984e-20, 2.569961e-20, 1.027984e-20, 2.006177e-36, 1.027984e-20, 
    5.139921e-21, 1.541976e-20, 5.139921e-21, 5.139921e-21, -1.027984e-20, 
    -2.006177e-36, 2.055969e-20, 2.569961e-20, 1.541976e-20, 1.027984e-20, 
    1.027984e-20, -1.541976e-20, 1.541976e-20, 5.139921e-21, -5.139921e-21, 
    -1.541976e-20, 2.569961e-20, 1.027984e-20, -2.569961e-20, -2.569961e-20, 
    -3.083953e-20, -1.027984e-20, -1.541976e-20, 3.597945e-20, 0, 
    2.006177e-36, 2.055969e-20, -5.139921e-21, 4.111937e-20, -5.139921e-21, 
    1.027984e-20, -2.006177e-36, 5.139921e-21, -2.055969e-20, 0, 
    -3.597945e-20, 5.139921e-21, -2.055969e-20, -1.027984e-20, -2.006177e-36, 
    -5.139921e-21, -5.139921e-21, 2.569961e-20, -1.027984e-20, 0, 
    5.139921e-21, -2.569961e-20, -1.027984e-20, 5.139921e-21, -1.027984e-20, 
    0, -2.006177e-36, -2.055969e-20, 5.139921e-21, -5.139921e-21, 
    -1.027984e-20, -2.055969e-20, 1.027984e-20, -5.139921e-21, 2.569961e-20, 
    -2.055969e-20, 2.055969e-20, 2.055969e-20, -2.055969e-20, -1.541976e-20, 
    5.139921e-21, -1.027984e-20, 0, 5.139921e-21, 2.569961e-20, 4.111937e-20, 
    0, 1.027984e-20, 1.541976e-20, -3.083953e-20, 0, -1.027984e-20, 
    2.006177e-36, -1.027984e-20, -2.569961e-20, -1.541976e-20, -5.139921e-21, 
    -2.055969e-20, -1.541976e-20, 2.055969e-20, 2.006177e-36, 0, 
    5.139921e-21, -2.006177e-36, -2.569961e-20, 1.541976e-20, -5.139921e-21, 
    -2.055969e-20, 1.027984e-20, -3.597945e-20, 5.139921e-21, -5.139921e-21, 
    -2.006177e-36, 0, -5.139921e-21, 3.083953e-20, 3.597945e-20, 
    1.027984e-20, -1.027984e-20, -1.027984e-20, -5.139921e-21, 5.139921e-21, 
    -3.597945e-20, -5.139921e-21, -2.569961e-20, -1.541976e-20, 
    -5.139921e-21, -5.139921e-21, -3.083953e-20, 5.139921e-21, 2.055969e-20, 
    5.139921e-21, 1.027984e-20, 1.027984e-20, -1.541976e-20, -2.569961e-20, 
    2.006177e-36, 2.055969e-20, 1.027984e-20, 3.597945e-20, -1.541976e-20, 
    3.597945e-20, -1.541976e-20, -1.027984e-20, -1.027984e-20, 4.111937e-20, 
    -3.083953e-20, -1.027984e-20, -2.569961e-20, -2.569961e-20, 
    -1.541976e-20, -3.597945e-20, 1.027984e-20, 2.569961e-20, 2.569961e-20, 
    -5.139921e-21, -1.541976e-20, -1.027984e-20, 5.139921e-21, -1.027984e-20, 
    -2.055969e-20, 1.541976e-20, 5.139921e-21, -3.083953e-20, -2.569961e-20, 
    -1.541976e-20, 2.055969e-20, 5.139921e-21, -5.139921e-21, 1.541976e-20, 
    5.139921e-21, -5.139921e-21, 0, 2.569961e-20, 2.055969e-20, 
    -2.055969e-20, -5.139921e-21, 1.541976e-20, -3.597945e-20, 3.597945e-20, 
    -3.597945e-20, 4.111937e-20, -2.006177e-36, 4.625929e-20, -2.569961e-20, 
    2.055969e-20, 3.597945e-20, 2.006177e-36, 2.006177e-36, 0, 0, 0, 
    2.055969e-20, -1.027984e-20, 0, -3.083953e-20, -1.541976e-20, 
    -1.027984e-20, -1.027984e-20, -5.139921e-21, 2.055969e-20, -4.111937e-20, 
    -1.541976e-20, -5.139921e-21, -2.055969e-20, 2.569961e-20, 5.139921e-21, 
    -1.027984e-20, -3.083953e-20, -4.625929e-20, 2.006177e-36, 1.027984e-20, 
    -1.541976e-20, -1.541976e-20, 1.027984e-20,
  1.027984e-20, -2.006177e-36, -5.139921e-21, -2.569961e-20, 1.027984e-20, 
    -1.541976e-20, 2.569961e-20, -5.139921e-21, 0, -1.541976e-20, 
    -1.027984e-20, -5.139921e-21, 1.541976e-20, 1.541976e-20, -1.027984e-20, 
    0, 5.139921e-21, 1.027984e-20, -5.139921e-21, -1.541976e-20, 
    -1.027984e-20, -2.569961e-20, 5.139921e-21, -2.006177e-36, 0, 
    2.055969e-20, -1.027984e-20, -5.139921e-21, 5.139921e-21, 1.541976e-20, 
    -2.055969e-20, -1.027984e-20, 1.541976e-20, 1.027984e-20, -1.027984e-20, 
    5.139921e-21, -5.139921e-21, -1.027984e-20, -5.139921e-21, -1.541976e-20, 
    1.027984e-20, 1.027984e-20, 2.055969e-20, -5.139921e-21, 5.139921e-21, 
    -3.083953e-20, 0, 5.139921e-21, 1.027984e-20, -5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, 1.541976e-20, -1.027984e-20, 
    0, 0, 0, -5.139921e-21, 5.139921e-21, 5.139921e-21, 3.597945e-20, 
    2.569961e-20, 2.569961e-20, 0, 2.569961e-20, 1.541976e-20, -3.083953e-20, 
    -1.541976e-20, -3.597945e-20, -1.541976e-20, 1.027984e-20, 1.541976e-20, 
    0, 1.027984e-20, -1.027984e-20, 1.541976e-20, -1.027984e-20, 
    3.083953e-20, -3.083953e-20, -2.569961e-20, -5.139921e-21, -5.139921e-21, 
    1.027984e-20, 3.083953e-20, -5.139921e-21, -2.055969e-20, -5.139921e-21, 
    2.055969e-20, 4.111937e-20, -1.027984e-20, 1.541976e-20, -5.139921e-21, 
    -1.027984e-20, 1.541976e-20, 2.569961e-20, 2.055969e-20, 2.569961e-20, 
    -5.139921e-21, 0, 3.083953e-20, -2.006177e-36, -1.541976e-20, 
    1.027984e-20, -2.055969e-20, 3.083953e-20, -1.027984e-20, 5.139921e-21, 
    -2.569961e-20, -5.139921e-21, 1.027984e-20, -5.139921e-21, -5.139921e-21, 
    5.139921e-21, 5.139921e-21, 2.569961e-20, -1.541976e-20, 2.006177e-36, 
    5.139921e-21, 5.139921e-21, -1.027984e-20, 5.139921e-21, 1.027984e-20, 
    2.055969e-20, 5.139921e-21, -2.569961e-20, 1.541976e-20, 5.139921e-21, 0, 
    5.139921e-21, -1.541976e-20, 5.139921e-21, 0, -5.139921e-21, 
    1.541976e-20, 2.006177e-36, -5.139921e-21, -5.139921e-21, -1.541976e-20, 
    -1.027984e-20, -1.541976e-20, -3.083953e-20, 1.027984e-20, -5.139921e-21, 
    2.006177e-36, -1.027984e-20, -5.139921e-21, 2.055969e-20, -2.569961e-20, 
    1.027984e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, -1.027984e-20, 
    -1.027984e-20, -5.139921e-20, 0, -5.139921e-21, 5.139921e-21, 0, 
    -5.139921e-21, 1.027984e-20, 1.541976e-20, -1.541976e-20, -2.055969e-20, 
    -1.027984e-20, -2.006177e-36, -2.055969e-20, 0, -1.027984e-20, 
    -5.139921e-21, 5.139921e-21, -1.027984e-20, 3.083953e-20, 1.027984e-20, 
    -1.027984e-20, -1.541976e-20, 1.027984e-20, -1.541976e-20, 1.027984e-20, 
    1.541976e-20, 3.083953e-20, -1.027984e-20, 5.139921e-21, -3.083953e-20, 
    -5.139921e-21, -5.139921e-21, -3.083953e-20, 5.139921e-21, 3.083953e-20, 
    -1.027984e-20, 3.083953e-20, 0, 2.569961e-20, 1.541976e-20, 
    -5.139921e-21, 5.139921e-21, 1.541976e-20, 5.139921e-20, 5.139921e-21, 
    1.027984e-20, -5.139921e-21, -3.083953e-20, -2.569961e-20, 3.597945e-20, 
    1.027984e-20, 0, 0, -2.006177e-36, -1.541976e-20, 1.541976e-20, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, 5.139921e-21, -2.055969e-20, 
    5.139921e-21, 2.569961e-20, -1.027984e-20, 1.541976e-20, -5.139921e-21, 
    5.139921e-21, 1.027984e-20, 5.139921e-21, 2.006177e-36, 1.027984e-20, 
    -1.027984e-20, 5.139921e-21, 1.541976e-20, 1.541976e-20, 2.055969e-20, 
    5.139921e-21, -1.027984e-20, -5.139921e-21, -5.139921e-21, 0, 
    -5.139921e-21, 1.541976e-20, -1.541976e-20, 2.055969e-20, -2.006177e-36, 
    -4.111937e-20, -5.139921e-21, -5.139921e-21, -3.083953e-20, 3.083953e-20, 
    5.139921e-21, 0, -5.139921e-21, -2.569961e-20, 1.027984e-20, 
    3.083953e-20, -1.027984e-20, -1.027984e-20, 1.541976e-20, -3.083953e-20, 
    3.083953e-20, 0, -5.139921e-21, 5.139921e-21, -5.139921e-21, 
    -3.597945e-20, -1.027984e-20, -5.139921e-21, -2.006177e-36, 2.006177e-36, 
    -1.541976e-20, -1.027984e-20, -2.055969e-20, -1.541976e-20, 1.027984e-20, 
    5.139921e-21, -1.027984e-20, -5.139921e-21, 1.027984e-20, -5.139921e-21, 
    5.139921e-21, -5.139921e-21, -1.027984e-20, 2.055969e-20, 5.139921e-21, 
    -1.541976e-20, -1.541976e-20, -5.139921e-21, 3.597945e-20, -1.541976e-20, 
    1.541976e-20, 1.541976e-20, 1.541976e-20, -2.055969e-20, -2.006177e-36, 
    -3.597945e-20, 5.139921e-21, -1.027984e-20, 3.083953e-20, 2.055969e-20, 
    0, 5.139921e-21, -2.569961e-20, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 2.006177e-36, 5.139921e-21, -5.139921e-21, 0, 
    -2.569961e-20, 3.083953e-20, -4.111937e-20, -1.541976e-20, 1.027984e-20, 
    1.027984e-20, -2.055969e-20, 1.027984e-20, 0, 5.139921e-21, 1.027984e-20, 
    -5.139921e-21, -1.027984e-20, -2.569961e-20, 5.139921e-21, -2.006177e-36, 
    -2.055969e-20, 1.027984e-20, 1.027984e-20, -1.027984e-20, 5.139921e-21, 
    -3.597945e-20, 1.027984e-20, -2.006177e-36, 5.139921e-21, 5.139921e-21, 
    1.541976e-20, 0, -1.541976e-20, -1.541976e-20, 1.541976e-20, 1.027984e-20,
  -1.027984e-20, 1.027984e-20, -5.139921e-21, -2.569961e-20, -5.139921e-21, 
    -1.027984e-20, -5.139921e-21, -1.541976e-20, 1.541976e-20, 4.111937e-20, 
    5.139921e-21, 1.541976e-20, 2.006177e-36, -5.139921e-21, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, 3.083953e-20, -1.027984e-20, 1.541976e-20, 
    1.027984e-20, 1.541976e-20, -1.027984e-20, 0, 5.139921e-21, 
    -2.006177e-36, -2.006177e-36, -1.027984e-20, 0, -5.139921e-21, 
    -1.027984e-20, 3.597945e-20, -5.139921e-21, -1.541976e-20, -5.139921e-21, 
    -2.569961e-20, -5.139921e-21, 2.055969e-20, 1.027984e-20, 0, 
    1.541976e-20, -1.541976e-20, -2.569961e-20, -2.569961e-20, 0, 
    -5.139921e-21, -2.569961e-20, 1.027984e-20, -2.569961e-20, -2.569961e-20, 
    5.139921e-21, 0, 3.597945e-20, -2.569961e-20, 5.139921e-21, 
    -1.027984e-20, -5.139921e-21, 1.027984e-20, -1.027984e-20, 5.139921e-21, 
    0, -5.139921e-21, 5.139921e-21, -5.139921e-21, -1.541976e-20, 
    2.055969e-20, -1.027984e-20, -1.541976e-20, -2.055969e-20, 2.006177e-36, 
    -3.597945e-20, -1.027984e-20, -2.055969e-20, 1.027984e-20, -1.027984e-20, 
    -2.006177e-36, -1.541976e-20, 2.055969e-20, -5.139921e-21, -5.139921e-21, 
    -1.027984e-20, -3.083953e-20, -1.541976e-20, 2.006177e-36, 1.541976e-20, 
    5.139921e-21, 0, 1.027984e-20, 3.083953e-20, -2.055969e-20, 1.541976e-20, 
    0, 5.139921e-21, -3.083953e-20, -5.139921e-21, 1.541976e-20, 
    5.139921e-21, -5.139921e-21, 1.541976e-20, -3.083953e-20, 1.027984e-20, 
    5.139921e-21, -5.139921e-21, 0, 0, 1.027984e-20, 5.139921e-21, 
    -5.139921e-21, 2.569961e-20, 1.541976e-20, -1.027984e-20, 1.541976e-20, 
    0, -1.027984e-20, -2.006177e-36, 5.139921e-21, 1.027984e-20, 
    2.055969e-20, 0, 5.139921e-21, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, 3.597945e-20, 1.541976e-20, -1.541976e-20, -5.139921e-21, 
    -5.139921e-21, -1.541976e-20, -2.569961e-20, -1.541976e-20, 
    -5.139921e-21, 2.055969e-20, -2.055969e-20, -5.139921e-21, 1.541976e-20, 
    5.139921e-21, -1.541976e-20, 5.139921e-21, 1.541976e-20, -5.139921e-21, 
    -1.541976e-20, 0, 1.541976e-20, 5.139921e-21, 1.541976e-20, 0, 
    -5.139921e-21, 2.055969e-20, -1.027984e-20, 0, 1.541976e-20, 
    -2.055969e-20, 0, -1.027984e-20, -2.569961e-20, 5.139921e-21, 
    -1.541976e-20, 1.027984e-20, 2.055969e-20, 0, -1.027984e-20, 
    3.083953e-20, 5.139921e-21, -1.027984e-20, -2.055969e-20, 0, 
    -5.139921e-21, -2.055969e-20, -1.541976e-20, -2.055969e-20, 
    -3.083953e-20, 1.027984e-20, 2.569961e-20, 2.055969e-20, -2.055969e-20, 
    1.027984e-20, 1.027984e-20, -1.541976e-20, 3.083953e-20, -1.027984e-20, 
    -2.055969e-20, -5.139921e-21, -1.541976e-20, 3.597945e-20, 0, 0, 
    -1.541976e-20, 5.139921e-21, 3.083953e-20, 2.569961e-20, -5.139921e-21, 
    2.055969e-20, -2.055969e-20, -5.139921e-21, -4.111937e-20, 1.541976e-20, 
    5.139921e-21, 1.027984e-20, 1.027984e-20, -2.006177e-36, 5.139921e-21, 
    1.027984e-20, -1.027984e-20, -5.139921e-21, 1.027984e-20, 1.027984e-20, 
    1.027984e-20, -5.139921e-21, 1.541976e-20, -1.027984e-20, 3.083953e-20, 
    1.027984e-20, 2.055969e-20, -5.139921e-21, 0, -4.111937e-20, 
    1.541976e-20, -2.055969e-20, -1.541976e-20, 0, 5.139921e-21, 
    1.027984e-20, 2.055969e-20, 1.541976e-20, -2.006177e-36, 1.027984e-20, 
    5.139921e-21, 5.139921e-21, -2.569961e-20, -5.139921e-21, -3.083953e-20, 
    0, -1.541976e-20, 5.139921e-21, 5.139921e-21, 1.027984e-20, 5.139921e-21, 
    2.055969e-20, 2.055969e-20, 2.006177e-36, 1.027984e-20, 0, -2.569961e-20, 
    -5.139921e-21, 5.139921e-21, -2.006177e-36, -2.569961e-20, -2.055969e-20, 
    -1.027984e-20, 1.027984e-20, 2.569961e-20, 1.541976e-20, -2.569961e-20, 
    5.139921e-21, -5.139921e-21, 0, 1.027984e-20, -1.541976e-20, 
    5.139921e-21, 5.139921e-21, -5.139921e-21, -5.139921e-21, 1.027984e-20, 
    -5.139921e-21, 2.055969e-20, -5.139921e-21, 2.006177e-36, 0, 
    -5.139921e-21, 1.541976e-20, -5.139921e-21, 5.139921e-21, -2.569961e-20, 
    -2.569961e-20, 1.027984e-20, 5.139921e-21, 1.541976e-20, -2.006177e-36, 
    -5.139921e-21, -2.055969e-20, 3.597945e-20, -1.027984e-20, -1.027984e-20, 
    5.139921e-21, -2.055969e-20, 1.027984e-20, -2.055969e-20, 1.027984e-20, 
    5.139921e-21, -5.139921e-21, 5.139921e-21, 2.055969e-20, 2.055969e-20, 
    -1.027984e-20, 1.541976e-20, -2.006177e-36, -5.139921e-21, -1.027984e-20, 
    1.027984e-20, 5.139921e-21, -2.569961e-20, -2.569961e-20, 1.541976e-20, 
    3.597945e-20, -1.027984e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -2.055969e-20, 0, 0, -5.139921e-21, 2.055969e-20, 0, -5.139921e-21, 
    5.139921e-21, -1.541976e-20, -1.027984e-20, -3.083953e-20, -5.139921e-21, 
    1.027984e-20, 1.027984e-20, 1.541976e-20, -5.139921e-21, -5.139921e-21, 
    2.055969e-20, -2.055969e-20, 2.006177e-36, 5.139921e-21, -1.541976e-20, 
    -2.006177e-36, 1.027984e-20, 1.027984e-20, 2.006177e-36, 3.597945e-20, 
    1.027984e-20, 2.055969e-20,
  -5.139921e-21, -5.139921e-21, -5.139921e-21, -3.083953e-20, -1.541976e-20, 
    -5.139921e-21, 1.027984e-20, 2.055969e-20, 7.709882e-20, -1.027984e-20, 
    -1.027984e-20, 0, -1.541976e-20, 1.541976e-20, 1.541976e-20, 
    -3.083953e-20, 2.055969e-20, 1.541976e-20, 2.055969e-20, -1.541976e-20, 
    -2.569961e-20, -1.027984e-20, -3.597945e-20, 1.541976e-20, 1.027984e-20, 
    -5.139921e-21, 1.027984e-20, 0, -5.139921e-21, 1.541976e-20, 
    1.541976e-20, 1.027984e-20, -5.139921e-21, -2.055969e-20, -2.055969e-20, 
    5.139921e-21, 1.541976e-20, 1.027984e-20, -3.597945e-20, -5.139921e-21, 
    1.541976e-20, -5.139921e-21, -5.139921e-21, 2.569961e-20, 1.541976e-20, 
    2.569961e-20, 3.083953e-20, -1.541976e-20, -1.541976e-20, 1.027984e-20, 
    -2.055969e-20, -1.541976e-20, -1.027984e-20, 2.569961e-20, -2.055969e-20, 
    -2.569961e-20, -1.027984e-20, -2.055969e-20, -3.597945e-20, 
    -5.139921e-21, -1.027984e-20, -3.597945e-20, -5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 1.027984e-20, 3.597945e-20, -1.541976e-20, 
    -4.111937e-20, 2.569961e-20, -2.569961e-20, -5.139921e-21, -2.055969e-20, 
    -2.055969e-20, 5.139921e-21, -4.111937e-20, 3.083953e-20, -3.597945e-20, 
    -2.006177e-36, -1.541976e-20, 5.139921e-21, 1.027984e-20, -3.083953e-20, 
    -2.055969e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, -1.027984e-20, 
    2.055969e-20, 2.569961e-20, -2.055969e-20, -1.027984e-20, -2.055969e-20, 
    1.541976e-20, -1.541976e-20, -1.027984e-20, -1.027984e-20, -5.139921e-21, 
    3.083953e-20, -1.027984e-20, -5.139921e-21, -5.139921e-21, -1.541976e-20, 
    1.027984e-20, 2.569961e-20, -2.055969e-20, -2.055969e-20, -1.027984e-20, 
    5.653913e-20, -3.083953e-20, 5.139921e-21, 1.027984e-20, -1.027984e-20, 
    -2.569961e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, 2.006177e-36, 
    -2.055969e-20, -5.139921e-21, -1.541976e-20, -1.027984e-20, 5.139921e-21, 
    -2.055969e-20, -5.139921e-21, -1.027984e-20, 5.139921e-21, -1.027984e-20, 
    -3.083953e-20, -2.006177e-36, -5.139921e-21, -2.055969e-20, 1.027984e-20, 
    -5.139921e-21, 1.541976e-20, 2.055969e-20, -1.027984e-20, -1.027984e-20, 
    -3.597945e-20, -2.055969e-20, -1.027984e-20, 5.139921e-21, 5.139921e-21, 
    -2.006177e-36, 5.139921e-21, 1.541976e-20, 1.027984e-20, 5.139921e-21, 
    -2.055969e-20, -5.139921e-21, -2.055969e-20, 3.597945e-20, -5.139921e-21, 
    -1.027984e-20, 4.111937e-20, 5.139921e-21, 5.139921e-21, 4.111937e-20, 
    5.139921e-21, -1.541976e-20, 5.139921e-21, -1.027984e-20, 5.139921e-21, 
    1.027984e-20, 3.083953e-20, 0, 4.111937e-20, 2.055969e-20, -2.006177e-36, 
    0, 1.541976e-20, -1.027984e-20, 1.027984e-20, 2.055969e-20, 0, 
    1.027984e-20, -2.055969e-20, 2.569961e-20, 2.055969e-20, 0, 
    -3.597945e-20, -5.139921e-21, 1.027984e-20, 1.027984e-20, 5.139921e-21, 
    3.597945e-20, -5.139921e-21, -1.541976e-20, 2.569961e-20, -5.139921e-21, 
    5.139921e-21, -2.055969e-20, 5.139921e-21, -5.139921e-20, 1.027984e-20, 
    -5.139921e-21, 1.027984e-20, 1.027984e-20, -5.139921e-21, 3.083953e-20, 
    -2.569961e-20, 1.541976e-20, -2.006177e-36, 5.139921e-21, 5.139921e-21, 
    -5.139921e-21, 5.139921e-21, 3.083953e-20, -5.139921e-21, -1.541976e-20, 
    -1.027984e-20, 2.569961e-20, 1.541976e-20, 0, 2.055969e-20, 2.569961e-20, 
    3.083953e-20, -5.139921e-21, -1.027984e-20, -1.027984e-20, -5.139921e-21, 
    2.569961e-20, 1.541976e-20, 5.139921e-21, 1.027984e-20, 4.111937e-20, 
    5.139921e-21, 5.139921e-21, -2.569961e-20, 2.569961e-20, -5.139921e-21, 
    -1.541976e-20, -2.569961e-20, 2.055969e-20, -3.597945e-20, 1.541976e-20, 
    1.027984e-20, -1.541976e-20, -5.139921e-21, 1.541976e-20, -1.027984e-20, 
    -5.139921e-21, -5.139921e-21, 2.569961e-20, -2.006177e-36, 1.541976e-20, 
    1.027984e-20, -2.055969e-20, 5.139921e-21, 1.027984e-20, -1.027984e-20, 
    -4.111937e-20, 5.139921e-21, -5.139921e-21, -1.541976e-20, -1.027984e-20, 
    2.055969e-20, 3.597945e-20, 1.541976e-20, 1.541976e-20, 5.139921e-21, 
    -2.055969e-20, 3.597945e-20, -1.027984e-20, -3.083953e-20, 2.006177e-36, 
    -3.083953e-20, 5.139921e-21, -4.625929e-20, 3.083953e-20, -1.541976e-20, 
    1.027984e-20, -5.139921e-21, 1.027984e-20, -1.541976e-20, 1.541976e-20, 
    2.569961e-20, -1.027984e-20, 2.055969e-20, -2.055969e-20, -2.055969e-20, 
    -5.139921e-21, 1.027984e-20, 3.597945e-20, 2.569961e-20, -2.055969e-20, 
    3.083953e-20, 1.027984e-20, -1.027984e-20, -2.569961e-20, -5.139921e-21, 
    -5.139921e-21, -1.027984e-20, 2.569961e-20, 5.139921e-21, 1.541976e-20, 
    1.027984e-20, -3.597945e-20, 0, -2.569961e-20, 5.139921e-21, 0, 
    2.006177e-36, 1.027984e-20, -2.006177e-36, 2.055969e-20, 5.139921e-21, 
    2.055969e-20, -2.055969e-20, -1.027984e-20, -2.055969e-20, 1.027984e-20, 
    1.027984e-20, 0, 1.541976e-20, 5.139921e-21, -1.541976e-20, 0, 
    3.597945e-20, -1.541976e-20, -2.569961e-20, 2.569961e-20, 1.027984e-20, 
    5.139921e-21, 0, -1.541976e-20, 0, 1.541976e-20, 2.569961e-20, 
    -1.541976e-20, -5.139921e-21, 1.027984e-20, 5.139921e-21, 0, 
    -2.055969e-20, 2.569961e-20, -5.139921e-21, 3.083953e-20,
  1.027984e-20, 5.139921e-21, 1.541976e-20, -3.083953e-20, -2.055969e-20, 
    3.083953e-20, -5.139921e-21, -2.006177e-36, -5.139921e-21, -2.055969e-20, 
    -5.139921e-21, 1.541976e-20, -2.569961e-20, -2.055969e-20, -5.139921e-21, 
    -1.541976e-20, 5.139921e-21, 1.541976e-20, -2.055969e-20, -2.055969e-20, 
    -2.055969e-20, 1.027984e-20, 1.027984e-20, -2.006177e-36, 2.569961e-20, 
    -1.027984e-20, -2.055969e-20, -1.541976e-20, 2.055969e-20, 1.027984e-20, 
    1.541976e-20, 0, 2.055969e-20, 1.541976e-20, 1.541976e-20, 1.541976e-20, 
    -2.055969e-20, -2.055969e-20, 3.597945e-20, 1.027984e-20, -5.139921e-21, 
    5.139921e-21, 1.027984e-20, -2.055969e-20, 2.055969e-20, -1.027984e-20, 
    3.597945e-20, -2.569961e-20, -1.541976e-20, 1.027984e-20, 0, 
    -3.597945e-20, -2.055969e-20, -1.541976e-20, 5.139921e-21, 0, 
    2.569961e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    3.083953e-20, 0, 2.006177e-36, 1.027984e-20, 1.541976e-20, 1.027984e-20, 
    0, 2.569961e-20, 3.597945e-20, 1.541976e-20, -3.597945e-20, 
    -5.139921e-21, -1.541976e-20, -1.027984e-20, 2.569961e-20, 5.139921e-21, 
    -5.139921e-21, -1.027984e-20, -1.027984e-20, 5.139921e-21, -1.541976e-20, 
    -1.027984e-20, 0, -5.139921e-21, -2.006177e-36, -3.083953e-20, 
    -1.541976e-20, -1.541976e-20, 1.027984e-20, -3.083953e-20, 2.055969e-20, 
    5.139921e-21, 5.139921e-21, 2.055969e-20, 2.569961e-20, 5.139921e-21, 
    2.569961e-20, 0, -1.027984e-20, 1.541976e-20, -5.139921e-21, 
    1.541976e-20, 1.027984e-20, 5.139921e-21, -1.541976e-20, 2.006177e-36, 0, 
    -5.139921e-21, -5.139921e-21, 0, 1.541976e-20, 1.027984e-20, 
    2.569961e-20, 2.569961e-20, 5.139921e-21, 5.139921e-21, 1.027984e-20, 
    -2.006177e-36, -1.027984e-20, 1.027984e-20, 4.625929e-20, -2.569961e-20, 
    -5.139921e-21, -2.055969e-20, -5.139921e-21, 1.541976e-20, -5.139921e-21, 
    -2.055969e-20, -1.541976e-20, -2.055969e-20, 5.139921e-21, 0, 
    5.139921e-21, 5.139921e-21, -3.597945e-20, -1.541976e-20, 1.541976e-20, 
    3.083953e-20, -1.027984e-20, -1.027984e-20, 4.625929e-20, -1.027984e-20, 
    2.055969e-20, 1.541976e-20, 5.139921e-21, 1.541976e-20, 1.027984e-20, 0, 
    -2.055969e-20, 2.055969e-20, -3.597945e-20, 2.006177e-36, -3.597945e-20, 
    1.541976e-20, 1.541976e-20, -1.027984e-20, -2.055969e-20, -1.541976e-20, 
    -5.139921e-21, 5.139921e-21, 1.541976e-20, 1.541976e-20, -1.027984e-20, 
    0, 2.569961e-20, 3.597945e-20, 0, 2.006177e-36, 0, 3.597945e-20, 0, 
    -2.569961e-20, -5.139921e-21, -1.027984e-20, 1.027984e-20, 2.055969e-20, 
    -5.139921e-21, -1.541976e-20, -1.541976e-20, 1.541976e-20, -5.139921e-21, 
    -3.597945e-20, 1.027984e-20, 2.055969e-20, 4.111937e-20, -5.139921e-21, 
    5.139921e-21, -1.027984e-20, 1.541976e-20, -1.027984e-20, 0, 
    -5.139921e-21, 2.055969e-20, 2.006177e-36, -5.139921e-21, 2.055969e-20, 
    -3.083953e-20, 1.541976e-20, -4.111937e-20, 2.569961e-20, 1.541976e-20, 
    -2.055969e-20, 1.027984e-20, 1.027984e-20, -1.027984e-20, -2.006177e-36, 
    2.006177e-36, -2.006177e-36, 1.027984e-20, -3.597945e-20, 2.055969e-20, 
    1.027984e-20, -5.653913e-20, -1.541976e-20, -5.139921e-21, 1.541976e-20, 
    -4.111937e-20, 5.139921e-21, -2.569961e-20, 2.006177e-36, 0, 
    2.055969e-20, 1.541976e-20, -2.569961e-20, 0, 5.139921e-21, 1.541976e-20, 
    1.541976e-20, -1.027984e-20, -2.055969e-20, 2.006177e-36, -1.027984e-20, 
    5.139921e-21, -2.055969e-20, 1.027984e-20, -1.541976e-20, 5.139921e-21, 
    -5.139921e-21, 2.055969e-20, 1.027984e-20, 2.055969e-20, -2.569961e-20, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, -2.055969e-20, -1.541976e-20, 
    -3.083953e-20, -1.027984e-20, -5.139921e-21, 5.139921e-21, 0, 
    1.541976e-20, 0, 5.139921e-21, 2.569961e-20, -1.541976e-20, 
    -1.027984e-20, 1.541976e-20, 1.541976e-20, 0, -1.027984e-20, 
    5.139921e-21, 2.006177e-36, -3.597945e-20, 5.139921e-21, -5.139921e-21, 
    1.027984e-20, -5.139921e-21, -5.139921e-21, -1.027984e-20, -4.625929e-20, 
    -2.055969e-20, 2.006177e-36, -5.139921e-21, 0, -5.139921e-21, 
    5.139921e-21, 5.139921e-21, 0, 2.006177e-36, 5.139921e-21, -2.006177e-36, 
    2.569961e-20, -3.083953e-20, 0, 1.541976e-20, -1.541976e-20, 
    2.055969e-20, 1.027984e-20, -1.027984e-20, -5.139921e-21, -2.006177e-36, 
    -2.569961e-20, -1.027984e-20, 2.055969e-20, -1.541976e-20, -5.139921e-21, 
    2.006177e-36, 5.139921e-21, 1.541976e-20, -1.541976e-20, 2.055969e-20, 
    5.139921e-21, 2.055969e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, 
    2.055969e-20, -2.055969e-20, -2.006177e-36, -1.027984e-20, 1.027984e-20, 
    -5.139921e-21, 2.569961e-20, -1.541976e-20, 5.139921e-21, 2.569961e-20, 
    -2.055969e-20, 5.139921e-21, 0, -2.055969e-20, -5.139921e-21, 
    1.027984e-20, 3.083953e-20, 1.027984e-20, 1.027984e-20, -5.139921e-21, 
    1.027984e-20, -2.055969e-20, 5.139921e-21, 2.055969e-20, 1.541976e-20, 
    2.006177e-36, 1.027984e-20, -5.139921e-21, 2.569961e-20,
  8.59741e-29, 8.59739e-29, 8.597394e-29, 8.597377e-29, 8.597386e-29, 
    8.597375e-29, 8.597406e-29, 8.597389e-29, 8.5974e-29, 8.597408e-29, 
    8.597344e-29, 8.597376e-29, 8.597311e-29, 8.597331e-29, 8.59728e-29, 
    8.597315e-29, 8.597274e-29, 8.597281e-29, 8.597258e-29, 8.597265e-29, 
    8.597235e-29, 8.597255e-29, 8.597219e-29, 8.597239e-29, 8.597236e-29, 
    8.597256e-29, 8.59737e-29, 8.597348e-29, 8.597371e-29, 8.597368e-29, 
    8.597369e-29, 8.597386e-29, 8.597395e-29, 8.597412e-29, 8.597409e-29, 
    8.597396e-29, 8.597366e-29, 8.597377e-29, 8.597351e-29, 8.597352e-29, 
    8.597324e-29, 8.597337e-29, 8.59729e-29, 8.597303e-29, 8.597265e-29, 
    8.597274e-29, 8.597265e-29, 8.597268e-29, 8.597265e-29, 8.597279e-29, 
    8.597273e-29, 8.597286e-29, 8.597334e-29, 8.59732e-29, 8.597363e-29, 
    8.597389e-29, 8.597405e-29, 8.597417e-29, 8.597416e-29, 8.597413e-29, 
    8.597396e-29, 8.59738e-29, 8.597368e-29, 8.59736e-29, 8.597352e-29, 
    8.597328e-29, 8.597315e-29, 8.597287e-29, 8.597292e-29, 8.597283e-29, 
    8.597275e-29, 8.597261e-29, 8.597263e-29, 8.597257e-29, 8.597283e-29, 
    8.597266e-29, 8.597295e-29, 8.597287e-29, 8.59735e-29, 8.597374e-29, 
    8.597384e-29, 8.597393e-29, 8.597414e-29, 8.597399e-29, 8.597405e-29, 
    8.597392e-29, 8.597383e-29, 8.597387e-29, 8.59736e-29, 8.597371e-29, 
    8.597315e-29, 8.597339e-29, 8.597276e-29, 8.597291e-29, 8.597272e-29, 
    8.597282e-29, 8.597266e-29, 8.59728e-29, 8.597255e-29, 8.59725e-29, 
    8.597253e-29, 8.597239e-29, 8.597281e-29, 8.597265e-29, 8.597387e-29, 
    8.597386e-29, 8.597383e-29, 8.597398e-29, 8.597399e-29, 8.597412e-29, 
    8.5974e-29, 8.597395e-29, 8.597382e-29, 8.597374e-29, 8.597367e-29, 
    8.597351e-29, 8.597333e-29, 8.597308e-29, 8.59729e-29, 8.597278e-29, 
    8.597285e-29, 8.597279e-29, 8.597286e-29, 8.597289e-29, 8.597251e-29, 
    8.597273e-29, 8.597241e-29, 8.597242e-29, 8.597257e-29, 8.597242e-29, 
    8.597386e-29, 8.59739e-29, 8.597404e-29, 8.597393e-29, 8.597414e-29, 
    8.597402e-29, 8.597396e-29, 8.59737e-29, 8.597365e-29, 8.597359e-29, 
    8.597349e-29, 8.597336e-29, 8.597313e-29, 8.597293e-29, 8.597274e-29, 
    8.597276e-29, 8.597275e-29, 8.597271e-29, 8.597281e-29, 8.597269e-29, 
    8.597268e-29, 8.597273e-29, 8.597243e-29, 8.597251e-29, 8.597242e-29, 
    8.597248e-29, 8.597389e-29, 8.597382e-29, 8.597386e-29, 8.597378e-29, 
    8.597383e-29, 8.597362e-29, 8.597355e-29, 8.597324e-29, 8.597336e-29, 
    8.597316e-29, 8.597334e-29, 8.597331e-29, 8.597315e-29, 8.597333e-29, 
    8.597294e-29, 8.597321e-29, 8.597271e-29, 8.597298e-29, 8.597269e-29, 
    8.597275e-29, 8.597266e-29, 8.597259e-29, 8.597249e-29, 8.597232e-29, 
    8.597235e-29, 8.597221e-29, 8.597371e-29, 8.597362e-29, 8.597363e-29, 
    8.597354e-29, 8.597346e-29, 8.597331e-29, 8.597307e-29, 8.597316e-29, 
    8.5973e-29, 8.597296e-29, 8.597322e-29, 8.597306e-29, 8.597356e-29, 
    8.597348e-29, 8.597353e-29, 8.597371e-29, 8.597314e-29, 8.597343e-29, 
    8.59729e-29, 8.597306e-29, 8.59726e-29, 8.597283e-29, 8.597238e-29, 
    8.597218e-29, 8.5972e-29, 8.597179e-29, 8.597357e-29, 8.597363e-29, 
    8.597352e-29, 8.597337e-29, 8.597323e-29, 8.597304e-29, 8.597303e-29, 
    8.597299e-29, 8.59729e-29, 8.597282e-29, 8.597298e-29, 8.59728e-29, 
    8.597346e-29, 8.597312e-29, 8.597366e-29, 8.597349e-29, 8.597338e-29, 
    8.597343e-29, 8.597318e-29, 8.597312e-29, 8.597286e-29, 8.5973e-29, 
    8.597223e-29, 8.597257e-29, 8.597163e-29, 8.597189e-29, 8.597366e-29, 
    8.597357e-29, 8.597328e-29, 8.597342e-29, 8.597303e-29, 8.597293e-29, 
    8.597286e-29, 8.597275e-29, 8.597275e-29, 8.597269e-29, 8.597278e-29, 
    8.597269e-29, 8.597304e-29, 8.597289e-29, 8.597332e-29, 8.597321e-29, 
    8.597326e-29, 8.597331e-29, 8.597315e-29, 8.597298e-29, 8.597297e-29, 
    8.597292e-29, 8.597276e-29, 8.597303e-29, 8.597219e-29, 8.597271e-29, 
    8.597348e-29, 8.597333e-29, 8.59733e-29, 8.597336e-29, 8.597295e-29, 
    8.59731e-29, 8.597269e-29, 8.59728e-29, 8.597262e-29, 8.597271e-29, 
    8.597272e-29, 8.597284e-29, 8.597291e-29, 8.597309e-29, 8.597324e-29, 
    8.597336e-29, 8.597333e-29, 8.59732e-29, 8.597297e-29, 8.597274e-29, 
    8.597279e-29, 8.597263e-29, 8.597306e-29, 8.597288e-29, 8.597295e-29, 
    8.597277e-29, 8.597316e-29, 8.597283e-29, 8.597325e-29, 8.597322e-29, 
    8.59731e-29, 8.597287e-29, 8.597281e-29, 8.597276e-29, 8.59728e-29, 
    8.597296e-29, 8.597299e-29, 8.59731e-29, 8.597313e-29, 8.597322e-29, 
    8.59733e-29, 8.597323e-29, 8.597316e-29, 8.597296e-29, 8.597278e-29, 
    8.597259e-29, 8.597254e-29, 8.597231e-29, 8.59725e-29, 8.597218e-29, 
    8.597245e-29, 8.5972e-29, 8.597281e-29, 8.597245e-29, 8.59731e-29, 
    8.597303e-29, 8.59729e-29, 8.597262e-29, 8.597277e-29, 8.597259e-29, 
    8.597299e-29, 8.597319e-29, 8.597325e-29, 8.597335e-29, 8.597325e-29, 
    8.597325e-29, 8.597316e-29, 8.597319e-29, 8.597295e-29, 8.597308e-29, 
    8.597272e-29, 8.597259e-29, 8.597222e-29, 8.5972e-29, 8.597176e-29, 
    8.597167e-29, 8.597163e-29, 8.597162e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N_TO_SOIL2N =
  1.397129e-08, 1.400952e-08, 1.400209e-08, 1.403292e-08, 1.401582e-08, 
    1.4036e-08, 1.397904e-08, 1.401103e-08, 1.399061e-08, 1.397473e-08, 
    1.409272e-08, 1.403429e-08, 1.415341e-08, 1.411616e-08, 1.420971e-08, 
    1.414761e-08, 1.422224e-08, 1.420793e-08, 1.4251e-08, 1.423866e-08, 
    1.429372e-08, 1.425669e-08, 1.432226e-08, 1.428488e-08, 1.429073e-08, 
    1.425547e-08, 1.404606e-08, 1.408544e-08, 1.404372e-08, 1.404934e-08, 
    1.404682e-08, 1.401617e-08, 1.400072e-08, 1.396837e-08, 1.397424e-08, 
    1.3998e-08, 1.405187e-08, 1.403359e-08, 1.407966e-08, 1.407862e-08, 
    1.412989e-08, 1.410678e-08, 1.419293e-08, 1.416845e-08, 1.423918e-08, 
    1.422139e-08, 1.423834e-08, 1.42332e-08, 1.423841e-08, 1.421232e-08, 
    1.42235e-08, 1.420055e-08, 1.41111e-08, 1.413739e-08, 1.405897e-08, 
    1.401178e-08, 1.398044e-08, 1.39582e-08, 1.396134e-08, 1.396734e-08, 
    1.399814e-08, 1.402711e-08, 1.404917e-08, 1.406393e-08, 1.407847e-08, 
    1.412246e-08, 1.414575e-08, 1.419787e-08, 1.418847e-08, 1.42044e-08, 
    1.421962e-08, 1.424517e-08, 1.424096e-08, 1.425222e-08, 1.420398e-08, 
    1.423604e-08, 1.418312e-08, 1.419759e-08, 1.40824e-08, 1.403852e-08, 
    1.401985e-08, 1.400352e-08, 1.396376e-08, 1.399121e-08, 1.398039e-08, 
    1.400614e-08, 1.40225e-08, 1.401441e-08, 1.406433e-08, 1.404493e-08, 
    1.414713e-08, 1.410312e-08, 1.421785e-08, 1.41904e-08, 1.422443e-08, 
    1.420707e-08, 1.423681e-08, 1.421004e-08, 1.425641e-08, 1.42665e-08, 
    1.42596e-08, 1.42861e-08, 1.420856e-08, 1.423834e-08, 1.401418e-08, 
    1.40155e-08, 1.402165e-08, 1.399462e-08, 1.399297e-08, 1.396821e-08, 
    1.399024e-08, 1.399963e-08, 1.402345e-08, 1.403754e-08, 1.405093e-08, 
    1.408036e-08, 1.411323e-08, 1.415918e-08, 1.419218e-08, 1.42143e-08, 
    1.420074e-08, 1.421271e-08, 1.419933e-08, 1.419305e-08, 1.426272e-08, 
    1.42236e-08, 1.428229e-08, 1.427904e-08, 1.425248e-08, 1.427941e-08, 
    1.401643e-08, 1.400884e-08, 1.398247e-08, 1.40031e-08, 1.396551e-08, 
    1.398655e-08, 1.399865e-08, 1.404533e-08, 1.405559e-08, 1.406509e-08, 
    1.408387e-08, 1.410796e-08, 1.415021e-08, 1.418696e-08, 1.422051e-08, 
    1.421805e-08, 1.421892e-08, 1.422641e-08, 1.420785e-08, 1.422945e-08, 
    1.423308e-08, 1.42236e-08, 1.427861e-08, 1.426289e-08, 1.427897e-08, 
    1.426874e-08, 1.401131e-08, 1.402408e-08, 1.401718e-08, 1.403016e-08, 
    1.402101e-08, 1.406167e-08, 1.407386e-08, 1.413088e-08, 1.410748e-08, 
    1.414472e-08, 1.411127e-08, 1.41172e-08, 1.414592e-08, 1.411308e-08, 
    1.418493e-08, 1.413621e-08, 1.42267e-08, 1.417805e-08, 1.422975e-08, 
    1.422036e-08, 1.42359e-08, 1.424981e-08, 1.426731e-08, 1.429959e-08, 
    1.429212e-08, 1.431911e-08, 1.404313e-08, 1.405969e-08, 1.405823e-08, 
    1.407557e-08, 1.408839e-08, 1.411617e-08, 1.416072e-08, 1.414397e-08, 
    1.417472e-08, 1.418089e-08, 1.413418e-08, 1.416285e-08, 1.407078e-08, 
    1.408565e-08, 1.40768e-08, 1.404443e-08, 1.414782e-08, 1.409477e-08, 
    1.419273e-08, 1.4164e-08, 1.424783e-08, 1.420614e-08, 1.4288e-08, 
    1.432297e-08, 1.43559e-08, 1.439434e-08, 1.406873e-08, 1.405748e-08, 
    1.407763e-08, 1.410551e-08, 1.413137e-08, 1.416575e-08, 1.416927e-08, 
    1.417571e-08, 1.419238e-08, 1.42064e-08, 1.417774e-08, 1.420992e-08, 
    1.40891e-08, 1.415243e-08, 1.405322e-08, 1.40831e-08, 1.410386e-08, 
    1.409476e-08, 1.414206e-08, 1.41532e-08, 1.419847e-08, 1.417507e-08, 
    1.431434e-08, 1.425274e-08, 1.442362e-08, 1.437589e-08, 1.405354e-08, 
    1.40687e-08, 1.412141e-08, 1.409633e-08, 1.416805e-08, 1.418569e-08, 
    1.420004e-08, 1.421837e-08, 1.422035e-08, 1.423121e-08, 1.421341e-08, 
    1.423051e-08, 1.416582e-08, 1.419473e-08, 1.411539e-08, 1.41347e-08, 
    1.412582e-08, 1.411607e-08, 1.414615e-08, 1.417819e-08, 1.417888e-08, 
    1.418915e-08, 1.421807e-08, 1.416834e-08, 1.432228e-08, 1.422722e-08, 
    1.408521e-08, 1.411438e-08, 1.411856e-08, 1.410726e-08, 1.418392e-08, 
    1.415615e-08, 1.423094e-08, 1.421073e-08, 1.424385e-08, 1.422739e-08, 
    1.422497e-08, 1.420384e-08, 1.419068e-08, 1.415742e-08, 1.413036e-08, 
    1.41089e-08, 1.411389e-08, 1.413746e-08, 1.418015e-08, 1.422052e-08, 
    1.421168e-08, 1.424133e-08, 1.416285e-08, 1.419576e-08, 1.418304e-08, 
    1.421621e-08, 1.414352e-08, 1.42054e-08, 1.41277e-08, 1.413452e-08, 
    1.41556e-08, 1.419799e-08, 1.420737e-08, 1.421738e-08, 1.421121e-08, 
    1.418123e-08, 1.417632e-08, 1.415509e-08, 1.414922e-08, 1.413303e-08, 
    1.411963e-08, 1.413187e-08, 1.414473e-08, 1.418125e-08, 1.421415e-08, 
    1.425001e-08, 1.425878e-08, 1.430065e-08, 1.426656e-08, 1.432281e-08, 
    1.427498e-08, 1.435777e-08, 1.4209e-08, 1.427358e-08, 1.415656e-08, 
    1.416917e-08, 1.419198e-08, 1.424428e-08, 1.421605e-08, 1.424907e-08, 
    1.417613e-08, 1.413827e-08, 1.412848e-08, 1.41102e-08, 1.41289e-08, 
    1.412738e-08, 1.414527e-08, 1.413952e-08, 1.418246e-08, 1.41594e-08, 
    1.422491e-08, 1.424881e-08, 1.431628e-08, 1.435763e-08, 1.439971e-08, 
    1.441828e-08, 1.442393e-08, 1.44263e-08 ;

 SOIL1N_TO_SOIL3N =
  1.657483e-10, 1.662021e-10, 1.661139e-10, 1.664798e-10, 1.662768e-10, 
    1.665164e-10, 1.658403e-10, 1.6622e-10, 1.659776e-10, 1.657892e-10, 
    1.671896e-10, 1.664961e-10, 1.679099e-10, 1.674678e-10, 1.685783e-10, 
    1.678411e-10, 1.687269e-10, 1.685571e-10, 1.690683e-10, 1.689219e-10, 
    1.695754e-10, 1.691359e-10, 1.699142e-10, 1.694705e-10, 1.695399e-10, 
    1.691214e-10, 1.666357e-10, 1.671032e-10, 1.66608e-10, 1.666747e-10, 
    1.666448e-10, 1.66281e-10, 1.660976e-10, 1.657136e-10, 1.657833e-10, 
    1.660654e-10, 1.667047e-10, 1.664877e-10, 1.670346e-10, 1.670222e-10, 
    1.676308e-10, 1.673564e-10, 1.68379e-10, 1.680884e-10, 1.68928e-10, 
    1.687169e-10, 1.68918e-10, 1.688571e-10, 1.689188e-10, 1.686092e-10, 
    1.687419e-10, 1.684694e-10, 1.674078e-10, 1.677198e-10, 1.66789e-10, 
    1.662289e-10, 1.65857e-10, 1.655929e-10, 1.656302e-10, 1.657014e-10, 
    1.66067e-10, 1.664108e-10, 1.666727e-10, 1.668479e-10, 1.670205e-10, 
    1.675426e-10, 1.67819e-10, 1.684377e-10, 1.683261e-10, 1.685152e-10, 
    1.686959e-10, 1.689991e-10, 1.689492e-10, 1.690828e-10, 1.685102e-10, 
    1.688907e-10, 1.682626e-10, 1.684344e-10, 1.670671e-10, 1.665463e-10, 
    1.663246e-10, 1.661308e-10, 1.656589e-10, 1.659848e-10, 1.658563e-10, 
    1.66162e-10, 1.663561e-10, 1.662601e-10, 1.668527e-10, 1.666223e-10, 
    1.678354e-10, 1.67313e-10, 1.686748e-10, 1.68349e-10, 1.687529e-10, 
    1.685468e-10, 1.688998e-10, 1.685821e-10, 1.691325e-10, 1.692523e-10, 
    1.691704e-10, 1.694849e-10, 1.685645e-10, 1.68918e-10, 1.662574e-10, 
    1.662731e-10, 1.66346e-10, 1.660253e-10, 1.660056e-10, 1.657117e-10, 
    1.659733e-10, 1.660846e-10, 1.663674e-10, 1.665346e-10, 1.666935e-10, 
    1.670429e-10, 1.67433e-10, 1.679784e-10, 1.683702e-10, 1.686327e-10, 
    1.684717e-10, 1.686138e-10, 1.68455e-10, 1.683805e-10, 1.692074e-10, 
    1.687431e-10, 1.694397e-10, 1.694012e-10, 1.690859e-10, 1.694055e-10, 
    1.662841e-10, 1.66194e-10, 1.65881e-10, 1.661259e-10, 1.656797e-10, 
    1.659295e-10, 1.66073e-10, 1.666271e-10, 1.667488e-10, 1.668617e-10, 
    1.670845e-10, 1.673705e-10, 1.67872e-10, 1.683082e-10, 1.687064e-10, 
    1.686772e-10, 1.686875e-10, 1.687764e-10, 1.685561e-10, 1.688126e-10, 
    1.688556e-10, 1.687431e-10, 1.69396e-10, 1.692095e-10, 1.694004e-10, 
    1.692789e-10, 1.662233e-10, 1.663749e-10, 1.66293e-10, 1.66447e-10, 
    1.663385e-10, 1.66821e-10, 1.669657e-10, 1.676425e-10, 1.673648e-10, 
    1.678068e-10, 1.674097e-10, 1.674801e-10, 1.678211e-10, 1.674312e-10, 
    1.682841e-10, 1.677058e-10, 1.687799e-10, 1.682025e-10, 1.68816e-10, 
    1.687047e-10, 1.688891e-10, 1.690542e-10, 1.692619e-10, 1.696451e-10, 
    1.695564e-10, 1.698768e-10, 1.666009e-10, 1.667975e-10, 1.667803e-10, 
    1.66986e-10, 1.671382e-10, 1.67468e-10, 1.679967e-10, 1.677979e-10, 
    1.681629e-10, 1.682361e-10, 1.676816e-10, 1.680221e-10, 1.669291e-10, 
    1.671057e-10, 1.670006e-10, 1.666164e-10, 1.678436e-10, 1.672139e-10, 
    1.683766e-10, 1.680356e-10, 1.690306e-10, 1.685358e-10, 1.695075e-10, 
    1.699226e-10, 1.703135e-10, 1.707698e-10, 1.669049e-10, 1.667713e-10, 
    1.670105e-10, 1.673413e-10, 1.676484e-10, 1.680564e-10, 1.680982e-10, 
    1.681746e-10, 1.683726e-10, 1.68539e-10, 1.681987e-10, 1.685807e-10, 
    1.671466e-10, 1.678983e-10, 1.667207e-10, 1.670754e-10, 1.673219e-10, 
    1.672138e-10, 1.677752e-10, 1.679075e-10, 1.684448e-10, 1.681671e-10, 
    1.698202e-10, 1.69089e-10, 1.711174e-10, 1.705507e-10, 1.667246e-10, 
    1.669044e-10, 1.675301e-10, 1.672325e-10, 1.680837e-10, 1.682931e-10, 
    1.684634e-10, 1.68681e-10, 1.687045e-10, 1.688334e-10, 1.686221e-10, 
    1.688251e-10, 1.680573e-10, 1.684004e-10, 1.674587e-10, 1.676879e-10, 
    1.675824e-10, 1.674668e-10, 1.678238e-10, 1.68204e-10, 1.682122e-10, 
    1.683341e-10, 1.686774e-10, 1.680871e-10, 1.699144e-10, 1.68786e-10, 
    1.671005e-10, 1.674467e-10, 1.674962e-10, 1.673621e-10, 1.682721e-10, 
    1.679424e-10, 1.688302e-10, 1.685904e-10, 1.689834e-10, 1.687881e-10, 
    1.687594e-10, 1.685085e-10, 1.683523e-10, 1.679575e-10, 1.676363e-10, 
    1.673816e-10, 1.674408e-10, 1.677206e-10, 1.682273e-10, 1.687066e-10, 
    1.686016e-10, 1.689535e-10, 1.68022e-10, 1.684126e-10, 1.682616e-10, 
    1.686553e-10, 1.677926e-10, 1.685271e-10, 1.676048e-10, 1.676857e-10, 
    1.679359e-10, 1.684391e-10, 1.685505e-10, 1.686693e-10, 1.68596e-10, 
    1.682402e-10, 1.681819e-10, 1.679298e-10, 1.678602e-10, 1.676681e-10, 
    1.67509e-10, 1.676543e-10, 1.678069e-10, 1.682404e-10, 1.686309e-10, 
    1.690565e-10, 1.691607e-10, 1.696577e-10, 1.69253e-10, 1.699206e-10, 
    1.693529e-10, 1.703356e-10, 1.685697e-10, 1.693364e-10, 1.679473e-10, 
    1.68097e-10, 1.683677e-10, 1.689885e-10, 1.686535e-10, 1.690454e-10, 
    1.681797e-10, 1.677302e-10, 1.67614e-10, 1.673971e-10, 1.67619e-10, 
    1.676009e-10, 1.678133e-10, 1.677451e-10, 1.682548e-10, 1.67981e-10, 
    1.687586e-10, 1.690423e-10, 1.698432e-10, 1.70334e-10, 1.708335e-10, 
    1.71054e-10, 1.711211e-10, 1.711491e-10 ;

 SOIL1N_vr =
  2.497551, 2.497545, 2.497546, 2.497541, 2.497544, 2.49754, 2.49755, 
    2.497545, 2.497548, 2.497551, 2.497531, 2.497541, 2.497521, 2.497527, 
    2.497512, 2.497522, 2.49751, 2.497512, 2.497505, 2.497507, 2.497498, 
    2.497504, 2.497494, 2.4975, 2.497499, 2.497505, 2.497539, 2.497532, 
    2.497539, 2.497538, 2.497539, 2.497544, 2.497546, 2.497552, 2.497551, 
    2.497547, 2.497538, 2.497541, 2.497533, 2.497534, 2.497525, 2.497529, 
    2.497515, 2.497519, 2.497507, 2.49751, 2.497507, 2.497508, 2.497507, 
    2.497512, 2.49751, 2.497514, 2.497528, 2.497524, 2.497537, 2.497545, 
    2.49755, 2.497553, 2.497553, 2.497552, 2.497547, 2.497542, 2.497538, 
    2.497536, 2.497534, 2.497526, 2.497523, 2.497514, 2.497516, 2.497513, 
    2.49751, 2.497506, 2.497507, 2.497505, 2.497513, 2.497508, 2.497516, 
    2.497514, 2.497533, 2.49754, 2.497543, 2.497546, 2.497552, 2.497548, 
    2.49755, 2.497545, 2.497543, 2.497544, 2.497536, 2.497539, 2.497522, 
    2.49753, 2.497511, 2.497515, 2.49751, 2.497513, 2.497508, 2.497512, 
    2.497504, 2.497503, 2.497504, 2.4975, 2.497512, 2.497507, 2.497544, 
    2.497544, 2.497543, 2.497547, 2.497548, 2.497552, 2.497548, 2.497546, 
    2.497543, 2.49754, 2.497538, 2.497533, 2.497528, 2.49752, 2.497515, 
    2.497511, 2.497514, 2.497512, 2.497514, 2.497515, 2.497504, 2.49751, 
    2.4975, 2.497501, 2.497505, 2.497501, 2.497544, 2.497545, 2.497549, 
    2.497546, 2.497552, 2.497549, 2.497547, 2.497539, 2.497537, 2.497536, 
    2.497533, 2.497529, 2.497522, 2.497516, 2.49751, 2.497511, 2.497511, 
    2.497509, 2.497512, 2.497509, 2.497508, 2.49751, 2.497501, 2.497503, 
    2.497501, 2.497502, 2.497545, 2.497543, 2.497544, 2.497541, 2.497543, 
    2.497536, 2.497534, 2.497525, 2.497529, 2.497523, 2.497528, 2.497527, 
    2.497523, 2.497528, 2.497516, 2.497524, 2.497509, 2.497517, 2.497509, 
    2.49751, 2.497508, 2.497505, 2.497503, 2.497497, 2.497499, 2.497494, 
    2.497539, 2.497537, 2.497537, 2.497534, 2.497532, 2.497527, 2.49752, 
    2.497523, 2.497518, 2.497517, 2.497524, 2.49752, 2.497535, 2.497532, 
    2.497534, 2.497539, 2.497522, 2.497531, 2.497515, 2.497519, 2.497506, 
    2.497513, 2.497499, 2.497494, 2.497488, 2.497482, 2.497535, 2.497537, 
    2.497534, 2.497529, 2.497525, 2.497519, 2.497519, 2.497518, 2.497515, 
    2.497513, 2.497517, 2.497512, 2.497532, 2.497521, 2.497538, 2.497533, 
    2.49753, 2.497531, 2.497523, 2.497521, 2.497514, 2.497518, 2.497495, 
    2.497505, 2.497477, 2.497485, 2.497538, 2.497535, 2.497527, 2.497531, 
    2.497519, 2.497516, 2.497514, 2.497511, 2.49751, 2.497509, 2.497511, 
    2.497509, 2.497519, 2.497514, 2.497528, 2.497524, 2.497526, 2.497527, 
    2.497523, 2.497517, 2.497517, 2.497515, 2.497511, 2.497519, 2.497494, 
    2.497509, 2.497532, 2.497528, 2.497527, 2.497529, 2.497516, 2.497521, 
    2.497509, 2.497512, 2.497507, 2.497509, 2.497509, 2.497513, 2.497515, 
    2.497521, 2.497525, 2.497529, 2.497528, 2.497524, 2.497517, 2.49751, 
    2.497512, 2.497507, 2.49752, 2.497514, 2.497516, 2.497511, 2.497523, 
    2.497513, 2.497525, 2.497524, 2.497521, 2.497514, 2.497513, 2.497511, 
    2.497512, 2.497517, 2.497518, 2.497521, 2.497522, 2.497525, 2.497527, 
    2.497525, 2.497523, 2.497517, 2.497511, 2.497505, 2.497504, 2.497497, 
    2.497503, 2.497494, 2.497501, 2.497488, 2.497512, 2.497502, 2.497521, 
    2.497519, 2.497515, 2.497506, 2.497511, 2.497506, 2.497518, 2.497524, 
    2.497525, 2.497528, 2.497525, 2.497525, 2.497523, 2.497524, 2.497517, 
    2.49752, 2.49751, 2.497506, 2.497495, 2.497488, 2.497481, 2.497478, 
    2.497477, 2.497477,
  2.497528, 2.497521, 2.497523, 2.497517, 2.49752, 2.497517, 2.497526, 
    2.497521, 2.497524, 2.497527, 2.497507, 2.497517, 2.497497, 2.497503, 
    2.497487, 2.497498, 2.497485, 2.497488, 2.49748, 2.497482, 2.497473, 
    2.497479, 2.497468, 2.497474, 2.497473, 2.497479, 2.497515, 2.497508, 
    2.497515, 2.497514, 2.497515, 2.49752, 2.497523, 2.497528, 2.497527, 
    2.497523, 2.497514, 2.497517, 2.497509, 2.497509, 2.497501, 2.497505, 
    2.49749, 2.497494, 2.497482, 2.497485, 2.497482, 2.497483, 2.497482, 
    2.497487, 2.497485, 2.497489, 2.497504, 2.497499, 2.497513, 2.497521, 
    2.497526, 2.49753, 2.49753, 2.497529, 2.497523, 2.497518, 2.497514, 
    2.497512, 2.497509, 2.497502, 2.497498, 2.497489, 2.497491, 2.497488, 
    2.497485, 2.497481, 2.497482, 2.49748, 2.497488, 2.497483, 2.497492, 
    2.497489, 2.497509, 2.497516, 2.497519, 2.497522, 2.497529, 2.497524, 
    2.497526, 2.497522, 2.497519, 2.49752, 2.497512, 2.497515, 2.497498, 
    2.497505, 2.497486, 2.49749, 2.497485, 2.497488, 2.497483, 2.497487, 
    2.497479, 2.497478, 2.497479, 2.497474, 2.497487, 2.497482, 2.49752, 
    2.49752, 2.497519, 2.497524, 2.497524, 2.497528, 2.497524, 2.497523, 
    2.497519, 2.497516, 2.497514, 2.497509, 2.497504, 2.497496, 2.49749, 
    2.497486, 2.497489, 2.497487, 2.497489, 2.49749, 2.497478, 2.497485, 
    2.497475, 2.497475, 2.49748, 2.497475, 2.49752, 2.497521, 2.497526, 
    2.497522, 2.497529, 2.497525, 2.497523, 2.497515, 2.497513, 2.497512, 
    2.497509, 2.497504, 2.497497, 2.497491, 2.497485, 2.497486, 2.497486, 
    2.497484, 2.497488, 2.497484, 2.497483, 2.497485, 2.497475, 2.497478, 
    2.497475, 2.497477, 2.497521, 2.497519, 2.49752, 2.497518, 2.497519, 
    2.497512, 2.49751, 2.497501, 2.497504, 2.497498, 2.497504, 2.497503, 
    2.497498, 2.497504, 2.497491, 2.4975, 2.497484, 2.497493, 2.497484, 
    2.497485, 2.497483, 2.49748, 2.497478, 2.497472, 2.497473, 2.497469, 
    2.497515, 2.497513, 2.497513, 2.49751, 2.497508, 2.497503, 2.497495, 
    2.497498, 2.497493, 2.497492, 2.4975, 2.497495, 2.497511, 2.497508, 
    2.49751, 2.497515, 2.497498, 2.497507, 2.49749, 2.497495, 2.497481, 
    2.497488, 2.497474, 2.497468, 2.497463, 2.497456, 2.497511, 2.497513, 
    2.49751, 2.497505, 2.4975, 2.497495, 2.497494, 2.497493, 2.49749, 
    2.497488, 2.497493, 2.497487, 2.497508, 2.497497, 2.497514, 2.497509, 
    2.497505, 2.497507, 2.497499, 2.497497, 2.497489, 2.497493, 2.497469, 
    2.49748, 2.497451, 2.497459, 2.497514, 2.497511, 2.497502, 2.497506, 
    2.497494, 2.497491, 2.497489, 2.497486, 2.497485, 2.497483, 2.497487, 
    2.497484, 2.497495, 2.49749, 2.497503, 2.4975, 2.497501, 2.497503, 
    2.497498, 2.497493, 2.497492, 2.497491, 2.497486, 2.497494, 2.497468, 
    2.497484, 2.497508, 2.497503, 2.497503, 2.497505, 2.497492, 2.497496, 
    2.497483, 2.497487, 2.497481, 2.497484, 2.497485, 2.497488, 2.49749, 
    2.497496, 2.497501, 2.497504, 2.497504, 2.497499, 2.497492, 2.497485, 
    2.497487, 2.497482, 2.497495, 2.497489, 2.497492, 2.497486, 2.497499, 
    2.497488, 2.497501, 2.4975, 2.497496, 2.497489, 2.497488, 2.497486, 
    2.497487, 2.497492, 2.497493, 2.497496, 2.497498, 2.4975, 2.497503, 
    2.4975, 2.497498, 2.497492, 2.497486, 2.49748, 2.497479, 2.497472, 
    2.497478, 2.497468, 2.497476, 2.497462, 2.497487, 2.497476, 2.497496, 
    2.497494, 2.49749, 2.497481, 2.497486, 2.497481, 2.497493, 2.497499, 
    2.497501, 2.497504, 2.497501, 2.497501, 2.497498, 2.497499, 2.497492, 
    2.497496, 2.497485, 2.497481, 2.497469, 2.497462, 2.497455, 2.497452, 
    2.497451, 2.497451,
  2.49752, 2.497513, 2.497514, 2.497509, 2.497512, 2.497509, 2.497518, 
    2.497513, 2.497516, 2.497519, 2.497499, 2.497509, 2.497488, 2.497495, 
    2.497478, 2.497489, 2.497476, 2.497479, 2.497471, 2.497473, 2.497464, 
    2.49747, 2.497459, 2.497466, 2.497464, 2.497471, 2.497507, 2.4975, 
    2.497507, 2.497506, 2.497507, 2.497512, 2.497514, 2.49752, 2.497519, 
    2.497515, 2.497506, 2.497509, 2.497501, 2.497501, 2.497492, 2.497496, 
    2.497481, 2.497486, 2.497473, 2.497476, 2.497473, 2.497474, 2.497473, 
    2.497478, 2.497476, 2.49748, 2.497495, 2.497491, 2.497504, 2.497513, 
    2.497518, 2.497522, 2.497521, 2.49752, 2.497515, 2.49751, 2.497506, 
    2.497504, 2.497501, 2.497494, 2.497489, 2.49748, 2.497482, 2.497479, 
    2.497477, 2.497472, 2.497473, 2.497471, 2.497479, 2.497474, 2.497483, 
    2.497481, 2.4975, 2.497508, 2.497511, 2.497514, 2.497521, 2.497516, 
    2.497518, 2.497514, 2.497511, 2.497512, 2.497504, 2.497507, 2.497489, 
    2.497497, 2.497477, 2.497482, 2.497476, 2.497479, 2.497474, 2.497478, 
    2.49747, 2.497469, 2.49747, 2.497465, 2.497479, 2.497473, 2.497512, 
    2.497512, 2.497511, 2.497516, 2.497516, 2.49752, 2.497516, 2.497515, 
    2.497511, 2.497508, 2.497506, 2.497501, 2.497495, 2.497487, 2.497482, 
    2.497478, 2.49748, 2.497478, 2.49748, 2.497481, 2.497469, 2.497476, 
    2.497466, 2.497467, 2.497471, 2.497467, 2.497512, 2.497513, 2.497518, 
    2.497514, 2.497521, 2.497517, 2.497515, 2.497507, 2.497505, 2.497504, 
    2.4975, 2.497496, 2.497489, 2.497482, 2.497477, 2.497477, 2.497477, 
    2.497476, 2.497479, 2.497475, 2.497474, 2.497476, 2.497467, 2.497469, 
    2.497467, 2.497468, 2.497513, 2.49751, 2.497512, 2.497509, 2.497511, 
    2.497504, 2.497502, 2.497492, 2.497496, 2.49749, 2.497495, 2.497494, 
    2.497489, 2.497495, 2.497483, 2.497491, 2.497476, 2.497484, 2.497475, 
    2.497477, 2.497474, 2.497472, 2.497468, 2.497463, 2.497464, 2.49746, 
    2.497507, 2.497504, 2.497505, 2.497502, 2.497499, 2.497495, 2.497487, 
    2.49749, 2.497484, 2.497483, 2.497492, 2.497487, 2.497502, 2.4975, 
    2.497501, 2.497507, 2.497489, 2.497498, 2.497481, 2.497486, 2.497472, 
    2.497479, 2.497465, 2.497459, 2.497453, 2.497447, 2.497503, 2.497505, 
    2.497501, 2.497496, 2.497492, 2.497486, 2.497485, 2.497484, 2.497481, 
    2.497479, 2.497484, 2.497478, 2.497499, 2.497488, 2.497505, 2.4975, 
    2.497497, 2.497498, 2.49749, 2.497488, 2.49748, 2.497484, 2.49746, 
    2.497471, 2.497442, 2.49745, 2.497505, 2.497503, 2.497494, 2.497498, 
    2.497486, 2.497483, 2.49748, 2.497477, 2.497477, 2.497475, 2.497478, 
    2.497475, 2.497486, 2.497481, 2.497495, 2.497491, 2.497493, 2.497495, 
    2.497489, 2.497484, 2.497484, 2.497482, 2.497477, 2.497486, 2.497459, 
    2.497475, 2.4975, 2.497495, 2.497494, 2.497496, 2.497483, 2.497488, 
    2.497475, 2.497478, 2.497473, 2.497475, 2.497476, 2.497479, 2.497482, 
    2.497488, 2.497492, 2.497496, 2.497495, 2.497491, 2.497483, 2.497477, 
    2.497478, 2.497473, 2.497487, 2.497481, 2.497483, 2.497477, 2.49749, 
    2.497479, 2.497493, 2.497491, 2.497488, 2.49748, 2.497479, 2.497477, 
    2.497478, 2.497483, 2.497484, 2.497488, 2.497489, 2.497492, 2.497494, 
    2.497492, 2.49749, 2.497483, 2.497478, 2.497472, 2.49747, 2.497463, 
    2.497469, 2.497459, 2.497467, 2.497453, 2.497478, 2.497468, 2.497488, 
    2.497485, 2.497482, 2.497473, 2.497477, 2.497472, 2.497484, 2.497491, 
    2.497493, 2.497496, 2.497492, 2.497493, 2.49749, 2.497491, 2.497483, 
    2.497487, 2.497476, 2.497472, 2.49746, 2.497453, 2.497446, 2.497442, 
    2.497442, 2.497441,
  2.497595, 2.497589, 2.49759, 2.497585, 2.497588, 2.497584, 2.497594, 
    2.497589, 2.497592, 2.497595, 2.497575, 2.497585, 2.497564, 2.497571, 
    2.497555, 2.497565, 2.497553, 2.497555, 2.497548, 2.49755, 2.49754, 
    2.497547, 2.497535, 2.497542, 2.497541, 2.497547, 2.497583, 2.497576, 
    2.497583, 2.497582, 2.497582, 2.497588, 2.49759, 2.497596, 2.497595, 
    2.497591, 2.497582, 2.497585, 2.497577, 2.497577, 2.497568, 2.497572, 
    2.497558, 2.497562, 2.49755, 2.497553, 2.49755, 2.497551, 2.49755, 
    2.497554, 2.497552, 2.497556, 2.497571, 2.497567, 2.497581, 2.497588, 
    2.497594, 2.497598, 2.497597, 2.497596, 2.497591, 2.497586, 2.497582, 
    2.49758, 2.497577, 2.49757, 2.497566, 2.497557, 2.497558, 2.497556, 
    2.497553, 2.497549, 2.497549, 2.497547, 2.497556, 2.49755, 2.497559, 
    2.497557, 2.497576, 2.497584, 2.497587, 2.49759, 2.497597, 2.497592, 
    2.497594, 2.497589, 2.497587, 2.497588, 2.49758, 2.497583, 2.497566, 
    2.497573, 2.497553, 2.497558, 2.497552, 2.497555, 2.49755, 2.497555, 
    2.497547, 2.497545, 2.497546, 2.497542, 2.497555, 2.49755, 2.497588, 
    2.497588, 2.497587, 2.497591, 2.497592, 2.497596, 2.497592, 2.497591, 
    2.497586, 2.497584, 2.497582, 2.497577, 2.497571, 2.497563, 2.497558, 
    2.497554, 2.497556, 2.497554, 2.497556, 2.497558, 2.497546, 2.497552, 
    2.497542, 2.497543, 2.497547, 2.497543, 2.497588, 2.497589, 2.497593, 
    2.49759, 2.497597, 2.497593, 2.497591, 2.497583, 2.497581, 2.497579, 
    2.497576, 2.497572, 2.497565, 2.497559, 2.497553, 2.497553, 2.497553, 
    2.497552, 2.497555, 2.497551, 2.497551, 2.497552, 2.497543, 2.497546, 
    2.497543, 2.497545, 2.497589, 2.497586, 2.497588, 2.497585, 2.497587, 
    2.49758, 2.497578, 2.497568, 2.497572, 2.497566, 2.497571, 2.497571, 
    2.497566, 2.497571, 2.497559, 2.497567, 2.497552, 2.49756, 2.497551, 
    2.497553, 2.49755, 2.497548, 2.497545, 2.49754, 2.497541, 2.497536, 
    2.497583, 2.49758, 2.497581, 2.497578, 2.497576, 2.497571, 2.497563, 
    2.497566, 2.497561, 2.49756, 2.497568, 2.497563, 2.497578, 2.497576, 
    2.497577, 2.497583, 2.497565, 2.497574, 2.497558, 2.497562, 2.497548, 
    2.497555, 2.497541, 2.497535, 2.49753, 2.497523, 2.497579, 2.497581, 
    2.497577, 2.497572, 2.497568, 2.497562, 2.497562, 2.497561, 2.497558, 
    2.497555, 2.49756, 2.497555, 2.497575, 2.497565, 2.497581, 2.497576, 
    2.497573, 2.497574, 2.497566, 2.497564, 2.497557, 2.497561, 2.497537, 
    2.497547, 2.497518, 2.497526, 2.497581, 2.497579, 2.49757, 2.497574, 
    2.497562, 2.497559, 2.497556, 2.497553, 2.497553, 2.497551, 2.497554, 
    2.497551, 2.497562, 2.497557, 2.497571, 2.497567, 2.497569, 2.497571, 
    2.497566, 2.49756, 2.49756, 2.497558, 2.497553, 2.497562, 2.497535, 
    2.497552, 2.497576, 2.497571, 2.49757, 2.497572, 2.497559, 2.497564, 
    2.497551, 2.497555, 2.497549, 2.497552, 2.497552, 2.497556, 2.497558, 
    2.497564, 2.497568, 2.497572, 2.497571, 2.497567, 2.49756, 2.497553, 
    2.497554, 2.497549, 2.497563, 2.497557, 2.497559, 2.497554, 2.497566, 
    2.497555, 2.497569, 2.497568, 2.497564, 2.497557, 2.497555, 2.497553, 
    2.497555, 2.49756, 2.497561, 2.497564, 2.497565, 2.497568, 2.49757, 
    2.497568, 2.497566, 2.49756, 2.497554, 2.497548, 2.497546, 2.497539, 
    2.497545, 2.497535, 2.497544, 2.49753, 2.497555, 2.497544, 2.497564, 
    2.497562, 2.497558, 2.497549, 2.497554, 2.497548, 2.497561, 2.497567, 
    2.497569, 2.497572, 2.497569, 2.497569, 2.497566, 2.497567, 2.497559, 
    2.497563, 2.497552, 2.497548, 2.497537, 2.49753, 2.497522, 2.497519, 
    2.497518, 2.497518,
  2.497849, 2.497843, 2.497844, 2.497839, 2.497842, 2.497839, 2.497848, 
    2.497843, 2.497846, 2.497849, 2.49783, 2.497839, 2.49782, 2.497826, 
    2.497811, 2.497821, 2.497809, 2.497812, 2.497805, 2.497807, 2.497798, 
    2.497804, 2.497793, 2.497799, 2.497798, 2.497804, 2.497837, 2.497831, 
    2.497838, 2.497837, 2.497837, 2.497842, 2.497844, 2.497849, 2.497849, 
    2.497845, 2.497836, 2.497839, 2.497832, 2.497832, 2.497824, 2.497828, 
    2.497814, 2.497818, 2.497807, 2.497809, 2.497807, 2.497808, 2.497807, 
    2.497811, 2.497809, 2.497813, 2.497827, 2.497823, 2.497835, 2.497843, 
    2.497848, 2.497851, 2.497851, 2.49785, 2.497845, 2.49784, 2.497837, 
    2.497834, 2.497832, 2.497825, 2.497822, 2.497813, 2.497815, 2.497812, 
    2.49781, 2.497806, 2.497806, 2.497805, 2.497812, 2.497807, 2.497816, 
    2.497813, 2.497832, 2.497838, 2.497841, 2.497844, 2.49785, 2.497846, 
    2.497848, 2.497844, 2.497841, 2.497842, 2.497834, 2.497838, 2.497821, 
    2.497828, 2.49781, 2.497814, 2.497809, 2.497812, 2.497807, 2.497811, 
    2.497804, 2.497802, 2.497803, 2.497799, 2.497812, 2.497807, 2.497842, 
    2.497842, 2.497841, 2.497845, 2.497846, 2.49785, 2.497846, 2.497845, 
    2.497841, 2.497839, 2.497837, 2.497832, 2.497827, 2.497819, 2.497814, 
    2.497811, 2.497813, 2.497811, 2.497813, 2.497814, 2.497803, 2.497809, 
    2.4978, 2.4978, 2.497804, 2.4978, 2.497842, 2.497843, 2.497847, 2.497844, 
    2.49785, 2.497847, 2.497845, 2.497837, 2.497836, 2.497834, 2.497831, 
    2.497828, 2.497821, 2.497815, 2.49781, 2.49781, 2.49781, 2.497809, 
    2.497812, 2.497808, 2.497808, 2.497809, 2.4978, 2.497803, 2.4978, 
    2.497802, 2.497843, 2.497841, 2.497842, 2.49784, 2.497841, 2.497835, 
    2.497833, 2.497824, 2.497828, 2.497822, 2.497827, 2.497826, 2.497821, 
    2.497827, 2.497815, 2.497823, 2.497809, 2.497816, 2.497808, 2.49781, 
    2.497807, 2.497805, 2.497802, 2.497797, 2.497798, 2.497794, 2.497838, 
    2.497835, 2.497835, 2.497833, 2.497831, 2.497826, 2.497819, 2.497822, 
    2.497817, 2.497816, 2.497823, 2.497819, 2.497833, 2.497831, 2.497832, 
    2.497838, 2.497821, 2.497829, 2.497814, 2.497818, 2.497805, 2.497812, 
    2.497799, 2.497793, 2.497788, 2.497782, 2.497834, 2.497835, 2.497832, 
    2.497828, 2.497824, 2.497818, 2.497818, 2.497817, 2.497814, 2.497812, 
    2.497816, 2.497811, 2.49783, 2.49782, 2.497836, 2.497831, 2.497828, 
    2.497829, 2.497822, 2.49782, 2.497813, 2.497817, 2.497795, 2.497804, 
    2.497777, 2.497785, 2.497836, 2.497834, 2.497825, 2.497829, 2.497818, 
    2.497815, 2.497813, 2.49781, 2.49781, 2.497808, 2.497811, 2.497808, 
    2.497818, 2.497814, 2.497826, 2.497823, 2.497825, 2.497826, 2.497821, 
    2.497816, 2.497816, 2.497815, 2.49781, 2.497818, 2.497793, 2.497808, 
    2.497831, 2.497826, 2.497826, 2.497828, 2.497815, 2.49782, 2.497808, 
    2.497811, 2.497806, 2.497808, 2.497809, 2.497812, 2.497814, 2.49782, 
    2.497824, 2.497827, 2.497827, 2.497823, 2.497816, 2.49781, 2.497811, 
    2.497806, 2.497819, 2.497813, 2.497816, 2.49781, 2.497822, 2.497812, 
    2.497824, 2.497823, 2.49782, 2.497813, 2.497812, 2.49781, 2.497811, 
    2.497816, 2.497817, 2.49782, 2.497821, 2.497823, 2.497826, 2.497824, 
    2.497822, 2.497816, 2.497811, 2.497805, 2.497803, 2.497797, 2.497802, 
    2.497793, 2.497801, 2.497788, 2.497811, 2.497801, 2.49782, 2.497818, 
    2.497814, 2.497806, 2.49781, 2.497805, 2.497817, 2.497823, 2.497824, 
    2.497827, 2.497824, 2.497824, 2.497822, 2.497823, 2.497816, 2.497819, 
    2.497809, 2.497805, 2.497794, 2.497788, 2.497781, 2.497778, 2.497777, 
    2.497777,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1_HR_S2 =
  7.36236e-08, 7.382512e-08, 7.378596e-08, 7.394845e-08, 7.385833e-08, 
    7.396471e-08, 7.366447e-08, 7.383311e-08, 7.372547e-08, 7.364176e-08, 
    7.426365e-08, 7.395571e-08, 7.458355e-08, 7.438722e-08, 7.488035e-08, 
    7.455299e-08, 7.494635e-08, 7.487094e-08, 7.509796e-08, 7.503293e-08, 
    7.532315e-08, 7.512797e-08, 7.547361e-08, 7.527657e-08, 7.530738e-08, 
    7.512153e-08, 7.401772e-08, 7.422531e-08, 7.400541e-08, 7.403502e-08, 
    7.402173e-08, 7.386018e-08, 7.377873e-08, 7.360821e-08, 7.363918e-08, 
    7.376443e-08, 7.404833e-08, 7.395199e-08, 7.419483e-08, 7.418935e-08, 
    7.445959e-08, 7.433776e-08, 7.479186e-08, 7.466283e-08, 7.503564e-08, 
    7.49419e-08, 7.503124e-08, 7.500415e-08, 7.503159e-08, 7.48941e-08, 
    7.495301e-08, 7.483202e-08, 7.436057e-08, 7.449915e-08, 7.408575e-08, 
    7.383704e-08, 7.367186e-08, 7.355461e-08, 7.357119e-08, 7.360278e-08, 
    7.376516e-08, 7.391782e-08, 7.403413e-08, 7.411192e-08, 7.418856e-08, 
    7.442042e-08, 7.454319e-08, 7.481793e-08, 7.476838e-08, 7.485234e-08, 
    7.493257e-08, 7.506723e-08, 7.504507e-08, 7.510438e-08, 7.485014e-08, 
    7.501911e-08, 7.474015e-08, 7.481646e-08, 7.420929e-08, 7.397799e-08, 
    7.387956e-08, 7.379348e-08, 7.358393e-08, 7.372864e-08, 7.36716e-08, 
    7.380733e-08, 7.389355e-08, 7.385091e-08, 7.411405e-08, 7.401175e-08, 
    7.455046e-08, 7.431847e-08, 7.492321e-08, 7.477855e-08, 7.495789e-08, 
    7.486639e-08, 7.502315e-08, 7.488207e-08, 7.512647e-08, 7.517966e-08, 
    7.51433e-08, 7.528298e-08, 7.487424e-08, 7.503122e-08, 7.384971e-08, 
    7.385666e-08, 7.388906e-08, 7.374661e-08, 7.37379e-08, 7.360736e-08, 
    7.372353e-08, 7.377298e-08, 7.389855e-08, 7.397279e-08, 7.404338e-08, 
    7.419853e-08, 7.437176e-08, 7.461396e-08, 7.478793e-08, 7.490451e-08, 
    7.483304e-08, 7.489614e-08, 7.482559e-08, 7.479253e-08, 7.515972e-08, 
    7.495355e-08, 7.526289e-08, 7.524578e-08, 7.510579e-08, 7.52477e-08, 
    7.386154e-08, 7.382153e-08, 7.368254e-08, 7.379131e-08, 7.359314e-08, 
    7.370407e-08, 7.376783e-08, 7.401387e-08, 7.406794e-08, 7.411804e-08, 
    7.421701e-08, 7.434399e-08, 7.456669e-08, 7.476042e-08, 7.493725e-08, 
    7.492429e-08, 7.492885e-08, 7.496833e-08, 7.487051e-08, 7.498439e-08, 
    7.50035e-08, 7.495354e-08, 7.524348e-08, 7.516066e-08, 7.524542e-08, 
    7.519149e-08, 7.383454e-08, 7.390187e-08, 7.386549e-08, 7.39339e-08, 
    7.38857e-08, 7.41e-08, 7.416425e-08, 7.446479e-08, 7.434149e-08, 
    7.453775e-08, 7.436144e-08, 7.439268e-08, 7.454411e-08, 7.437097e-08, 
    7.474972e-08, 7.449292e-08, 7.496987e-08, 7.471347e-08, 7.498593e-08, 
    7.493648e-08, 7.501837e-08, 7.509169e-08, 7.518394e-08, 7.535409e-08, 
    7.53147e-08, 7.5457e-08, 7.400226e-08, 7.408956e-08, 7.40819e-08, 
    7.417327e-08, 7.424084e-08, 7.438729e-08, 7.462208e-08, 7.45338e-08, 
    7.469588e-08, 7.47284e-08, 7.448218e-08, 7.463335e-08, 7.414801e-08, 
    7.422642e-08, 7.417975e-08, 7.400914e-08, 7.455412e-08, 7.427447e-08, 
    7.47908e-08, 7.463937e-08, 7.508123e-08, 7.48615e-08, 7.529301e-08, 
    7.547735e-08, 7.56509e-08, 7.585354e-08, 7.413723e-08, 7.407792e-08, 
    7.418414e-08, 7.433106e-08, 7.446741e-08, 7.46486e-08, 7.466715e-08, 
    7.470108e-08, 7.4789e-08, 7.48629e-08, 7.471179e-08, 7.488142e-08, 
    7.424457e-08, 7.45784e-08, 7.405547e-08, 7.421294e-08, 7.432241e-08, 
    7.427441e-08, 7.452372e-08, 7.458246e-08, 7.48211e-08, 7.469776e-08, 
    7.543184e-08, 7.510715e-08, 7.600787e-08, 7.575625e-08, 7.405718e-08, 
    7.413704e-08, 7.441488e-08, 7.42827e-08, 7.46607e-08, 7.475371e-08, 
    7.482933e-08, 7.492595e-08, 7.493639e-08, 7.499364e-08, 7.489983e-08, 
    7.498994e-08, 7.464899e-08, 7.480137e-08, 7.438316e-08, 7.448496e-08, 
    7.443813e-08, 7.438675e-08, 7.454531e-08, 7.471417e-08, 7.471781e-08, 
    7.477194e-08, 7.492439e-08, 7.466225e-08, 7.547367e-08, 7.49726e-08, 
    7.422411e-08, 7.437784e-08, 7.439984e-08, 7.434029e-08, 7.474439e-08, 
    7.459799e-08, 7.499224e-08, 7.488572e-08, 7.506026e-08, 7.497353e-08, 
    7.496077e-08, 7.484937e-08, 7.477999e-08, 7.46047e-08, 7.446205e-08, 
    7.434893e-08, 7.437524e-08, 7.449949e-08, 7.47245e-08, 7.493733e-08, 
    7.489071e-08, 7.5047e-08, 7.463331e-08, 7.480678e-08, 7.473973e-08, 
    7.491457e-08, 7.453146e-08, 7.485761e-08, 7.444805e-08, 7.448397e-08, 
    7.459509e-08, 7.481853e-08, 7.486801e-08, 7.492076e-08, 7.488821e-08, 
    7.473022e-08, 7.470435e-08, 7.459239e-08, 7.456146e-08, 7.447616e-08, 
    7.44055e-08, 7.447004e-08, 7.453782e-08, 7.473029e-08, 7.490371e-08, 
    7.509272e-08, 7.513899e-08, 7.535969e-08, 7.518e-08, 7.547646e-08, 
    7.522436e-08, 7.566075e-08, 7.487656e-08, 7.5217e-08, 7.460015e-08, 
    7.466664e-08, 7.478685e-08, 7.506254e-08, 7.491375e-08, 7.508777e-08, 
    7.470334e-08, 7.450377e-08, 7.445216e-08, 7.43558e-08, 7.445436e-08, 
    7.444635e-08, 7.454064e-08, 7.451035e-08, 7.473669e-08, 7.461512e-08, 
    7.496044e-08, 7.50864e-08, 7.544207e-08, 7.566e-08, 7.588183e-08, 
    7.597973e-08, 7.600952e-08, 7.602198e-08 ;

 SOIL1_HR_S3 =
  8.73601e-10, 8.759933e-10, 8.755285e-10, 8.774574e-10, 8.763876e-10, 
    8.776506e-10, 8.740862e-10, 8.760881e-10, 8.748103e-10, 8.738166e-10, 
    8.811994e-10, 8.775436e-10, 8.849971e-10, 8.826664e-10, 8.885207e-10, 
    8.846343e-10, 8.893043e-10, 8.884091e-10, 8.911042e-10, 8.903322e-10, 
    8.937778e-10, 8.914605e-10, 8.95564e-10, 8.932247e-10, 8.935905e-10, 
    8.91384e-10, 8.782798e-10, 8.807443e-10, 8.781337e-10, 8.784852e-10, 
    8.783275e-10, 8.764096e-10, 8.754426e-10, 8.734184e-10, 8.73786e-10, 
    8.752729e-10, 8.786432e-10, 8.774995e-10, 8.803824e-10, 8.803173e-10, 
    8.835256e-10, 8.820792e-10, 8.874701e-10, 8.859383e-10, 8.903644e-10, 
    8.892515e-10, 8.903121e-10, 8.899905e-10, 8.903163e-10, 8.88684e-10, 
    8.893833e-10, 8.87947e-10, 8.8235e-10, 8.839951e-10, 8.790875e-10, 
    8.761348e-10, 8.74174e-10, 8.727821e-10, 8.729789e-10, 8.733539e-10, 
    8.752816e-10, 8.770938e-10, 8.784746e-10, 8.793981e-10, 8.80308e-10, 
    8.830606e-10, 8.84518e-10, 8.877796e-10, 8.871914e-10, 8.881881e-10, 
    8.891408e-10, 8.907393e-10, 8.904763e-10, 8.911805e-10, 8.881621e-10, 
    8.901681e-10, 8.868563e-10, 8.877621e-10, 8.80554e-10, 8.778082e-10, 
    8.766397e-10, 8.756178e-10, 8.731302e-10, 8.74848e-10, 8.741708e-10, 
    8.757821e-10, 8.768056e-10, 8.762995e-10, 8.794234e-10, 8.78209e-10, 
    8.846043e-10, 8.818501e-10, 8.890296e-10, 8.873122e-10, 8.894412e-10, 
    8.88355e-10, 8.902161e-10, 8.885411e-10, 8.914426e-10, 8.920742e-10, 
    8.916426e-10, 8.933008e-10, 8.884483e-10, 8.903119e-10, 8.762853e-10, 
    8.763678e-10, 8.767524e-10, 8.750614e-10, 8.749579e-10, 8.734083e-10, 
    8.747873e-10, 8.753744e-10, 8.768651e-10, 8.777465e-10, 8.785844e-10, 
    8.804263e-10, 8.824829e-10, 8.853581e-10, 8.874235e-10, 8.888076e-10, 
    8.87959e-10, 8.887082e-10, 8.878707e-10, 8.874781e-10, 8.918374e-10, 
    8.893898e-10, 8.930623e-10, 8.928592e-10, 8.911972e-10, 8.92882e-10, 
    8.764258e-10, 8.759508e-10, 8.743008e-10, 8.75592e-10, 8.732395e-10, 
    8.745563e-10, 8.753132e-10, 8.78234e-10, 8.78876e-10, 8.794708e-10, 
    8.806457e-10, 8.821532e-10, 8.847971e-10, 8.870969e-10, 8.891962e-10, 
    8.890424e-10, 8.890966e-10, 8.895653e-10, 8.88404e-10, 8.89756e-10, 
    8.899828e-10, 8.893896e-10, 8.92832e-10, 8.918487e-10, 8.928548e-10, 
    8.922147e-10, 8.761052e-10, 8.769045e-10, 8.764726e-10, 8.772848e-10, 
    8.767125e-10, 8.792566e-10, 8.800193e-10, 8.835873e-10, 8.821234e-10, 
    8.844535e-10, 8.823602e-10, 8.827312e-10, 8.84529e-10, 8.824735e-10, 
    8.869699e-10, 8.839213e-10, 8.895835e-10, 8.865395e-10, 8.897743e-10, 
    8.891871e-10, 8.901593e-10, 8.910297e-10, 8.92125e-10, 8.941451e-10, 
    8.936775e-10, 8.953668e-10, 8.780963e-10, 8.791327e-10, 8.790417e-10, 
    8.801264e-10, 8.809286e-10, 8.826671e-10, 8.854545e-10, 8.844065e-10, 
    8.863307e-10, 8.867169e-10, 8.837937e-10, 8.855884e-10, 8.798265e-10, 
    8.807574e-10, 8.802034e-10, 8.781779e-10, 8.846477e-10, 8.813278e-10, 
    8.874576e-10, 8.856598e-10, 8.909056e-10, 8.882969e-10, 8.934199e-10, 
    8.956085e-10, 8.976689e-10, 9.000749e-10, 8.796986e-10, 8.789944e-10, 
    8.802555e-10, 8.819996e-10, 8.836183e-10, 8.857694e-10, 8.859897e-10, 
    8.863925e-10, 8.874362e-10, 8.883135e-10, 8.865197e-10, 8.885335e-10, 
    8.809729e-10, 8.84936e-10, 8.787279e-10, 8.805974e-10, 8.818969e-10, 
    8.813271e-10, 8.842868e-10, 8.849841e-10, 8.878173e-10, 8.86353e-10, 
    8.950681e-10, 8.912133e-10, 9.019072e-10, 8.989198e-10, 8.787482e-10, 
    8.796963e-10, 8.829948e-10, 8.814255e-10, 8.859132e-10, 8.870173e-10, 
    8.879151e-10, 8.890621e-10, 8.891861e-10, 8.898657e-10, 8.88752e-10, 
    8.898218e-10, 8.857741e-10, 8.875831e-10, 8.826181e-10, 8.838267e-10, 
    8.832708e-10, 8.826608e-10, 8.845432e-10, 8.865478e-10, 8.86591e-10, 
    8.872337e-10, 8.890436e-10, 8.859314e-10, 8.955648e-10, 8.89616e-10, 
    8.8073e-10, 8.825551e-10, 8.828162e-10, 8.821092e-10, 8.869066e-10, 
    8.851686e-10, 8.898492e-10, 8.885845e-10, 8.906567e-10, 8.89627e-10, 
    8.894755e-10, 8.881529e-10, 8.873293e-10, 8.852482e-10, 8.835547e-10, 
    8.822118e-10, 8.825241e-10, 8.839992e-10, 8.866706e-10, 8.891972e-10, 
    8.886437e-10, 8.904992e-10, 8.855879e-10, 8.876474e-10, 8.868513e-10, 
    8.88927e-10, 8.843787e-10, 8.882508e-10, 8.833885e-10, 8.83815e-10, 
    8.851341e-10, 8.877868e-10, 8.883742e-10, 8.890005e-10, 8.886141e-10, 
    8.867384e-10, 8.864312e-10, 8.851021e-10, 8.847349e-10, 8.837222e-10, 
    8.828834e-10, 8.836497e-10, 8.844542e-10, 8.867393e-10, 8.88798e-10, 
    8.910421e-10, 8.915914e-10, 8.942115e-10, 8.920782e-10, 8.955979e-10, 
    8.926048e-10, 8.977859e-10, 8.884757e-10, 8.925174e-10, 8.851943e-10, 
    8.859836e-10, 8.874107e-10, 8.906837e-10, 8.889173e-10, 8.909833e-10, 
    8.864192e-10, 8.840499e-10, 8.834373e-10, 8.822933e-10, 8.834634e-10, 
    8.833683e-10, 8.844878e-10, 8.84128e-10, 8.868152e-10, 8.853719e-10, 
    8.894716e-10, 8.909671e-10, 8.951897e-10, 8.97777e-10, 9.004107e-10, 
    9.01573e-10, 9.019268e-10, 9.020746e-10 ;

 SOIL2C =
  5.784273, 5.784277, 5.784276, 5.78428, 5.784278, 5.784281, 5.784274, 
    5.784278, 5.784276, 5.784274, 5.784287, 5.784281, 5.784295, 5.78429, 
    5.784302, 5.784294, 5.784303, 5.784301, 5.784307, 5.784305, 5.784312, 
    5.784307, 5.784315, 5.784311, 5.784311, 5.784307, 5.784282, 5.784286, 
    5.784282, 5.784282, 5.784282, 5.784278, 5.784276, 5.784273, 5.784273, 
    5.784276, 5.784283, 5.78428, 5.784286, 5.784286, 5.784292, 5.784289, 
    5.784299, 5.784297, 5.784305, 5.784303, 5.784305, 5.784305, 5.784305, 
    5.784302, 5.784303, 5.7843, 5.78429, 5.784293, 5.784284, 5.784278, 
    5.784274, 5.784271, 5.784272, 5.784273, 5.784276, 5.78428, 5.784282, 
    5.784284, 5.784286, 5.784291, 5.784294, 5.7843, 5.784299, 5.784301, 
    5.784303, 5.784306, 5.784306, 5.784307, 5.784301, 5.784305, 5.784298, 
    5.7843, 5.784286, 5.784281, 5.784279, 5.784277, 5.784272, 5.784276, 
    5.784274, 5.784277, 5.784279, 5.784278, 5.784284, 5.784282, 5.784294, 
    5.784289, 5.784303, 5.784299, 5.784303, 5.784301, 5.784305, 5.784302, 
    5.784307, 5.784308, 5.784307, 5.784311, 5.784301, 5.784305, 5.784278, 
    5.784278, 5.784279, 5.784276, 5.784276, 5.784273, 5.784275, 5.784276, 
    5.784279, 5.784281, 5.784283, 5.784286, 5.78429, 5.784296, 5.784299, 
    5.784302, 5.7843, 5.784302, 5.7843, 5.784299, 5.784308, 5.784303, 
    5.78431, 5.78431, 5.784307, 5.78431, 5.784278, 5.784277, 5.784275, 
    5.784277, 5.784272, 5.784275, 5.784276, 5.784282, 5.784283, 5.784284, 
    5.784286, 5.784289, 5.784295, 5.784299, 5.784303, 5.784303, 5.784303, 
    5.784304, 5.784301, 5.784304, 5.784305, 5.784303, 5.78431, 5.784308, 
    5.78431, 5.784308, 5.784278, 5.784279, 5.784278, 5.78428, 5.784279, 
    5.784284, 5.784286, 5.784292, 5.784289, 5.784294, 5.78429, 5.78429, 
    5.784294, 5.78429, 5.784298, 5.784293, 5.784304, 5.784298, 5.784304, 
    5.784303, 5.784305, 5.784307, 5.784308, 5.784312, 5.784311, 5.784315, 
    5.784282, 5.784284, 5.784284, 5.784286, 5.784287, 5.78429, 5.784296, 
    5.784294, 5.784297, 5.784298, 5.784293, 5.784296, 5.784285, 5.784286, 
    5.784286, 5.784282, 5.784294, 5.784288, 5.784299, 5.784296, 5.784306, 
    5.784301, 5.784311, 5.784315, 5.784319, 5.784324, 5.784285, 5.784283, 
    5.784286, 5.784289, 5.784292, 5.784297, 5.784297, 5.784297, 5.784299, 
    5.784301, 5.784298, 5.784302, 5.784287, 5.784295, 5.784283, 5.784286, 
    5.784289, 5.784288, 5.784294, 5.784295, 5.7843, 5.784297, 5.784314, 
    5.784307, 5.784327, 5.784321, 5.784283, 5.784285, 5.784291, 5.784288, 
    5.784297, 5.784299, 5.7843, 5.784303, 5.784303, 5.784304, 5.784302, 
    5.784304, 5.784297, 5.7843, 5.78429, 5.784293, 5.784292, 5.78429, 
    5.784294, 5.784298, 5.784298, 5.784299, 5.784303, 5.784297, 5.784315, 
    5.784304, 5.784286, 5.78429, 5.784291, 5.784289, 5.784298, 5.784295, 
    5.784304, 5.784302, 5.784306, 5.784304, 5.784303, 5.784301, 5.784299, 
    5.784296, 5.784292, 5.784289, 5.78429, 5.784293, 5.784298, 5.784303, 
    5.784302, 5.784306, 5.784296, 5.7843, 5.784298, 5.784302, 5.784294, 
    5.784301, 5.784292, 5.784293, 5.784295, 5.7843, 5.784301, 5.784303, 
    5.784302, 5.784298, 5.784297, 5.784295, 5.784294, 5.784292, 5.784291, 
    5.784292, 5.784294, 5.784298, 5.784302, 5.784307, 5.784307, 5.784313, 
    5.784308, 5.784315, 5.784309, 5.784319, 5.784301, 5.784309, 5.784295, 
    5.784297, 5.784299, 5.784306, 5.784302, 5.784307, 5.784297, 5.784293, 
    5.784292, 5.78429, 5.784292, 5.784292, 5.784294, 5.784293, 5.784298, 
    5.784296, 5.784303, 5.784306, 5.784314, 5.784319, 5.784324, 5.784327, 
    5.784327, 5.784328 ;

 SOIL2C_TO_SOIL1C =
  1.302853e-09, 1.306423e-09, 1.305729e-09, 1.308607e-09, 1.307011e-09, 
    1.308895e-09, 1.303577e-09, 1.306564e-09, 1.304658e-09, 1.303175e-09, 
    1.31419e-09, 1.308736e-09, 1.319856e-09, 1.316379e-09, 1.325113e-09, 
    1.319315e-09, 1.326282e-09, 1.324946e-09, 1.328967e-09, 1.327816e-09, 
    1.332956e-09, 1.329499e-09, 1.335621e-09, 1.332131e-09, 1.332677e-09, 
    1.329385e-09, 1.309834e-09, 1.313511e-09, 1.309616e-09, 1.31014e-09, 
    1.309905e-09, 1.307044e-09, 1.305601e-09, 1.302581e-09, 1.303129e-09, 
    1.305348e-09, 1.310376e-09, 1.30867e-09, 1.312971e-09, 1.312874e-09, 
    1.317661e-09, 1.315503e-09, 1.323546e-09, 1.32126e-09, 1.327864e-09, 
    1.326203e-09, 1.327786e-09, 1.327306e-09, 1.327792e-09, 1.325357e-09, 
    1.3264e-09, 1.324257e-09, 1.315907e-09, 1.318361e-09, 1.311039e-09, 
    1.306634e-09, 1.303708e-09, 1.301631e-09, 1.301925e-09, 1.302485e-09, 
    1.305361e-09, 1.308065e-09, 1.310125e-09, 1.311503e-09, 1.31286e-09, 
    1.316967e-09, 1.319141e-09, 1.324007e-09, 1.32313e-09, 1.324617e-09, 
    1.326038e-09, 1.328423e-09, 1.328031e-09, 1.329081e-09, 1.324578e-09, 
    1.327571e-09, 1.32263e-09, 1.323981e-09, 1.313227e-09, 1.30913e-09, 
    1.307387e-09, 1.305862e-09, 1.302151e-09, 1.304714e-09, 1.303704e-09, 
    1.306108e-09, 1.307635e-09, 1.306879e-09, 1.31154e-09, 1.309728e-09, 
    1.31927e-09, 1.315161e-09, 1.325872e-09, 1.32331e-09, 1.326486e-09, 
    1.324866e-09, 1.327642e-09, 1.325144e-09, 1.329472e-09, 1.330414e-09, 
    1.329771e-09, 1.332244e-09, 1.325005e-09, 1.327785e-09, 1.306858e-09, 
    1.306981e-09, 1.307555e-09, 1.305032e-09, 1.304878e-09, 1.302566e-09, 
    1.304623e-09, 1.305499e-09, 1.307723e-09, 1.309038e-09, 1.310288e-09, 
    1.313037e-09, 1.316105e-09, 1.320395e-09, 1.323476e-09, 1.325541e-09, 
    1.324275e-09, 1.325393e-09, 1.324143e-09, 1.323558e-09, 1.330061e-09, 
    1.32641e-09, 1.331889e-09, 1.331586e-09, 1.329106e-09, 1.33162e-09, 
    1.307068e-09, 1.306359e-09, 1.303897e-09, 1.305824e-09, 1.302314e-09, 
    1.304279e-09, 1.305408e-09, 1.309766e-09, 1.310724e-09, 1.311611e-09, 
    1.313364e-09, 1.315613e-09, 1.319558e-09, 1.322989e-09, 1.326121e-09, 
    1.325891e-09, 1.325972e-09, 1.326671e-09, 1.324939e-09, 1.326956e-09, 
    1.327294e-09, 1.326409e-09, 1.331545e-09, 1.330078e-09, 1.331579e-09, 
    1.330624e-09, 1.30659e-09, 1.307782e-09, 1.307138e-09, 1.30835e-09, 
    1.307496e-09, 1.311291e-09, 1.312429e-09, 1.317753e-09, 1.315569e-09, 
    1.319045e-09, 1.315922e-09, 1.316475e-09, 1.319158e-09, 1.316091e-09, 
    1.322799e-09, 1.318251e-09, 1.326699e-09, 1.322157e-09, 1.326983e-09, 
    1.326107e-09, 1.327558e-09, 1.328856e-09, 1.33049e-09, 1.333504e-09, 
    1.332806e-09, 1.335327e-09, 1.30956e-09, 1.311107e-09, 1.310971e-09, 
    1.312589e-09, 1.313786e-09, 1.31638e-09, 1.320539e-09, 1.318975e-09, 
    1.321846e-09, 1.322422e-09, 1.318061e-09, 1.320738e-09, 1.312142e-09, 
    1.313531e-09, 1.312704e-09, 1.309682e-09, 1.319335e-09, 1.314382e-09, 
    1.323527e-09, 1.320845e-09, 1.328671e-09, 1.324779e-09, 1.332422e-09, 
    1.335687e-09, 1.338761e-09, 1.34235e-09, 1.311951e-09, 1.3109e-09, 
    1.312782e-09, 1.315384e-09, 1.317799e-09, 1.321008e-09, 1.321337e-09, 
    1.321938e-09, 1.323495e-09, 1.324804e-09, 1.322128e-09, 1.325132e-09, 
    1.313852e-09, 1.319765e-09, 1.310503e-09, 1.313292e-09, 1.315231e-09, 
    1.314381e-09, 1.318796e-09, 1.319837e-09, 1.324064e-09, 1.321879e-09, 
    1.334881e-09, 1.32913e-09, 1.345084e-09, 1.340627e-09, 1.310533e-09, 
    1.311947e-09, 1.316869e-09, 1.314527e-09, 1.321223e-09, 1.32287e-09, 
    1.324209e-09, 1.325921e-09, 1.326106e-09, 1.32712e-09, 1.325458e-09, 
    1.327054e-09, 1.321015e-09, 1.323714e-09, 1.316307e-09, 1.31811e-09, 
    1.31728e-09, 1.31637e-09, 1.319179e-09, 1.32217e-09, 1.322234e-09, 
    1.323193e-09, 1.325893e-09, 1.32125e-09, 1.335622e-09, 1.326747e-09, 
    1.31349e-09, 1.316213e-09, 1.316602e-09, 1.315547e-09, 1.322705e-09, 
    1.320112e-09, 1.327095e-09, 1.325208e-09, 1.3283e-09, 1.326763e-09, 
    1.326537e-09, 1.324564e-09, 1.323335e-09, 1.320231e-09, 1.317704e-09, 
    1.3157e-09, 1.316167e-09, 1.318367e-09, 1.322353e-09, 1.326122e-09, 
    1.325297e-09, 1.328065e-09, 1.320737e-09, 1.32381e-09, 1.322622e-09, 
    1.325719e-09, 1.318933e-09, 1.32471e-09, 1.317456e-09, 1.318092e-09, 
    1.320061e-09, 1.324018e-09, 1.324894e-09, 1.325829e-09, 1.325252e-09, 
    1.322454e-09, 1.321996e-09, 1.320013e-09, 1.319465e-09, 1.317954e-09, 
    1.316703e-09, 1.317846e-09, 1.319046e-09, 1.322455e-09, 1.325527e-09, 
    1.328875e-09, 1.329694e-09, 1.333603e-09, 1.33042e-09, 1.335671e-09, 
    1.331206e-09, 1.338936e-09, 1.325046e-09, 1.331076e-09, 1.32015e-09, 
    1.321328e-09, 1.323457e-09, 1.32834e-09, 1.325705e-09, 1.328787e-09, 
    1.321978e-09, 1.318443e-09, 1.317529e-09, 1.315822e-09, 1.317568e-09, 
    1.317426e-09, 1.319096e-09, 1.318559e-09, 1.322568e-09, 1.320415e-09, 
    1.326532e-09, 1.328763e-09, 1.335062e-09, 1.338922e-09, 1.342851e-09, 
    1.344585e-09, 1.345113e-09, 1.345334e-09 ;

 SOIL2C_TO_SOIL3C =
  9.306095e-11, 9.331591e-11, 9.326637e-11, 9.347194e-11, 9.335793e-11, 
    9.349252e-11, 9.311267e-11, 9.332601e-11, 9.318984e-11, 9.308394e-11, 
    9.387072e-11, 9.348113e-11, 9.427543e-11, 9.402705e-11, 9.465093e-11, 
    9.423677e-11, 9.473443e-11, 9.463903e-11, 9.492624e-11, 9.484397e-11, 
    9.521114e-11, 9.496421e-11, 9.540149e-11, 9.515221e-11, 9.519119e-11, 
    9.495606e-11, 9.355958e-11, 9.382221e-11, 9.354401e-11, 9.358146e-11, 
    9.356466e-11, 9.336026e-11, 9.325721e-11, 9.304149e-11, 9.308067e-11, 
    9.323912e-11, 9.359831e-11, 9.347642e-11, 9.378365e-11, 9.377672e-11, 
    9.411862e-11, 9.396448e-11, 9.453897e-11, 9.437574e-11, 9.48474e-11, 
    9.47288e-11, 9.484183e-11, 9.480756e-11, 9.484227e-11, 9.466833e-11, 
    9.474285e-11, 9.458979e-11, 9.399333e-11, 9.416865e-11, 9.364565e-11, 
    9.333099e-11, 9.312202e-11, 9.297368e-11, 9.299465e-11, 9.303462e-11, 
    9.324005e-11, 9.343319e-11, 9.358034e-11, 9.367875e-11, 9.377572e-11, 
    9.406906e-11, 9.422437e-11, 9.457195e-11, 9.450928e-11, 9.461549e-11, 
    9.471701e-11, 9.488735e-11, 9.485933e-11, 9.493437e-11, 9.461271e-11, 
    9.482649e-11, 9.447356e-11, 9.457009e-11, 9.380194e-11, 9.350931e-11, 
    9.338479e-11, 9.327589e-11, 9.301077e-11, 9.319385e-11, 9.312168e-11, 
    9.329339e-11, 9.340248e-11, 9.334854e-11, 9.368144e-11, 9.355203e-11, 
    9.423357e-11, 9.394007e-11, 9.470516e-11, 9.452214e-11, 9.474903e-11, 
    9.463327e-11, 9.48316e-11, 9.46531e-11, 9.496231e-11, 9.50296e-11, 
    9.498361e-11, 9.516032e-11, 9.464321e-11, 9.484181e-11, 9.334702e-11, 
    9.335582e-11, 9.339681e-11, 9.321659e-11, 9.320556e-11, 9.304042e-11, 
    9.318738e-11, 9.324994e-11, 9.340881e-11, 9.350274e-11, 9.359204e-11, 
    9.378833e-11, 9.400749e-11, 9.43139e-11, 9.453401e-11, 9.468151e-11, 
    9.459107e-11, 9.467091e-11, 9.458166e-11, 9.453983e-11, 9.500438e-11, 
    9.474355e-11, 9.513491e-11, 9.511326e-11, 9.493615e-11, 9.511569e-11, 
    9.336199e-11, 9.331137e-11, 9.313553e-11, 9.327314e-11, 9.302243e-11, 
    9.316276e-11, 9.324343e-11, 9.35547e-11, 9.362312e-11, 9.36865e-11, 
    9.381171e-11, 9.397236e-11, 9.425411e-11, 9.44992e-11, 9.472291e-11, 
    9.470653e-11, 9.471229e-11, 9.476225e-11, 9.463849e-11, 9.478256e-11, 
    9.480673e-11, 9.474353e-11, 9.511036e-11, 9.500557e-11, 9.51128e-11, 
    9.504458e-11, 9.332783e-11, 9.341301e-11, 9.336698e-11, 9.345354e-11, 
    9.339255e-11, 9.366367e-11, 9.374495e-11, 9.412519e-11, 9.396919e-11, 
    9.421749e-11, 9.399443e-11, 9.403395e-11, 9.422554e-11, 9.40065e-11, 
    9.448566e-11, 9.416078e-11, 9.476418e-11, 9.44398e-11, 9.478451e-11, 
    9.472195e-11, 9.482555e-11, 9.491831e-11, 9.503502e-11, 9.525029e-11, 
    9.520046e-11, 9.538048e-11, 9.354002e-11, 9.365047e-11, 9.364078e-11, 
    9.375637e-11, 9.384185e-11, 9.402713e-11, 9.432418e-11, 9.42125e-11, 
    9.441755e-11, 9.44587e-11, 9.414719e-11, 9.433844e-11, 9.372441e-11, 
    9.382362e-11, 9.376457e-11, 9.354872e-11, 9.42382e-11, 9.38844e-11, 
    9.453763e-11, 9.434606e-11, 9.490508e-11, 9.462708e-11, 9.517302e-11, 
    9.540622e-11, 9.562579e-11, 9.588218e-11, 9.371078e-11, 9.363573e-11, 
    9.377013e-11, 9.3956e-11, 9.41285e-11, 9.435774e-11, 9.43812e-11, 
    9.442414e-11, 9.453536e-11, 9.462885e-11, 9.443769e-11, 9.465229e-11, 
    9.384658e-11, 9.426891e-11, 9.360734e-11, 9.380656e-11, 9.394505e-11, 
    9.388433e-11, 9.419974e-11, 9.427405e-11, 9.457597e-11, 9.441992e-11, 
    9.534865e-11, 9.493787e-11, 9.607742e-11, 9.575909e-11, 9.36095e-11, 
    9.371053e-11, 9.406205e-11, 9.389482e-11, 9.437305e-11, 9.449072e-11, 
    9.458639e-11, 9.470862e-11, 9.472184e-11, 9.479426e-11, 9.467558e-11, 
    9.478958e-11, 9.435823e-11, 9.455101e-11, 9.402191e-11, 9.41507e-11, 
    9.409146e-11, 9.402646e-11, 9.422706e-11, 9.444068e-11, 9.444529e-11, 
    9.451377e-11, 9.470665e-11, 9.437499e-11, 9.540158e-11, 9.476765e-11, 
    9.382069e-11, 9.401519e-11, 9.404302e-11, 9.396767e-11, 9.447892e-11, 
    9.42937e-11, 9.47925e-11, 9.465773e-11, 9.487855e-11, 9.476882e-11, 
    9.475267e-11, 9.461174e-11, 9.452397e-11, 9.430219e-11, 9.412172e-11, 
    9.397861e-11, 9.40119e-11, 9.416909e-11, 9.445376e-11, 9.472301e-11, 
    9.466404e-11, 9.486176e-11, 9.433839e-11, 9.455786e-11, 9.447303e-11, 
    9.469422e-11, 9.420953e-11, 9.462216e-11, 9.4104e-11, 9.414945e-11, 
    9.429003e-11, 9.457272e-11, 9.463531e-11, 9.470207e-11, 9.466088e-11, 
    9.4461e-11, 9.442826e-11, 9.428662e-11, 9.424749e-11, 9.413956e-11, 
    9.405018e-11, 9.413183e-11, 9.421758e-11, 9.446109e-11, 9.468049e-11, 
    9.491962e-11, 9.497816e-11, 9.525736e-11, 9.503003e-11, 9.54051e-11, 
    9.508615e-11, 9.563825e-11, 9.464614e-11, 9.507684e-11, 9.429644e-11, 
    9.438055e-11, 9.453264e-11, 9.488143e-11, 9.469319e-11, 9.491335e-11, 
    9.442698e-11, 9.417449e-11, 9.410921e-11, 9.39873e-11, 9.4112e-11, 
    9.410185e-11, 9.422115e-11, 9.418282e-11, 9.446918e-11, 9.431537e-11, 
    9.475226e-11, 9.491163e-11, 9.53616e-11, 9.563731e-11, 9.591796e-11, 
    9.604181e-11, 9.607951e-11, 9.609526e-11 ;

 SOIL2C_vr =
  20.00613, 20.00614, 20.00614, 20.00615, 20.00614, 20.00615, 20.00613, 
    20.00614, 20.00613, 20.00613, 20.00618, 20.00615, 20.0062, 20.00619, 
    20.00622, 20.0062, 20.00623, 20.00622, 20.00624, 20.00624, 20.00626, 
    20.00624, 20.00627, 20.00625, 20.00626, 20.00624, 20.00616, 20.00617, 
    20.00616, 20.00616, 20.00616, 20.00614, 20.00614, 20.00612, 20.00613, 
    20.00614, 20.00616, 20.00615, 20.00617, 20.00617, 20.00619, 20.00618, 
    20.00622, 20.00621, 20.00624, 20.00623, 20.00624, 20.00623, 20.00624, 
    20.00623, 20.00623, 20.00622, 20.00618, 20.00619, 20.00616, 20.00614, 
    20.00613, 20.00612, 20.00612, 20.00612, 20.00614, 20.00615, 20.00616, 
    20.00616, 20.00617, 20.00619, 20.0062, 20.00622, 20.00621, 20.00622, 
    20.00623, 20.00624, 20.00624, 20.00624, 20.00622, 20.00624, 20.00621, 
    20.00622, 20.00617, 20.00615, 20.00615, 20.00614, 20.00612, 20.00613, 
    20.00613, 20.00614, 20.00615, 20.00614, 20.00616, 20.00616, 20.0062, 
    20.00618, 20.00623, 20.00622, 20.00623, 20.00622, 20.00624, 20.00622, 
    20.00624, 20.00625, 20.00624, 20.00625, 20.00622, 20.00624, 20.00614, 
    20.00614, 20.00615, 20.00614, 20.00613, 20.00612, 20.00613, 20.00614, 
    20.00615, 20.00615, 20.00616, 20.00617, 20.00618, 20.0062, 20.00622, 
    20.00623, 20.00622, 20.00623, 20.00622, 20.00622, 20.00624, 20.00623, 
    20.00625, 20.00625, 20.00624, 20.00625, 20.00614, 20.00614, 20.00613, 
    20.00614, 20.00612, 20.00613, 20.00614, 20.00616, 20.00616, 20.00616, 
    20.00617, 20.00618, 20.0062, 20.00621, 20.00623, 20.00623, 20.00623, 
    20.00623, 20.00622, 20.00623, 20.00623, 20.00623, 20.00625, 20.00624, 
    20.00625, 20.00625, 20.00614, 20.00615, 20.00615, 20.00615, 20.00615, 
    20.00616, 20.00617, 20.00619, 20.00618, 20.0062, 20.00618, 20.00619, 
    20.0062, 20.00618, 20.00621, 20.00619, 20.00623, 20.00621, 20.00623, 
    20.00623, 20.00624, 20.00624, 20.00625, 20.00626, 20.00626, 20.00627, 
    20.00616, 20.00616, 20.00616, 20.00617, 20.00617, 20.00619, 20.0062, 
    20.0062, 20.00621, 20.00621, 20.00619, 20.0062, 20.00617, 20.00617, 
    20.00617, 20.00616, 20.0062, 20.00618, 20.00622, 20.0062, 20.00624, 
    20.00622, 20.00626, 20.00627, 20.00628, 20.0063, 20.00617, 20.00616, 
    20.00617, 20.00618, 20.00619, 20.00621, 20.00621, 20.00621, 20.00622, 
    20.00622, 20.00621, 20.00622, 20.00617, 20.0062, 20.00616, 20.00617, 
    20.00618, 20.00618, 20.0062, 20.0062, 20.00622, 20.00621, 20.00627, 
    20.00624, 20.00631, 20.00629, 20.00616, 20.00617, 20.00619, 20.00618, 
    20.00621, 20.00621, 20.00622, 20.00623, 20.00623, 20.00623, 20.00623, 
    20.00623, 20.00621, 20.00622, 20.00619, 20.00619, 20.00619, 20.00619, 
    20.0062, 20.00621, 20.00621, 20.00622, 20.00623, 20.00621, 20.00627, 
    20.00623, 20.00617, 20.00619, 20.00619, 20.00618, 20.00621, 20.0062, 
    20.00623, 20.00622, 20.00624, 20.00623, 20.00623, 20.00622, 20.00622, 
    20.0062, 20.00619, 20.00618, 20.00618, 20.00619, 20.00621, 20.00623, 
    20.00622, 20.00624, 20.0062, 20.00622, 20.00621, 20.00623, 20.0062, 
    20.00622, 20.00619, 20.00619, 20.0062, 20.00622, 20.00622, 20.00623, 
    20.00622, 20.00621, 20.00621, 20.0062, 20.0062, 20.00619, 20.00619, 
    20.00619, 20.0062, 20.00621, 20.00623, 20.00624, 20.00624, 20.00626, 
    20.00625, 20.00627, 20.00625, 20.00628, 20.00622, 20.00625, 20.0062, 
    20.00621, 20.00622, 20.00624, 20.00623, 20.00624, 20.00621, 20.0062, 
    20.00619, 20.00618, 20.00619, 20.00619, 20.0062, 20.0062, 20.00621, 
    20.0062, 20.00623, 20.00624, 20.00627, 20.00628, 20.0063, 20.00631, 
    20.00631, 20.00631,
  20.00632, 20.00634, 20.00633, 20.00635, 20.00634, 20.00635, 20.00632, 
    20.00634, 20.00633, 20.00632, 20.00637, 20.00635, 20.0064, 20.00638, 
    20.00642, 20.0064, 20.00643, 20.00642, 20.00644, 20.00644, 20.00646, 
    20.00644, 20.00647, 20.00646, 20.00646, 20.00644, 20.00635, 20.00637, 
    20.00635, 20.00635, 20.00635, 20.00634, 20.00633, 20.00632, 20.00632, 
    20.00633, 20.00636, 20.00635, 20.00637, 20.00637, 20.00639, 20.00638, 
    20.00642, 20.0064, 20.00644, 20.00643, 20.00644, 20.00643, 20.00644, 
    20.00642, 20.00643, 20.00642, 20.00638, 20.00639, 20.00636, 20.00634, 
    20.00632, 20.00631, 20.00632, 20.00632, 20.00633, 20.00634, 20.00635, 
    20.00636, 20.00637, 20.00639, 20.0064, 20.00642, 20.00641, 20.00642, 
    20.00643, 20.00644, 20.00644, 20.00644, 20.00642, 20.00644, 20.00641, 
    20.00642, 20.00637, 20.00635, 20.00634, 20.00633, 20.00632, 20.00633, 
    20.00632, 20.00633, 20.00634, 20.00634, 20.00636, 20.00635, 20.0064, 
    20.00638, 20.00643, 20.00641, 20.00643, 20.00642, 20.00644, 20.00642, 
    20.00644, 20.00645, 20.00644, 20.00646, 20.00642, 20.00644, 20.00634, 
    20.00634, 20.00634, 20.00633, 20.00633, 20.00632, 20.00633, 20.00633, 
    20.00634, 20.00635, 20.00636, 20.00637, 20.00638, 20.0064, 20.00642, 
    20.00643, 20.00642, 20.00643, 20.00642, 20.00642, 20.00645, 20.00643, 
    20.00645, 20.00645, 20.00644, 20.00645, 20.00634, 20.00634, 20.00632, 
    20.00633, 20.00632, 20.00633, 20.00633, 20.00635, 20.00636, 20.00636, 
    20.00637, 20.00638, 20.0064, 20.00641, 20.00643, 20.00643, 20.00643, 
    20.00643, 20.00642, 20.00643, 20.00643, 20.00643, 20.00645, 20.00645, 
    20.00645, 20.00645, 20.00634, 20.00634, 20.00634, 20.00635, 20.00634, 
    20.00636, 20.00636, 20.00639, 20.00638, 20.0064, 20.00638, 20.00638, 
    20.0064, 20.00638, 20.00641, 20.00639, 20.00643, 20.00641, 20.00643, 
    20.00643, 20.00644, 20.00644, 20.00645, 20.00646, 20.00646, 20.00647, 
    20.00635, 20.00636, 20.00636, 20.00636, 20.00637, 20.00638, 20.0064, 
    20.0064, 20.00641, 20.00641, 20.00639, 20.0064, 20.00636, 20.00637, 
    20.00637, 20.00635, 20.0064, 20.00637, 20.00642, 20.0064, 20.00644, 
    20.00642, 20.00646, 20.00647, 20.00649, 20.0065, 20.00636, 20.00636, 
    20.00637, 20.00638, 20.00639, 20.0064, 20.00641, 20.00641, 20.00642, 
    20.00642, 20.00641, 20.00642, 20.00637, 20.0064, 20.00636, 20.00637, 
    20.00638, 20.00637, 20.00639, 20.0064, 20.00642, 20.00641, 20.00647, 
    20.00644, 20.00652, 20.0065, 20.00636, 20.00636, 20.00639, 20.00637, 
    20.0064, 20.00641, 20.00642, 20.00643, 20.00643, 20.00643, 20.00643, 
    20.00643, 20.0064, 20.00642, 20.00638, 20.00639, 20.00639, 20.00638, 
    20.0064, 20.00641, 20.00641, 20.00641, 20.00643, 20.0064, 20.00647, 
    20.00643, 20.00637, 20.00638, 20.00638, 20.00638, 20.00641, 20.0064, 
    20.00643, 20.00642, 20.00644, 20.00643, 20.00643, 20.00642, 20.00642, 
    20.0064, 20.00639, 20.00638, 20.00638, 20.00639, 20.00641, 20.00643, 
    20.00642, 20.00644, 20.0064, 20.00642, 20.00641, 20.00643, 20.0064, 
    20.00642, 20.00639, 20.00639, 20.0064, 20.00642, 20.00642, 20.00643, 
    20.00642, 20.00641, 20.00641, 20.0064, 20.0064, 20.00639, 20.00638, 
    20.00639, 20.0064, 20.00641, 20.00643, 20.00644, 20.00644, 20.00646, 
    20.00645, 20.00647, 20.00645, 20.00649, 20.00642, 20.00645, 20.0064, 
    20.00641, 20.00642, 20.00644, 20.00643, 20.00644, 20.00641, 20.00639, 
    20.00639, 20.00638, 20.00639, 20.00639, 20.0064, 20.00639, 20.00641, 
    20.0064, 20.00643, 20.00644, 20.00647, 20.00649, 20.00651, 20.00651, 
    20.00652, 20.00652,
  20.00634, 20.00636, 20.00636, 20.00637, 20.00636, 20.00637, 20.00634, 
    20.00636, 20.00635, 20.00634, 20.0064, 20.00637, 20.00642, 20.0064, 
    20.00645, 20.00642, 20.00645, 20.00644, 20.00646, 20.00646, 20.00648, 
    20.00647, 20.0065, 20.00648, 20.00648, 20.00647, 20.00637, 20.00639, 
    20.00637, 20.00637, 20.00637, 20.00636, 20.00635, 20.00634, 20.00634, 
    20.00635, 20.00638, 20.00637, 20.00639, 20.00639, 20.00641, 20.0064, 
    20.00644, 20.00643, 20.00646, 20.00645, 20.00646, 20.00646, 20.00646, 
    20.00645, 20.00645, 20.00644, 20.0064, 20.00641, 20.00638, 20.00636, 
    20.00635, 20.00633, 20.00634, 20.00634, 20.00635, 20.00636, 20.00637, 
    20.00638, 20.00639, 20.00641, 20.00642, 20.00644, 20.00644, 20.00644, 
    20.00645, 20.00646, 20.00646, 20.00646, 20.00644, 20.00646, 20.00643, 
    20.00644, 20.00639, 20.00637, 20.00636, 20.00636, 20.00634, 20.00635, 
    20.00635, 20.00636, 20.00636, 20.00636, 20.00638, 20.00637, 20.00642, 
    20.0064, 20.00645, 20.00644, 20.00645, 20.00644, 20.00646, 20.00645, 
    20.00647, 20.00647, 20.00647, 20.00648, 20.00644, 20.00646, 20.00636, 
    20.00636, 20.00636, 20.00635, 20.00635, 20.00634, 20.00635, 20.00635, 
    20.00636, 20.00637, 20.00638, 20.00639, 20.0064, 20.00642, 20.00644, 
    20.00645, 20.00644, 20.00645, 20.00644, 20.00644, 20.00647, 20.00645, 
    20.00648, 20.00648, 20.00646, 20.00648, 20.00636, 20.00636, 20.00635, 
    20.00636, 20.00634, 20.00635, 20.00635, 20.00637, 20.00638, 20.00638, 
    20.00639, 20.0064, 20.00642, 20.00644, 20.00645, 20.00645, 20.00645, 
    20.00645, 20.00644, 20.00645, 20.00646, 20.00645, 20.00648, 20.00647, 
    20.00648, 20.00647, 20.00636, 20.00636, 20.00636, 20.00637, 20.00636, 
    20.00638, 20.00639, 20.00641, 20.0064, 20.00642, 20.0064, 20.0064, 
    20.00642, 20.0064, 20.00644, 20.00641, 20.00645, 20.00643, 20.00645, 
    20.00645, 20.00646, 20.00646, 20.00647, 20.00648, 20.00648, 20.00649, 
    20.00637, 20.00638, 20.00638, 20.00639, 20.00639, 20.0064, 20.00642, 
    20.00642, 20.00643, 20.00643, 20.00641, 20.00643, 20.00638, 20.00639, 
    20.00639, 20.00637, 20.00642, 20.0064, 20.00644, 20.00643, 20.00646, 
    20.00644, 20.00648, 20.0065, 20.00651, 20.00653, 20.00638, 20.00638, 
    20.00639, 20.0064, 20.00641, 20.00643, 20.00643, 20.00643, 20.00644, 
    20.00644, 20.00643, 20.00645, 20.00639, 20.00642, 20.00638, 20.00639, 
    20.0064, 20.0064, 20.00642, 20.00642, 20.00644, 20.00643, 20.00649, 
    20.00647, 20.00654, 20.00652, 20.00638, 20.00638, 20.00641, 20.0064, 
    20.00643, 20.00644, 20.00644, 20.00645, 20.00645, 20.00646, 20.00645, 
    20.00645, 20.00643, 20.00644, 20.0064, 20.00641, 20.00641, 20.0064, 
    20.00642, 20.00643, 20.00643, 20.00644, 20.00645, 20.00643, 20.0065, 
    20.00645, 20.00639, 20.0064, 20.00641, 20.0064, 20.00644, 20.00642, 
    20.00645, 20.00645, 20.00646, 20.00645, 20.00645, 20.00644, 20.00644, 
    20.00642, 20.00641, 20.0064, 20.0064, 20.00641, 20.00643, 20.00645, 
    20.00645, 20.00646, 20.00643, 20.00644, 20.00643, 20.00645, 20.00642, 
    20.00644, 20.00641, 20.00641, 20.00642, 20.00644, 20.00644, 20.00645, 
    20.00645, 20.00643, 20.00643, 20.00642, 20.00642, 20.00641, 20.00641, 
    20.00641, 20.00642, 20.00643, 20.00645, 20.00646, 20.00647, 20.00649, 
    20.00647, 20.0065, 20.00648, 20.00651, 20.00644, 20.00647, 20.00642, 
    20.00643, 20.00644, 20.00646, 20.00645, 20.00646, 20.00643, 20.00641, 
    20.00641, 20.0064, 20.00641, 20.00641, 20.00642, 20.00641, 20.00643, 
    20.00642, 20.00645, 20.00646, 20.00649, 20.00651, 20.00653, 20.00654, 
    20.00654, 20.00654,
  20.00615, 20.00616, 20.00616, 20.00617, 20.00617, 20.00618, 20.00615, 
    20.00616, 20.00616, 20.00615, 20.0062, 20.00617, 20.00623, 20.00621, 
    20.00625, 20.00622, 20.00626, 20.00625, 20.00627, 20.00626, 20.00629, 
    20.00627, 20.0063, 20.00628, 20.00629, 20.00627, 20.00618, 20.0062, 
    20.00618, 20.00618, 20.00618, 20.00617, 20.00616, 20.00615, 20.00615, 
    20.00616, 20.00618, 20.00617, 20.0062, 20.00619, 20.00622, 20.00621, 
    20.00624, 20.00623, 20.00626, 20.00626, 20.00626, 20.00626, 20.00626, 
    20.00625, 20.00626, 20.00625, 20.00621, 20.00622, 20.00619, 20.00616, 
    20.00615, 20.00614, 20.00614, 20.00615, 20.00616, 20.00617, 20.00618, 
    20.00619, 20.00619, 20.00621, 20.00622, 20.00625, 20.00624, 20.00625, 
    20.00626, 20.00627, 20.00627, 20.00627, 20.00625, 20.00626, 20.00624, 
    20.00625, 20.0062, 20.00618, 20.00617, 20.00616, 20.00614, 20.00616, 
    20.00615, 20.00616, 20.00617, 20.00617, 20.00619, 20.00618, 20.00622, 
    20.0062, 20.00625, 20.00624, 20.00626, 20.00625, 20.00626, 20.00625, 
    20.00627, 20.00628, 20.00627, 20.00628, 20.00625, 20.00626, 20.00617, 
    20.00617, 20.00617, 20.00616, 20.00616, 20.00615, 20.00616, 20.00616, 
    20.00617, 20.00618, 20.00618, 20.0062, 20.00621, 20.00623, 20.00624, 
    20.00625, 20.00625, 20.00625, 20.00625, 20.00624, 20.00627, 20.00626, 
    20.00628, 20.00628, 20.00627, 20.00628, 20.00617, 20.00616, 20.00615, 
    20.00616, 20.00615, 20.00615, 20.00616, 20.00618, 20.00618, 20.00619, 
    20.0062, 20.00621, 20.00623, 20.00624, 20.00626, 20.00625, 20.00625, 
    20.00626, 20.00625, 20.00626, 20.00626, 20.00626, 20.00628, 20.00628, 
    20.00628, 20.00628, 20.00616, 20.00617, 20.00617, 20.00617, 20.00617, 
    20.00619, 20.00619, 20.00622, 20.00621, 20.00622, 20.00621, 20.00621, 
    20.00622, 20.00621, 20.00624, 20.00622, 20.00626, 20.00624, 20.00626, 
    20.00626, 20.00626, 20.00627, 20.00628, 20.00629, 20.00629, 20.0063, 
    20.00618, 20.00619, 20.00619, 20.00619, 20.0062, 20.00621, 20.00623, 
    20.00622, 20.00624, 20.00624, 20.00622, 20.00623, 20.00619, 20.0062, 
    20.00619, 20.00618, 20.00622, 20.0062, 20.00624, 20.00623, 20.00627, 
    20.00625, 20.00628, 20.0063, 20.00632, 20.00633, 20.00619, 20.00619, 
    20.00619, 20.00621, 20.00622, 20.00623, 20.00623, 20.00624, 20.00624, 
    20.00625, 20.00624, 20.00625, 20.0062, 20.00623, 20.00618, 20.0062, 
    20.0062, 20.0062, 20.00622, 20.00623, 20.00625, 20.00624, 20.0063, 
    20.00627, 20.00634, 20.00632, 20.00618, 20.00619, 20.00621, 20.0062, 
    20.00623, 20.00624, 20.00625, 20.00625, 20.00626, 20.00626, 20.00625, 
    20.00626, 20.00623, 20.00624, 20.00621, 20.00622, 20.00621, 20.00621, 
    20.00622, 20.00624, 20.00624, 20.00624, 20.00625, 20.00623, 20.0063, 
    20.00626, 20.0062, 20.00621, 20.00621, 20.00621, 20.00624, 20.00623, 
    20.00626, 20.00625, 20.00627, 20.00626, 20.00626, 20.00625, 20.00624, 
    20.00623, 20.00622, 20.00621, 20.00621, 20.00622, 20.00624, 20.00626, 
    20.00625, 20.00627, 20.00623, 20.00624, 20.00624, 20.00625, 20.00622, 
    20.00625, 20.00622, 20.00622, 20.00623, 20.00625, 20.00625, 20.00625, 
    20.00625, 20.00624, 20.00624, 20.00623, 20.00623, 20.00622, 20.00621, 
    20.00622, 20.00622, 20.00624, 20.00625, 20.00627, 20.00627, 20.00629, 
    20.00628, 20.0063, 20.00628, 20.00632, 20.00625, 20.00628, 20.00623, 
    20.00623, 20.00624, 20.00627, 20.00625, 20.00627, 20.00624, 20.00622, 
    20.00622, 20.00621, 20.00622, 20.00622, 20.00622, 20.00622, 20.00624, 
    20.00623, 20.00626, 20.00627, 20.0063, 20.00632, 20.00633, 20.00634, 
    20.00634, 20.00635,
  20.00526, 20.00528, 20.00527, 20.00529, 20.00528, 20.00529, 20.00526, 
    20.00528, 20.00527, 20.00526, 20.00531, 20.00529, 20.00533, 20.00532, 
    20.00535, 20.00533, 20.00536, 20.00535, 20.00537, 20.00537, 20.00539, 
    20.00537, 20.0054, 20.00538, 20.00539, 20.00537, 20.00529, 20.00531, 
    20.00529, 20.00529, 20.00529, 20.00528, 20.00527, 20.00526, 20.00526, 
    20.00527, 20.00529, 20.00529, 20.0053, 20.0053, 20.00532, 20.00531, 
    20.00535, 20.00534, 20.00537, 20.00536, 20.00537, 20.00536, 20.00537, 
    20.00536, 20.00536, 20.00535, 20.00532, 20.00533, 20.00529, 20.00528, 
    20.00527, 20.00526, 20.00526, 20.00526, 20.00527, 20.00528, 20.00529, 
    20.0053, 20.0053, 20.00532, 20.00533, 20.00535, 20.00535, 20.00535, 
    20.00536, 20.00537, 20.00537, 20.00537, 20.00535, 20.00537, 20.00534, 
    20.00535, 20.0053, 20.00529, 20.00528, 20.00527, 20.00526, 20.00527, 
    20.00527, 20.00528, 20.00528, 20.00528, 20.0053, 20.00529, 20.00533, 
    20.00531, 20.00536, 20.00535, 20.00536, 20.00535, 20.00537, 20.00535, 
    20.00537, 20.00538, 20.00537, 20.00538, 20.00535, 20.00537, 20.00528, 
    20.00528, 20.00528, 20.00527, 20.00527, 20.00526, 20.00527, 20.00527, 
    20.00528, 20.00529, 20.00529, 20.0053, 20.00532, 20.00533, 20.00535, 
    20.00536, 20.00535, 20.00536, 20.00535, 20.00535, 20.00537, 20.00536, 
    20.00538, 20.00538, 20.00537, 20.00538, 20.00528, 20.00528, 20.00527, 
    20.00527, 20.00526, 20.00527, 20.00527, 20.00529, 20.00529, 20.0053, 
    20.00531, 20.00531, 20.00533, 20.00535, 20.00536, 20.00536, 20.00536, 
    20.00536, 20.00535, 20.00536, 20.00536, 20.00536, 20.00538, 20.00537, 
    20.00538, 20.00538, 20.00528, 20.00528, 20.00528, 20.00529, 20.00528, 
    20.0053, 20.0053, 20.00532, 20.00531, 20.00533, 20.00532, 20.00532, 
    20.00533, 20.00532, 20.00534, 20.00533, 20.00536, 20.00534, 20.00536, 
    20.00536, 20.00536, 20.00537, 20.00538, 20.00539, 20.00539, 20.0054, 
    20.00529, 20.0053, 20.00529, 20.0053, 20.00531, 20.00532, 20.00533, 
    20.00533, 20.00534, 20.00534, 20.00533, 20.00534, 20.0053, 20.00531, 
    20.0053, 20.00529, 20.00533, 20.00531, 20.00535, 20.00534, 20.00537, 
    20.00535, 20.00538, 20.0054, 20.00541, 20.00543, 20.0053, 20.00529, 
    20.0053, 20.00531, 20.00532, 20.00534, 20.00534, 20.00534, 20.00535, 
    20.00535, 20.00534, 20.00535, 20.00531, 20.00533, 20.00529, 20.0053, 
    20.00531, 20.00531, 20.00533, 20.00533, 20.00535, 20.00534, 20.00539, 
    20.00537, 20.00544, 20.00542, 20.00529, 20.0053, 20.00532, 20.00531, 
    20.00534, 20.00534, 20.00535, 20.00536, 20.00536, 20.00536, 20.00536, 
    20.00536, 20.00534, 20.00535, 20.00532, 20.00533, 20.00532, 20.00532, 
    20.00533, 20.00534, 20.00534, 20.00535, 20.00536, 20.00534, 20.0054, 
    20.00536, 20.00531, 20.00532, 20.00532, 20.00531, 20.00534, 20.00533, 
    20.00536, 20.00535, 20.00537, 20.00536, 20.00536, 20.00535, 20.00535, 
    20.00533, 20.00532, 20.00532, 20.00532, 20.00533, 20.00534, 20.00536, 
    20.00536, 20.00537, 20.00534, 20.00535, 20.00534, 20.00536, 20.00533, 
    20.00535, 20.00532, 20.00533, 20.00533, 20.00535, 20.00535, 20.00536, 
    20.00535, 20.00534, 20.00534, 20.00533, 20.00533, 20.00533, 20.00532, 
    20.00532, 20.00533, 20.00534, 20.00536, 20.00537, 20.00537, 20.00539, 
    20.00538, 20.0054, 20.00538, 20.00541, 20.00535, 20.00538, 20.00533, 
    20.00534, 20.00535, 20.00537, 20.00536, 20.00537, 20.00534, 20.00533, 
    20.00532, 20.00532, 20.00532, 20.00532, 20.00533, 20.00533, 20.00534, 
    20.00533, 20.00536, 20.00537, 20.0054, 20.00541, 20.00543, 20.00544, 
    20.00544, 20.00544,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N =
  0.525843, 0.5258434, 0.5258433, 0.5258437, 0.5258435, 0.5258437, 0.5258431, 
    0.5258434, 0.5258432, 0.525843, 0.5258443, 0.5258437, 0.525845, 
    0.5258446, 0.5258456, 0.5258449, 0.5258457, 0.5258456, 0.5258461, 
    0.5258459, 0.5258465, 0.5258461, 0.5258468, 0.5258464, 0.5258465, 
    0.5258461, 0.5258438, 0.5258442, 0.5258438, 0.5258439, 0.5258438, 
    0.5258435, 0.5258433, 0.525843, 0.525843, 0.5258433, 0.5258439, 
    0.5258437, 0.5258442, 0.5258442, 0.5258448, 0.5258445, 0.5258454, 
    0.5258452, 0.5258459, 0.5258457, 0.5258459, 0.5258459, 0.5258459, 
    0.5258456, 0.5258458, 0.5258455, 0.5258445, 0.5258448, 0.525844, 
    0.5258434, 0.5258431, 0.5258428, 0.5258429, 0.525843, 0.5258433, 
    0.5258436, 0.5258439, 0.525844, 0.5258442, 0.5258446, 0.5258449, 
    0.5258455, 0.5258453, 0.5258455, 0.5258457, 0.525846, 0.5258459, 
    0.5258461, 0.5258455, 0.5258459, 0.5258453, 0.5258455, 0.5258442, 
    0.5258437, 0.5258435, 0.5258434, 0.5258429, 0.5258432, 0.5258431, 
    0.5258434, 0.5258436, 0.5258435, 0.525844, 0.5258438, 0.5258449, 
    0.5258445, 0.5258457, 0.5258454, 0.5258458, 0.5258456, 0.5258459, 
    0.5258456, 0.5258461, 0.5258462, 0.5258461, 0.5258464, 0.5258456, 
    0.5258459, 0.5258434, 0.5258435, 0.5258436, 0.5258433, 0.5258433, 
    0.525843, 0.5258432, 0.5258433, 0.5258436, 0.5258437, 0.5258439, 
    0.5258442, 0.5258446, 0.5258451, 0.5258454, 0.5258456, 0.5258455, 
    0.5258456, 0.5258455, 0.5258454, 0.5258462, 0.5258458, 0.5258464, 
    0.5258464, 0.5258461, 0.5258464, 0.5258435, 0.5258434, 0.5258431, 
    0.5258433, 0.525843, 0.5258431, 0.5258433, 0.5258438, 0.5258439, 
    0.525844, 0.5258442, 0.5258445, 0.5258449, 0.5258453, 0.5258457, 
    0.5258457, 0.5258457, 0.5258458, 0.5258456, 0.5258458, 0.5258458, 
    0.5258458, 0.5258464, 0.5258462, 0.5258464, 0.5258462, 0.5258434, 
    0.5258436, 0.5258435, 0.5258436, 0.5258436, 0.525844, 0.5258441, 
    0.5258448, 0.5258445, 0.5258449, 0.5258445, 0.5258446, 0.5258449, 
    0.5258446, 0.5258453, 0.5258448, 0.5258458, 0.5258452, 0.5258458, 
    0.5258457, 0.5258459, 0.5258461, 0.5258462, 0.5258466, 0.5258465, 
    0.5258468, 0.5258438, 0.525844, 0.525844, 0.5258442, 0.5258443, 
    0.5258446, 0.5258451, 0.5258449, 0.5258452, 0.5258453, 0.5258448, 
    0.5258451, 0.5258441, 0.5258443, 0.5258442, 0.5258438, 0.5258449, 
    0.5258443, 0.5258454, 0.5258451, 0.525846, 0.5258456, 0.5258465, 
    0.5258468, 0.5258472, 0.5258476, 0.525844, 0.5258439, 0.5258442, 
    0.5258445, 0.5258448, 0.5258451, 0.5258452, 0.5258452, 0.5258454, 
    0.5258456, 0.5258452, 0.5258456, 0.5258443, 0.525845, 0.5258439, 
    0.5258442, 0.5258445, 0.5258443, 0.5258449, 0.525845, 0.5258455, 
    0.5258452, 0.5258467, 0.5258461, 0.5258479, 0.5258474, 0.5258439, 
    0.525844, 0.5258446, 0.5258443, 0.5258452, 0.5258453, 0.5258455, 
    0.5258457, 0.5258457, 0.5258458, 0.5258456, 0.5258458, 0.5258451, 
    0.5258454, 0.5258446, 0.5258448, 0.5258447, 0.5258446, 0.5258449, 
    0.5258452, 0.5258453, 0.5258453, 0.5258457, 0.5258452, 0.5258468, 
    0.5258458, 0.5258442, 0.5258446, 0.5258446, 0.5258445, 0.5258453, 
    0.525845, 0.5258458, 0.5258456, 0.5258459, 0.5258458, 0.5258458, 
    0.5258455, 0.5258454, 0.5258451, 0.5258448, 0.5258445, 0.5258446, 
    0.5258448, 0.5258453, 0.5258457, 0.5258456, 0.5258459, 0.5258451, 
    0.5258455, 0.5258453, 0.5258456, 0.5258449, 0.5258455, 0.5258447, 
    0.5258448, 0.525845, 0.5258455, 0.5258456, 0.5258457, 0.5258456, 
    0.5258453, 0.5258452, 0.525845, 0.5258449, 0.5258448, 0.5258446, 
    0.5258448, 0.5258449, 0.5258453, 0.5258456, 0.5258461, 0.5258461, 
    0.5258466, 0.5258462, 0.5258468, 0.5258463, 0.5258472, 0.5258456, 
    0.5258463, 0.525845, 0.5258452, 0.5258454, 0.525846, 0.5258456, 0.525846, 
    0.5258452, 0.5258448, 0.5258447, 0.5258445, 0.5258447, 0.5258447, 
    0.5258449, 0.5258448, 0.5258453, 0.5258451, 0.5258458, 0.525846, 
    0.5258468, 0.5258472, 0.5258477, 0.5258479, 0.5258479, 0.525848 ;

 SOIL2N_TNDNCY_VERT_TRANS =
  -2.312965e-20, -1.28498e-20, 1.027984e-20, 0, -1.027984e-20, 7.709882e-21, 
    -2.569961e-21, 1.541976e-20, -7.709882e-21, -1.003089e-36, -2.055969e-20, 
    2.569961e-21, -1.003089e-36, 1.541976e-20, 1.027984e-20, 5.139921e-21, 
    -1.027984e-20, -1.003089e-36, -2.569961e-21, -2.569961e-20, 5.139921e-21, 
    2.312965e-20, 1.541976e-20, 2.569961e-21, 7.709882e-21, 2.569961e-21, 
    -2.055969e-20, 1.798972e-20, -7.709882e-21, 1.027984e-20, 1.027984e-20, 
    1.003089e-36, -2.312965e-20, 1.027984e-20, 1.28498e-20, -1.003089e-36, 
    1.003089e-36, 5.139921e-21, -1.027984e-20, 7.709882e-21, 1.28498e-20, 
    1.28498e-20, 1.541976e-20, 2.569961e-21, -5.139921e-21, 2.569961e-21, 
    5.139921e-21, 7.709882e-21, -1.003089e-36, -2.569961e-21, -1.541976e-20, 
    2.569961e-21, -7.709882e-21, 0, 0, 2.569961e-21, -1.027984e-20, 0, 
    5.139921e-21, 5.139921e-21, -1.027984e-20, 0, -1.027984e-20, 
    1.003089e-36, 5.139921e-21, -1.027984e-20, 2.569961e-21, 2.569961e-21, 
    -7.709882e-21, -2.569961e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, 
    -5.139921e-21, -7.709882e-21, 7.709882e-21, -1.798972e-20, -1.027984e-20, 
    -2.569961e-21, 7.709882e-21, -1.003089e-36, -1.027984e-20, 2.569961e-21, 
    -1.541976e-20, -5.139921e-21, -7.709882e-21, 1.027984e-20, -1.027984e-20, 
    -1.003089e-36, -1.798972e-20, 1.003089e-36, -2.569961e-21, 5.139921e-21, 
    -1.28498e-20, 2.569961e-21, 7.709882e-21, 1.28498e-20, -2.569961e-21, 
    -5.139921e-21, -7.709882e-21, 7.709882e-21, -5.139921e-21, 1.541976e-20, 
    -7.709882e-21, -1.003089e-36, 2.569961e-21, -2.569961e-21, -2.569961e-21, 
    -1.003089e-36, -1.28498e-20, -1.003089e-36, 1.28498e-20, 2.569961e-21, 
    -2.569961e-21, -1.027984e-20, 5.139921e-21, 0, -7.709882e-21, 
    -7.709882e-21, 0, 1.027984e-20, 5.139921e-21, -1.541976e-20, 
    -5.139921e-21, -1.003089e-36, 0, 1.28498e-20, 2.569961e-21, 5.139921e-21, 
    -7.709882e-21, -1.027984e-20, 1.28498e-20, -7.709882e-21, 2.569961e-21, 
    -1.28498e-20, 7.709882e-21, -7.709882e-21, -2.569961e-21, -2.569961e-21, 
    1.027984e-20, -1.003089e-36, 1.003089e-36, -1.003089e-36, 7.709882e-21, 
    2.569961e-21, 1.003089e-36, -1.798972e-20, 2.569961e-21, -1.027984e-20, 
    2.569961e-21, 2.569961e-21, 1.027984e-20, 1.798972e-20, 5.139921e-21, 
    -1.027984e-20, 1.28498e-20, -1.003089e-36, 1.003089e-36, -1.027984e-20, 
    0, 1.541976e-20, 1.003089e-36, 2.569961e-21, -2.569961e-21, 5.139921e-21, 
    -2.569961e-21, -1.027984e-20, 0, 1.027984e-20, 2.569961e-21, 
    -7.709882e-21, 2.569961e-21, 7.709882e-21, 2.569961e-21, -7.709882e-21, 
    -2.569961e-21, -5.139921e-21, -1.027984e-20, -7.709882e-21, 5.139921e-21, 
    1.027984e-20, -2.569961e-21, 7.709882e-21, -5.139921e-21, -1.027984e-20, 
    2.569961e-21, -2.312965e-20, 7.709882e-21, 1.027984e-20, 1.027984e-20, 
    -2.569961e-21, -2.569961e-21, -1.027984e-20, -5.139921e-21, 2.569961e-21, 
    2.055969e-20, 1.003089e-36, -2.826957e-20, -2.569961e-21, 1.798972e-20, 
    7.709882e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, -1.003089e-36, 
    7.709882e-21, 7.709882e-21, 5.139921e-21, 1.28498e-20, -1.027984e-20, 
    2.569961e-21, -5.139921e-21, 5.139921e-21, 1.003089e-36, -2.569961e-21, 
    -5.139921e-21, 1.027984e-20, 1.28498e-20, 1.28498e-20, -1.027984e-20, 0, 
    1.28498e-20, -1.027984e-20, -2.569961e-21, -2.569961e-21, 1.027984e-20, 
    -1.003089e-36, -2.569961e-21, -1.28498e-20, -2.569961e-21, -2.055969e-20, 
    -7.709882e-21, -1.541976e-20, -2.569961e-21, 1.798972e-20, -2.569961e-21, 
    1.28498e-20, -5.139921e-21, -2.569961e-21, -5.139921e-21, -1.003089e-36, 
    -7.709882e-21, 0, 2.569961e-21, -7.709882e-21, 2.569961e-21, 
    2.569961e-21, -5.139921e-21, 1.027984e-20, -5.139921e-21, -1.003089e-36, 
    -5.139921e-21, -2.569961e-21, -2.569961e-21, 0, 7.709882e-21, 
    -1.027984e-20, 1.28498e-20, 1.28498e-20, 5.139921e-21, 1.541976e-20, 
    -1.28498e-20, -2.569961e-21, 7.709882e-21, 2.569961e-21, -1.541976e-20, 
    -2.569961e-21, -5.139921e-21, 1.003089e-36, 1.003089e-36, -7.709882e-21, 
    -7.709882e-21, -1.003089e-36, 7.709882e-21, -2.312965e-20, 2.569961e-21, 
    -1.541976e-20, 2.569961e-21, -1.027984e-20, -2.569961e-21, -5.139921e-21, 
    7.709882e-21, -1.28498e-20, -2.569961e-21, 1.28498e-20, -2.569961e-21, 
    7.709882e-21, -2.569961e-21, -5.139921e-21, -7.709882e-21, -2.569961e-21, 
    -5.139921e-21, 5.139921e-21, 1.027984e-20, 5.139921e-21, -1.003089e-36, 
    1.027984e-20, 1.541976e-20, -1.027984e-20, 5.139921e-21, 0, 2.569961e-21, 
    -2.569961e-21, -1.027984e-20, 2.569961e-21, -1.541976e-20, 7.709882e-21, 
    -5.139921e-21, 5.139921e-21, -1.28498e-20, 2.569961e-21, 2.569961e-21, 
    -7.709882e-21, -2.569961e-21, -5.139921e-21, 5.139921e-21, -1.003089e-36, 
    2.055969e-20, -1.003089e-36, 0, 1.027984e-20, -5.139921e-21, 
    1.027984e-20, -5.139921e-21, -2.569961e-21, 2.569961e-21, -2.569961e-21, 
    1.003089e-36, -1.027984e-20, 1.027984e-20, -1.798972e-20, 7.709882e-21, 
    -2.055969e-20, 2.055969e-20, 1.798972e-20, 2.569961e-21, 2.569961e-21, 
    2.569961e-21,
  7.709882e-21, 1.28498e-20, 1.027984e-20, -1.003089e-36, 5.139921e-21, 0, 
    7.709882e-21, 1.027984e-20, -2.569961e-21, -2.569961e-21, 2.569961e-21, 
    5.139921e-21, 1.798972e-20, 1.28498e-20, 1.28498e-20, -5.139921e-21, 
    -7.709882e-21, -1.28498e-20, 2.569961e-21, -1.541976e-20, 2.569961e-21, 
    2.569961e-21, -5.139921e-21, -1.027984e-20, -7.709882e-21, -2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -5.139921e-21, 0, -7.709882e-21, 0, 
    5.139921e-21, 2.569961e-21, 1.003089e-36, 1.027984e-20, 2.312965e-20, 
    1.541976e-20, 1.003089e-36, 2.569961e-21, -7.709882e-21, 2.569961e-21, 
    -2.569961e-21, -7.709882e-21, -5.139921e-21, -7.709882e-21, 0, 
    -7.709882e-21, 5.139921e-21, 5.139921e-21, -1.027984e-20, -1.28498e-20, 
    -1.003089e-36, 5.139921e-21, 5.139921e-21, -7.709882e-21, -2.569961e-21, 
    -1.027984e-20, -1.28498e-20, 2.569961e-21, -2.569961e-21, -1.027984e-20, 
    -1.28498e-20, -2.569961e-21, -2.569961e-21, -5.139921e-21, -2.569961e-21, 
    -1.003089e-36, -7.709882e-21, 5.139921e-21, -1.027984e-20, 1.027984e-20, 
    -2.569961e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, -5.139921e-21, 
    -1.027984e-20, 1.027984e-20, -1.541976e-20, 7.709882e-21, 5.139921e-21, 
    -5.139921e-21, 1.28498e-20, 0, 1.28498e-20, -1.027984e-20, 0, 
    -1.541976e-20, 1.798972e-20, 7.709882e-21, -1.027984e-20, 2.569961e-21, 
    0, -1.28498e-20, 2.569961e-21, -7.709882e-21, 2.569961e-21, 5.139921e-21, 
    1.541976e-20, -2.569961e-21, -2.569961e-21, 7.709882e-21, -7.709882e-21, 
    5.139921e-21, -7.709882e-21, 1.541976e-20, -5.139921e-21, -2.569961e-21, 
    7.709882e-21, 7.709882e-21, 7.709882e-21, 2.569961e-21, 5.139921e-21, 
    1.003089e-36, 1.28498e-20, 5.139921e-21, 1.027984e-20, 1.027984e-20, 
    -2.569961e-21, 2.569961e-21, 5.139921e-21, -1.28498e-20, -5.139921e-21, 
    -1.027984e-20, -7.709882e-21, 0, 2.569961e-21, -2.569961e-21, 
    7.709882e-21, 0, 7.709882e-21, 1.28498e-20, 0, -7.709882e-21, 0, 
    2.569961e-21, 0, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    -5.139921e-21, -1.28498e-20, 2.569961e-21, -5.139921e-21, 2.569961e-21, 
    -2.569961e-21, 1.027984e-20, 2.569961e-21, -7.709882e-21, -1.003089e-36, 
    1.541976e-20, 5.139921e-21, 1.541976e-20, -5.139921e-21, -5.139921e-21, 
    5.139921e-21, -5.139921e-21, 0, 7.709882e-21, 0, -2.569961e-21, 
    7.709882e-21, 5.139921e-21, -2.569961e-21, -5.139921e-21, -5.139921e-21, 
    1.798972e-20, 2.569961e-21, 1.28498e-20, 0, 1.28498e-20, -1.027984e-20, 
    0, 7.709882e-21, -5.139921e-21, 5.139921e-21, 5.139921e-21, 0, 
    1.027984e-20, -1.003089e-36, -1.28498e-20, 1.003089e-36, 1.027984e-20, 
    7.709882e-21, -2.569961e-21, -1.28498e-20, 5.139921e-21, 5.139921e-21, 
    2.569961e-21, 7.709882e-21, 5.139921e-21, 7.709882e-21, -5.139921e-21, 
    2.312965e-20, 0, -5.139921e-21, 1.027984e-20, 7.709882e-21, 
    -5.139921e-21, -5.139921e-21, -2.569961e-21, 2.569961e-21, -1.541976e-20, 
    -5.139921e-21, 1.003089e-36, -1.28498e-20, -5.139921e-21, -2.569961e-21, 
    -2.569961e-21, -1.027984e-20, 5.139921e-21, 2.569961e-21, 7.709882e-21, 
    -5.139921e-21, 1.027984e-20, 5.139921e-21, 1.28498e-20, 5.139921e-21, 
    -5.139921e-21, 7.709882e-21, -1.027984e-20, 7.709882e-21, 7.709882e-21, 
    7.709882e-21, -1.027984e-20, 0, 1.28498e-20, 5.139921e-21, -1.027984e-20, 
    -1.541976e-20, 1.027984e-20, -1.027984e-20, -7.709882e-21, 1.027984e-20, 
    2.569961e-21, -2.569961e-21, 0, -1.28498e-20, 5.139921e-21, 
    -2.569961e-21, -7.709882e-21, 7.709882e-21, 7.709882e-21, 1.027984e-20, 
    2.569961e-21, -1.027984e-20, 1.003089e-36, -5.139921e-21, 2.569961e-21, 
    1.003089e-36, 0, 1.003089e-36, 2.569961e-21, -7.709882e-21, 
    -5.139921e-21, 1.28498e-20, 5.139921e-21, 1.541976e-20, -7.709882e-21, 
    7.709882e-21, 7.709882e-21, 1.027984e-20, -1.027984e-20, 2.569961e-21, 
    -1.003089e-36, -1.28498e-20, 0, -2.569961e-21, 0, -2.312965e-20, 
    -5.139921e-21, -1.027984e-20, -2.569961e-21, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, 5.139921e-21, -1.003089e-36, 0, 
    -1.28498e-20, -5.139921e-21, 0, 2.569961e-21, -7.709882e-21, 
    7.709882e-21, -1.541976e-20, 0, -7.709882e-21, -1.28498e-20, 
    -1.28498e-20, -2.569961e-21, -1.027984e-20, 5.139921e-21, 5.139921e-21, 
    -2.569961e-21, -7.709882e-21, -1.027984e-20, 1.003089e-36, -1.28498e-20, 
    -1.28498e-20, 2.569961e-21, -1.003089e-36, 1.003089e-36, -7.709882e-21, 
    7.709882e-21, 5.139921e-21, 0, 0, -2.569961e-21, -7.709882e-21, 
    -7.709882e-21, -1.003089e-36, -5.139921e-21, 0, 1.027984e-20, 
    7.709882e-21, -5.139921e-21, -7.709882e-21, -2.569961e-21, -2.569961e-21, 
    -7.709882e-21, -2.569961e-21, -5.139921e-21, -2.569961e-21, 7.709882e-21, 
    5.139921e-21, -1.027984e-20, -1.027984e-20, -5.139921e-21, 0, 
    -1.003089e-36, 5.139921e-21, 1.027984e-20, -7.709882e-21, 5.139921e-21, 
    0, -2.569961e-21,
  7.709882e-21, -2.569961e-21, 2.569961e-21, -1.003089e-36, -1.027984e-20, 
    2.055969e-20, 1.003089e-36, -5.139921e-21, 7.709882e-21, 1.798972e-20, 
    7.709882e-21, -5.139921e-21, -2.569961e-21, 5.139921e-21, 2.569961e-21, 
    -1.027984e-20, 1.027984e-20, 0, 1.798972e-20, 7.709882e-21, 5.139921e-21, 
    0, 1.28498e-20, -7.709882e-21, -1.027984e-20, -2.569961e-21, 0, 
    -5.139921e-21, 5.139921e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, 
    2.569961e-21, 1.003089e-36, -1.541976e-20, -2.569961e-21, 7.709882e-21, 
    -7.709882e-21, 0, -2.055969e-20, 2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 0, -5.139921e-21, -5.139921e-21, 7.709882e-21, 
    2.569961e-21, -1.541976e-20, -2.569961e-21, -5.139921e-21, -2.569961e-21, 
    -1.003089e-36, -1.28498e-20, -1.28498e-20, -2.569961e-21, 0, 
    2.569961e-21, 1.28498e-20, -5.139921e-21, 1.027984e-20, 1.027984e-20, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, 5.139921e-21, 2.569961e-21, 
    -2.569961e-21, -7.709882e-21, 0, 2.569961e-21, 2.569961e-21, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, -5.139921e-21, -2.569961e-21, 
    -7.709882e-21, 1.541976e-20, -5.139921e-21, 7.709882e-21, -2.569961e-21, 
    1.003089e-36, -1.027984e-20, -2.569961e-21, 5.139921e-21, 2.569961e-21, 
    1.28498e-20, 2.569961e-21, -7.709882e-21, 5.139921e-21, -5.139921e-21, 
    2.569961e-21, -1.28498e-20, 2.569961e-21, 2.569961e-21, 7.709882e-21, 
    -2.569961e-21, -7.709882e-21, 7.709882e-21, 5.139921e-21, -5.139921e-21, 
    1.003089e-36, -2.569961e-21, -1.798972e-20, -5.139921e-21, -5.139921e-21, 
    1.28498e-20, -1.28498e-20, 2.569961e-21, 5.139921e-21, -2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -1.027984e-20, -1.798972e-20, -1.027984e-20, 
    1.541976e-20, -1.027984e-20, 7.709882e-21, 1.798972e-20, -5.139921e-21, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, -2.569961e-21, -7.709882e-21, 
    5.139921e-21, -7.709882e-21, -1.798972e-20, 5.139921e-21, -1.027984e-20, 
    1.003089e-36, -1.28498e-20, -2.569961e-21, 7.709882e-21, -1.027984e-20, 
    -5.139921e-21, -1.003089e-36, -1.027984e-20, -7.709882e-21, 5.139921e-21, 
    -7.709882e-21, 2.569961e-21, -1.027984e-20, 2.569961e-21, 1.027984e-20, 
    2.569961e-21, -5.139921e-21, 5.139921e-21, -5.139921e-21, 0, 
    -1.28498e-20, -1.027984e-20, -1.027984e-20, 1.027984e-20, -5.139921e-21, 
    1.027984e-20, 1.28498e-20, -5.139921e-21, -5.139921e-21, -2.569961e-21, 
    1.003089e-36, -5.139921e-21, -5.139921e-21, -5.139921e-21, -2.569961e-21, 
    -1.28498e-20, -5.139921e-21, 1.027984e-20, -5.139921e-21, 7.709882e-21, 
    7.709882e-21, 5.139921e-21, -1.027984e-20, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 1.003089e-36, 7.709882e-21, 2.569961e-21, 0, 
    5.139921e-21, 0, 7.709882e-21, 7.709882e-21, -2.569961e-21, 
    -5.139921e-21, -7.709882e-21, -2.569961e-21, 7.709882e-21, -1.027984e-20, 
    1.541976e-20, -2.569961e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, 
    -2.312965e-20, 1.027984e-20, 1.027984e-20, 7.709882e-21, 7.709882e-21, 
    -2.569961e-21, 7.709882e-21, 7.709882e-21, -5.139921e-21, -7.709882e-21, 
    -1.027984e-20, 7.709882e-21, -5.139921e-21, -7.709882e-21, 0, 0, 
    2.569961e-21, 7.709882e-21, 1.003089e-36, -1.28498e-20, 2.569961e-21, 
    -2.569961e-21, -1.003089e-36, 5.139921e-21, -7.709882e-21, -1.003089e-36, 
    7.709882e-21, 5.139921e-21, -1.027984e-20, 7.709882e-21, 1.027984e-20, 
    -5.139921e-21, 0, -1.541976e-20, 0, -1.027984e-20, 1.027984e-20, 
    1.28498e-20, -7.709882e-21, -2.569961e-21, 5.139921e-21, -1.027984e-20, 
    2.569961e-21, 2.569961e-21, 0, 7.709882e-21, 2.569961e-21, -1.003089e-36, 
    -1.027984e-20, 0, -2.569961e-21, -1.027984e-20, -1.541976e-20, 
    1.027984e-20, 1.027984e-20, -7.709882e-21, -1.027984e-20, -5.139921e-21, 
    -5.139921e-21, -1.28498e-20, -7.709882e-21, -5.139921e-21, 1.027984e-20, 
    1.027984e-20, -5.139921e-21, 7.709882e-21, -2.569961e-21, -5.139921e-21, 
    -5.139921e-21, -7.709882e-21, 2.569961e-21, -2.055969e-20, -2.569961e-21, 
    1.027984e-20, 5.139921e-21, -2.569961e-21, -7.709882e-21, 1.28498e-20, 
    2.569961e-21, 5.139921e-21, -7.709882e-21, -1.027984e-20, -1.027984e-20, 
    -5.139921e-21, -1.027984e-20, -7.709882e-21, 5.139921e-21, -1.003089e-36, 
    1.003089e-36, -2.569961e-21, 7.709882e-21, 2.569961e-21, 5.139921e-21, 0, 
    -7.709882e-21, -2.569961e-21, 0, -5.139921e-21, 5.139921e-21, 
    2.569961e-21, 1.027984e-20, 1.027984e-20, -7.709882e-21, 5.139921e-21, 
    -1.541976e-20, -5.139921e-21, 7.709882e-21, 2.569961e-21, 1.003089e-36, 
    -7.709882e-21, 2.569961e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, 
    0, 1.003089e-36, 5.139921e-21, 2.569961e-21, -7.709882e-21, -1.28498e-20, 
    -1.027984e-20, 7.709882e-21, 2.569961e-21, 7.709882e-21, 5.139921e-21, 
    -1.28498e-20, 1.28498e-20, -2.569961e-21, -2.569961e-21, 0, 
    -2.569961e-21, 1.28498e-20, 5.139921e-21, -1.003089e-36, 0, 
    -7.709882e-21, -1.027984e-20, 1.027984e-20, 2.569961e-21, -7.709882e-21,
  -2.569961e-21, -2.569961e-21, -7.709882e-21, 0, -5.139921e-21, 
    -1.027984e-20, -2.055969e-20, -1.027984e-20, -5.139921e-21, 7.709882e-21, 
    7.709882e-21, -2.055969e-20, -2.569961e-21, -5.139921e-21, 1.28498e-20, 
    -2.569961e-21, 7.709882e-21, 1.003089e-36, -5.139921e-21, 1.28498e-20, 
    -5.139921e-21, 1.28498e-20, -2.312965e-20, 1.027984e-20, 7.709882e-21, 
    1.027984e-20, 7.709882e-21, 2.569961e-21, -7.709882e-21, -1.003089e-36, 
    -5.139921e-21, -1.28498e-20, -2.055969e-20, 5.139921e-21, -5.139921e-21, 
    0, -7.709882e-21, 2.569961e-21, -1.003089e-36, -2.569961e-21, 
    -1.027984e-20, 5.139921e-21, -7.709882e-21, 5.139921e-21, 7.709882e-21, 
    0, 1.28498e-20, 1.541976e-20, 1.541976e-20, 5.139921e-21, -5.139921e-21, 
    1.003089e-36, 0, 0, -2.569961e-21, 0, -5.139921e-21, -5.139921e-21, 
    1.28498e-20, 1.798972e-20, 1.027984e-20, 2.569961e-21, 2.569961e-21, 0, 
    -1.28498e-20, 1.28498e-20, -7.709882e-21, 0, 0, 2.569961e-21, 
    -2.569961e-21, -1.541976e-20, 7.709882e-21, -1.28498e-20, 7.709882e-21, 
    7.709882e-21, 5.139921e-21, -1.28498e-20, -2.312965e-20, -2.569961e-21, 
    -5.139921e-21, -1.541976e-20, -7.709882e-21, -1.28498e-20, -1.003089e-36, 
    -1.027984e-20, -7.709882e-21, -1.28498e-20, -2.569961e-21, 1.28498e-20, 
    -2.569961e-20, -5.139921e-21, 2.569961e-21, -2.569961e-21, -2.569961e-21, 
    0, 1.541976e-20, -2.569961e-21, 5.139921e-21, -5.139921e-21, 
    -7.709882e-21, -5.139921e-21, -7.709882e-21, 5.139921e-21, 7.709882e-21, 
    2.569961e-21, -7.709882e-21, -5.139921e-21, -1.541976e-20, 5.139921e-21, 
    -1.027984e-20, -5.139921e-21, 2.569961e-21, -1.798972e-20, -7.709882e-21, 
    -5.139921e-21, 2.569961e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, 
    -1.541976e-20, 5.139921e-21, 7.709882e-21, -2.569961e-21, -7.709882e-21, 
    -2.055969e-20, -7.709882e-21, 1.28498e-20, -7.709882e-21, 2.569961e-21, 
    2.569961e-21, 2.569961e-21, -1.027984e-20, -1.28498e-20, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, 1.027984e-20, 2.055969e-20, 1.798972e-20, 
    2.569961e-21, 1.28498e-20, -7.709882e-21, -1.28498e-20, -5.139921e-21, 
    -7.709882e-21, 2.569961e-21, 1.541976e-20, 2.569961e-21, -1.28498e-20, 
    2.569961e-21, 7.709882e-21, 5.139921e-21, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, 5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 7.709882e-21, -1.027984e-20, -2.569961e-21, 
    -1.027984e-20, 1.027984e-20, -5.139921e-21, -1.003089e-36, -2.569961e-21, 
    -2.569961e-21, 5.139921e-21, -1.027984e-20, -2.569961e-21, -7.709882e-21, 
    -5.139921e-21, 2.569961e-21, 1.798972e-20, -7.709882e-21, 2.569961e-21, 
    -2.055969e-20, 1.28498e-20, 2.569961e-21, -2.569961e-21, -7.709882e-21, 
    -5.139921e-21, 2.055969e-20, -1.798972e-20, -1.798972e-20, -1.003089e-36, 
    1.28498e-20, 7.709882e-21, -7.709882e-21, 2.569961e-20, 0, -7.709882e-21, 
    2.569961e-21, 0, -1.541976e-20, -7.709882e-21, -1.027984e-20, 
    2.569961e-21, 7.709882e-21, 7.709882e-21, 5.139921e-21, 5.139921e-21, 
    1.003089e-36, -7.709882e-21, -5.139921e-21, 1.003089e-36, 1.027984e-20, 
    2.826957e-20, 5.139921e-21, 1.003089e-36, 1.027984e-20, 2.569961e-21, 
    -7.709882e-21, -5.139921e-21, -7.709882e-21, 1.003089e-36, 1.28498e-20, 
    -2.569961e-21, 1.541976e-20, 2.569961e-21, 2.569961e-21, -7.709882e-21, 
    1.541976e-20, 7.709882e-21, 5.139921e-21, -5.139921e-21, 5.139921e-21, 
    -1.003089e-36, -2.569961e-21, -7.709882e-21, 1.027984e-20, 7.709882e-21, 
    7.709882e-21, 1.027984e-20, 1.027984e-20, -2.569961e-21, 0, 0, 
    2.055969e-20, 7.709882e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, 
    1.541976e-20, -2.569961e-21, 5.139921e-21, -5.139921e-21, 2.569961e-21, 
    -1.027984e-20, 2.569961e-21, -7.709882e-21, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, -2.569961e-21, -1.003089e-36, 5.139921e-21, -2.569961e-21, 
    -5.139921e-21, -1.027984e-20, -5.139921e-21, -1.003089e-36, 
    -2.312965e-20, -7.709882e-21, -2.569961e-21, 1.541976e-20, 1.027984e-20, 
    -7.709882e-21, 7.709882e-21, -1.28498e-20, -2.569961e-21, 1.798972e-20, 
    1.003089e-36, -2.569961e-21, 7.709882e-21, -7.709882e-21, -2.569961e-21, 
    -5.139921e-21, -1.027984e-20, -7.709882e-21, 1.027984e-20, 7.709882e-21, 
    0, -2.569961e-21, 1.28498e-20, -5.139921e-21, -1.027984e-20, 
    -1.798972e-20, -1.28498e-20, 1.027984e-20, -7.709882e-21, 1.28498e-20, 
    1.003089e-36, 1.541976e-20, 0, -2.569961e-21, 1.027984e-20, 
    -5.139921e-21, -2.569961e-21, 7.709882e-21, -7.709882e-21, -1.027984e-20, 
    -5.139921e-21, 1.798972e-20, 1.027984e-20, 1.027984e-20, -5.139921e-21, 
    -1.027984e-20, 5.139921e-21, 1.798972e-20, -1.027984e-20, 0, 
    -2.569961e-21, -1.28498e-20, -5.139921e-21, -7.709882e-21, 2.569961e-21, 
    -2.055969e-20, -1.798972e-20, 7.709882e-21, 1.027984e-20, -2.569961e-21, 
    2.055969e-20, -1.798972e-20, 7.709882e-21, -1.541976e-20, 5.139921e-21, 
    -5.139921e-21, -1.28498e-20, 1.027984e-20, -5.139921e-21, -1.027984e-20, 
    -7.709882e-21, -7.709882e-21,
  0, 1.027984e-20, -1.798972e-20, -1.28498e-20, 2.312965e-20, -7.709882e-21, 
    -2.055969e-20, 2.569961e-21, -5.139921e-21, -1.798972e-20, -1.28498e-20, 
    1.003089e-36, -1.798972e-20, -2.569961e-21, 1.027984e-20, 2.569961e-21, 
    1.027984e-20, 2.569961e-21, -5.139921e-21, -5.139921e-21, -7.709882e-21, 
    -7.709882e-21, 1.28498e-20, -7.709882e-21, -5.139921e-21, 2.312965e-20, 
    -1.798972e-20, -2.055969e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, 
    2.569961e-21, -5.139921e-21, 2.569961e-21, 5.139921e-21, 0, 
    -5.139921e-21, -2.569961e-21, -1.027984e-20, -7.709882e-21, 
    -5.139921e-21, 2.055969e-20, -7.709882e-21, -1.027984e-20, -1.28498e-20, 
    -5.139921e-21, -2.569961e-21, 7.709882e-21, 1.541976e-20, 5.139921e-21, 
    -1.003089e-36, -7.709882e-21, -5.139921e-21, -2.569961e-21, 2.055969e-20, 
    1.28498e-20, -2.826957e-20, 2.569961e-21, -1.003089e-36, 2.055969e-20, 
    1.28498e-20, 5.139921e-21, -7.709882e-21, 0, 1.003089e-36, 1.003089e-36, 
    1.28498e-20, 7.709882e-21, -1.28498e-20, -7.709882e-21, -5.139921e-21, 
    -1.28498e-20, 2.569961e-21, -2.569961e-21, -5.139921e-21, 5.139921e-21, 
    -1.798972e-20, -5.139921e-21, -2.055969e-20, -1.541976e-20, 1.541976e-20, 
    2.569961e-21, 7.709882e-21, 2.569961e-21, 7.709882e-21, -7.709882e-21, 
    -1.027984e-20, -1.28498e-20, 5.139921e-21, 7.709882e-21, 1.027984e-20, 
    -2.006177e-36, 2.569961e-20, -2.569961e-21, 5.139921e-21, 1.027984e-20, 
    2.569961e-21, -5.139921e-21, 1.027984e-20, 1.027984e-20, -1.798972e-20, 
    -1.28498e-20, -1.28498e-20, -7.709882e-21, -1.027984e-20, -1.027984e-20, 
    7.709882e-21, -2.569961e-21, 1.28498e-20, 2.569961e-21, 7.709882e-21, 
    1.28498e-20, 2.569961e-21, -1.027984e-20, -2.569961e-21, -5.139921e-21, 
    -1.027984e-20, 1.027984e-20, -1.027984e-20, 7.709882e-21, -7.709882e-21, 
    7.709882e-21, -2.569961e-21, -2.569961e-21, 2.055969e-20, 5.139921e-21, 
    2.569961e-21, -2.569961e-21, -5.139921e-21, 5.139921e-21, 2.569961e-21, 
    1.798972e-20, 5.139921e-21, 2.569961e-21, -7.709882e-21, 2.569961e-21, 
    5.139921e-21, -1.798972e-20, 5.139921e-21, 2.569961e-21, -1.798972e-20, 
    1.28498e-20, 1.798972e-20, 2.055969e-20, 7.709882e-21, -2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -2.569961e-21, -1.027984e-20, 7.709882e-21, 7.709882e-21, 1.28498e-20, 
    -1.28498e-20, -1.798972e-20, 0, 3.009266e-36, -7.709882e-21, 
    2.569961e-21, -2.569961e-21, -1.28498e-20, 2.569961e-21, -2.569961e-21, 
    -5.139921e-21, -5.139921e-21, 1.28498e-20, 1.541976e-20, 1.003089e-36, 
    -1.027984e-20, 1.798972e-20, 5.139921e-21, -1.798972e-20, 2.569961e-21, 
    5.139921e-21, -5.139921e-21, -1.003089e-36, -1.28498e-20, 0, 
    7.709882e-21, 2.569961e-21, -5.139921e-21, 5.139921e-21, 1.541976e-20, 
    1.027984e-20, 3.083953e-20, 2.569961e-21, 2.055969e-20, 7.709882e-21, 
    -1.027984e-20, -1.027984e-20, 1.027984e-20, 2.569961e-21, -1.027984e-20, 
    1.003089e-36, -1.28498e-20, -1.003089e-36, 7.709882e-21, 5.139921e-21, 
    -1.003089e-36, -2.569961e-21, 7.709882e-21, 2.569961e-21, -1.003089e-36, 
    7.709882e-21, 2.569961e-21, -1.28498e-20, 2.569961e-21, -2.569961e-21, 
    7.709882e-21, 1.541976e-20, 1.027984e-20, 5.139921e-21, 5.139921e-21, 
    -1.027984e-20, 7.709882e-21, -2.569961e-21, -5.139921e-21, -7.709882e-21, 
    1.798972e-20, 0, 1.027984e-20, 5.139921e-21, -5.139921e-21, 1.027984e-20, 
    0, -1.541976e-20, -5.139921e-21, 0, 2.312965e-20, 1.003089e-36, 
    1.541976e-20, 2.569961e-21, -2.569961e-21, -2.569961e-21, 1.027984e-20, 
    -1.003089e-36, -1.003089e-36, -7.709882e-21, 1.027984e-20, -1.541976e-20, 
    -2.569961e-21, 0, 1.541976e-20, 7.709882e-21, -5.139921e-21, 
    2.569961e-21, -7.709882e-21, 1.003089e-36, -7.709882e-21, -2.569961e-21, 
    -1.027984e-20, -7.709882e-21, 2.569961e-21, 2.569961e-21, 1.798972e-20, 
    2.055969e-20, 2.569961e-21, -7.709882e-21, -1.28498e-20, -7.709882e-21, 
    2.569961e-21, 5.139921e-21, 7.709882e-21, 1.027984e-20, -1.541976e-20, 
    2.569961e-21, 2.055969e-20, -1.28498e-20, -1.541976e-20, -7.709882e-21, 
    1.027984e-20, -1.027984e-20, 2.569961e-21, -7.709882e-21, -1.027984e-20, 
    -7.709882e-21, -2.569961e-21, 2.055969e-20, -2.569961e-21, 1.28498e-20, 
    5.139921e-21, 5.139921e-21, 2.569961e-21, 1.003089e-36, 2.569961e-21, 
    3.009266e-36, -5.139921e-21, -5.139921e-21, -5.139921e-21, 2.312965e-20, 
    5.139921e-21, -1.28498e-20, 1.003089e-36, 2.569961e-21, -7.709882e-21, 0, 
    -7.709882e-21, 7.709882e-21, -2.055969e-20, 2.055969e-20, 1.28498e-20, 
    -1.798972e-20, 5.139921e-21, -1.027984e-20, 7.709882e-21, -1.541976e-20, 
    1.027984e-20, 5.139921e-21, -5.139921e-21, 7.709882e-21, -1.541976e-20, 
    -2.569961e-21, -5.139921e-21, 7.709882e-21, -5.139921e-21, 7.709882e-21, 
    2.569961e-21, 5.139921e-21, 1.798972e-20, -5.139921e-21, -7.709882e-21, 
    1.28498e-20, -2.569961e-21, -1.28498e-20, 1.027984e-20, 2.569961e-21, 0, 
    5.139921e-21, -1.28498e-20, -5.139921e-21, -1.798972e-20, -5.139921e-21, 
    -1.027984e-20, 5.139921e-21, 1.003089e-36,
  6.259693e-29, 6.259697e-29, 6.259697e-29, 6.2597e-29, 6.259698e-29, 
    6.259701e-29, 6.259694e-29, 6.259698e-29, 6.259695e-29, 6.259693e-29, 
    6.259707e-29, 6.2597e-29, 6.259715e-29, 6.25971e-29, 6.259722e-29, 
    6.259714e-29, 6.259723e-29, 6.259721e-29, 6.259727e-29, 6.259725e-29, 
    6.259732e-29, 6.259727e-29, 6.259735e-29, 6.259731e-29, 6.259732e-29, 
    6.259727e-29, 6.259702e-29, 6.259707e-29, 6.259701e-29, 6.259702e-29, 
    6.259702e-29, 6.259698e-29, 6.259696e-29, 6.259692e-29, 6.259693e-29, 
    6.259696e-29, 6.259703e-29, 6.2597e-29, 6.259706e-29, 6.259706e-29, 
    6.259712e-29, 6.259709e-29, 6.259719e-29, 6.259716e-29, 6.259726e-29, 
    6.259723e-29, 6.259725e-29, 6.259724e-29, 6.259725e-29, 6.259722e-29, 
    6.259723e-29, 6.259721e-29, 6.25971e-29, 6.259713e-29, 6.259703e-29, 
    6.259698e-29, 6.259694e-29, 6.259691e-29, 6.259692e-29, 6.259692e-29, 
    6.259696e-29, 6.2597e-29, 6.259702e-29, 6.259704e-29, 6.259706e-29, 
    6.259711e-29, 6.259714e-29, 6.25972e-29, 6.259719e-29, 6.259721e-29, 
    6.259723e-29, 6.259726e-29, 6.259726e-29, 6.259727e-29, 6.259721e-29, 
    6.259725e-29, 6.259718e-29, 6.25972e-29, 6.259706e-29, 6.259701e-29, 
    6.259698e-29, 6.259697e-29, 6.259692e-29, 6.259695e-29, 6.259694e-29, 
    6.259697e-29, 6.259699e-29, 6.259698e-29, 6.259704e-29, 6.259701e-29, 
    6.259714e-29, 6.259709e-29, 6.259723e-29, 6.259719e-29, 6.259724e-29, 
    6.259721e-29, 6.259725e-29, 6.259722e-29, 6.259727e-29, 6.259729e-29, 
    6.259728e-29, 6.259731e-29, 6.259721e-29, 6.259725e-29, 6.259698e-29, 
    6.259698e-29, 6.259699e-29, 6.259695e-29, 6.259695e-29, 6.259692e-29, 
    6.259695e-29, 6.259696e-29, 6.259699e-29, 6.259701e-29, 6.259703e-29, 
    6.259706e-29, 6.25971e-29, 6.259715e-29, 6.259719e-29, 6.259723e-29, 
    6.259721e-29, 6.259722e-29, 6.259721e-29, 6.259719e-29, 6.259728e-29, 
    6.259723e-29, 6.25973e-29, 6.25973e-29, 6.259727e-29, 6.25973e-29, 
    6.259698e-29, 6.259697e-29, 6.259694e-29, 6.259697e-29, 6.259692e-29, 
    6.259695e-29, 6.259696e-29, 6.259701e-29, 6.259703e-29, 6.259704e-29, 
    6.259706e-29, 6.259709e-29, 6.259715e-29, 6.259719e-29, 6.259723e-29, 
    6.259723e-29, 6.259723e-29, 6.259724e-29, 6.259721e-29, 6.259724e-29, 
    6.259724e-29, 6.259723e-29, 6.25973e-29, 6.259728e-29, 6.25973e-29, 
    6.259729e-29, 6.259698e-29, 6.259699e-29, 6.259698e-29, 6.2597e-29, 
    6.259699e-29, 6.259704e-29, 6.259705e-29, 6.259712e-29, 6.259709e-29, 
    6.259714e-29, 6.25971e-29, 6.25971e-29, 6.259714e-29, 6.25971e-29, 
    6.259719e-29, 6.259713e-29, 6.259724e-29, 6.259718e-29, 6.259724e-29, 
    6.259723e-29, 6.259725e-29, 6.259727e-29, 6.259729e-29, 6.259733e-29, 
    6.259732e-29, 6.259735e-29, 6.259701e-29, 6.259703e-29, 6.259703e-29, 
    6.259706e-29, 6.259707e-29, 6.25971e-29, 6.259716e-29, 6.259713e-29, 
    6.259718e-29, 6.259718e-29, 6.259712e-29, 6.259716e-29, 6.259705e-29, 
    6.259707e-29, 6.259706e-29, 6.259701e-29, 6.259714e-29, 6.259707e-29, 
    6.259719e-29, 6.259716e-29, 6.259726e-29, 6.259721e-29, 6.259731e-29, 
    6.259736e-29, 6.259739e-29, 6.259744e-29, 6.259704e-29, 6.259703e-29, 
    6.259706e-29, 6.259709e-29, 6.259712e-29, 6.259716e-29, 6.259716e-29, 
    6.259718e-29, 6.259719e-29, 6.259721e-29, 6.259718e-29, 6.259722e-29, 
    6.259707e-29, 6.259715e-29, 6.259703e-29, 6.259706e-29, 6.259709e-29, 
    6.259707e-29, 6.259713e-29, 6.259715e-29, 6.25972e-29, 6.259718e-29, 
    6.259735e-29, 6.259727e-29, 6.259748e-29, 6.259742e-29, 6.259703e-29, 
    6.259704e-29, 6.259711e-29, 6.259708e-29, 6.259716e-29, 6.259719e-29, 
    6.259721e-29, 6.259723e-29, 6.259723e-29, 6.259724e-29, 6.259722e-29, 
    6.259724e-29, 6.259716e-29, 6.25972e-29, 6.25971e-29, 6.259712e-29, 
    6.259712e-29, 6.25971e-29, 6.259714e-29, 6.259718e-29, 6.259718e-29, 
    6.259719e-29, 6.259723e-29, 6.259716e-29, 6.259735e-29, 6.259724e-29, 
    6.259707e-29, 6.25971e-29, 6.25971e-29, 6.259709e-29, 6.259718e-29, 
    6.259715e-29, 6.259724e-29, 6.259722e-29, 6.259726e-29, 6.259724e-29, 
    6.259724e-29, 6.259721e-29, 6.259719e-29, 6.259715e-29, 6.259712e-29, 
    6.259709e-29, 6.25971e-29, 6.259713e-29, 6.259718e-29, 6.259723e-29, 
    6.259722e-29, 6.259726e-29, 6.259716e-29, 6.25972e-29, 6.259718e-29, 
    6.259723e-29, 6.259713e-29, 6.259721e-29, 6.259712e-29, 6.259712e-29, 
    6.259715e-29, 6.25972e-29, 6.259721e-29, 6.259723e-29, 6.259722e-29, 
    6.259718e-29, 6.259718e-29, 6.259715e-29, 6.259714e-29, 6.259712e-29, 
    6.25971e-29, 6.259712e-29, 6.259714e-29, 6.259718e-29, 6.259723e-29, 
    6.259727e-29, 6.259728e-29, 6.259733e-29, 6.259729e-29, 6.259735e-29, 
    6.25973e-29, 6.25974e-29, 6.259721e-29, 6.25973e-29, 6.259715e-29, 
    6.259716e-29, 6.259719e-29, 6.259726e-29, 6.259723e-29, 6.259727e-29, 
    6.259718e-29, 6.259713e-29, 6.259712e-29, 6.25971e-29, 6.259712e-29, 
    6.259712e-29, 6.259714e-29, 6.259713e-29, 6.259718e-29, 6.259715e-29, 
    6.259724e-29, 6.259727e-29, 6.259735e-29, 6.25974e-29, 6.259745e-29, 
    6.259747e-29, 6.259748e-29, 6.259748e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N_TO_SOIL1N =
  2.632027e-10, 2.639238e-10, 2.637837e-10, 2.643651e-10, 2.640426e-10, 
    2.644233e-10, 2.63349e-10, 2.639524e-10, 2.635672e-10, 2.632677e-10, 
    2.65493e-10, 2.643911e-10, 2.666376e-10, 2.659351e-10, 2.676996e-10, 
    2.665282e-10, 2.679358e-10, 2.676659e-10, 2.684782e-10, 2.682456e-10, 
    2.69284e-10, 2.685857e-10, 2.698224e-10, 2.691173e-10, 2.692276e-10, 
    2.685626e-10, 2.646129e-10, 2.653558e-10, 2.645689e-10, 2.646748e-10, 
    2.646273e-10, 2.640492e-10, 2.637578e-10, 2.631477e-10, 2.632584e-10, 
    2.637066e-10, 2.647225e-10, 2.643778e-10, 2.652467e-10, 2.652271e-10, 
    2.661941e-10, 2.657581e-10, 2.673829e-10, 2.669213e-10, 2.682553e-10, 
    2.679199e-10, 2.682395e-10, 2.681426e-10, 2.682408e-10, 2.677488e-10, 
    2.679596e-10, 2.675267e-10, 2.658397e-10, 2.663356e-10, 2.648564e-10, 
    2.639664e-10, 2.633754e-10, 2.629559e-10, 2.630152e-10, 2.631282e-10, 
    2.637092e-10, 2.642555e-10, 2.646717e-10, 2.6495e-10, 2.652243e-10, 
    2.660539e-10, 2.664932e-10, 2.674762e-10, 2.67299e-10, 2.675994e-10, 
    2.678865e-10, 2.683683e-10, 2.68289e-10, 2.685012e-10, 2.675915e-10, 
    2.681961e-10, 2.671979e-10, 2.67471e-10, 2.652984e-10, 2.644708e-10, 
    2.641186e-10, 2.638106e-10, 2.630608e-10, 2.635786e-10, 2.633745e-10, 
    2.638601e-10, 2.641686e-10, 2.640161e-10, 2.649576e-10, 2.645916e-10, 
    2.665192e-10, 2.656891e-10, 2.67853e-10, 2.673353e-10, 2.679771e-10, 
    2.676497e-10, 2.682106e-10, 2.677057e-10, 2.685803e-10, 2.687706e-10, 
    2.686405e-10, 2.691403e-10, 2.676778e-10, 2.682395e-10, 2.640118e-10, 
    2.640367e-10, 2.641526e-10, 2.636429e-10, 2.636117e-10, 2.631446e-10, 
    2.635603e-10, 2.637372e-10, 2.641865e-10, 2.644522e-10, 2.647047e-10, 
    2.652599e-10, 2.658798e-10, 2.667464e-10, 2.673689e-10, 2.677861e-10, 
    2.675303e-10, 2.677561e-10, 2.675037e-10, 2.673854e-10, 2.686993e-10, 
    2.679615e-10, 2.690684e-10, 2.690072e-10, 2.685063e-10, 2.690141e-10, 
    2.640541e-10, 2.639109e-10, 2.634136e-10, 2.638028e-10, 2.630937e-10, 
    2.634906e-10, 2.637188e-10, 2.645991e-10, 2.647926e-10, 2.649719e-10, 
    2.65326e-10, 2.657804e-10, 2.665773e-10, 2.672705e-10, 2.679032e-10, 
    2.678568e-10, 2.678732e-10, 2.680144e-10, 2.676644e-10, 2.680719e-10, 
    2.681403e-10, 2.679615e-10, 2.68999e-10, 2.687026e-10, 2.690059e-10, 
    2.688129e-10, 2.639575e-10, 2.641984e-10, 2.640682e-10, 2.64313e-10, 
    2.641405e-10, 2.649073e-10, 2.651372e-10, 2.662127e-10, 2.657715e-10, 
    2.664737e-10, 2.658428e-10, 2.659546e-10, 2.664965e-10, 2.65877e-10, 
    2.672322e-10, 2.663133e-10, 2.680199e-10, 2.671025e-10, 2.680774e-10, 
    2.679005e-10, 2.681935e-10, 2.684558e-10, 2.687859e-10, 2.693948e-10, 
    2.692538e-10, 2.69763e-10, 2.645576e-10, 2.6487e-10, 2.648426e-10, 
    2.651696e-10, 2.654113e-10, 2.659353e-10, 2.667755e-10, 2.664596e-10, 
    2.670395e-10, 2.671559e-10, 2.662749e-10, 2.668158e-10, 2.650792e-10, 
    2.653597e-10, 2.651927e-10, 2.645822e-10, 2.665323e-10, 2.655317e-10, 
    2.673792e-10, 2.668373e-10, 2.684184e-10, 2.676322e-10, 2.691762e-10, 
    2.698358e-10, 2.704568e-10, 2.711819e-10, 2.650406e-10, 2.648283e-10, 
    2.652084e-10, 2.657341e-10, 2.66222e-10, 2.668704e-10, 2.669368e-10, 
    2.670582e-10, 2.673727e-10, 2.676372e-10, 2.670965e-10, 2.677034e-10, 
    2.654247e-10, 2.666191e-10, 2.64748e-10, 2.653115e-10, 2.657032e-10, 
    2.655314e-10, 2.664235e-10, 2.666337e-10, 2.674876e-10, 2.670462e-10, 
    2.69673e-10, 2.685111e-10, 2.717341e-10, 2.708338e-10, 2.647541e-10, 
    2.650399e-10, 2.660341e-10, 2.655611e-10, 2.669137e-10, 2.672465e-10, 
    2.675171e-10, 2.678628e-10, 2.679001e-10, 2.68105e-10, 2.677693e-10, 
    2.680917e-10, 2.668717e-10, 2.67417e-10, 2.659205e-10, 2.662848e-10, 
    2.661173e-10, 2.659334e-10, 2.665008e-10, 2.67105e-10, 2.67118e-10, 
    2.673117e-10, 2.678572e-10, 2.669192e-10, 2.698226e-10, 2.680297e-10, 
    2.653515e-10, 2.659016e-10, 2.659803e-10, 2.657672e-10, 2.672131e-10, 
    2.666893e-10, 2.681e-10, 2.677188e-10, 2.683434e-10, 2.68033e-10, 
    2.679874e-10, 2.675888e-10, 2.673405e-10, 2.667133e-10, 2.662028e-10, 
    2.657981e-10, 2.658922e-10, 2.663368e-10, 2.67142e-10, 2.679035e-10, 
    2.677367e-10, 2.682959e-10, 2.668157e-10, 2.674364e-10, 2.671965e-10, 
    2.67822e-10, 2.664512e-10, 2.676182e-10, 2.661527e-10, 2.662813e-10, 
    2.666789e-10, 2.674784e-10, 2.676554e-10, 2.678442e-10, 2.677278e-10, 
    2.671624e-10, 2.670698e-10, 2.666692e-10, 2.665586e-10, 2.662533e-10, 
    2.660005e-10, 2.662315e-10, 2.66474e-10, 2.671627e-10, 2.677832e-10, 
    2.684595e-10, 2.686251e-10, 2.694148e-10, 2.687718e-10, 2.698326e-10, 
    2.689305e-10, 2.70492e-10, 2.67686e-10, 2.689042e-10, 2.66697e-10, 
    2.669349e-10, 2.67365e-10, 2.683515e-10, 2.678191e-10, 2.684418e-10, 
    2.670662e-10, 2.663521e-10, 2.661674e-10, 2.658227e-10, 2.661753e-10, 
    2.661467e-10, 2.664841e-10, 2.663756e-10, 2.671856e-10, 2.667506e-10, 
    2.679862e-10, 2.684369e-10, 2.697096e-10, 2.704894e-10, 2.712831e-10, 
    2.716334e-10, 2.7174e-10, 2.717846e-10 ;

 SOIL2N_TO_SOIL3N =
  1.880019e-11, 1.88517e-11, 1.884169e-11, 1.888322e-11, 1.886019e-11, 
    1.888738e-11, 1.881064e-11, 1.885374e-11, 1.882623e-11, 1.880483e-11, 
    1.896378e-11, 1.888508e-11, 1.904554e-11, 1.899536e-11, 1.91214e-11, 
    1.903773e-11, 1.913827e-11, 1.9119e-11, 1.917702e-11, 1.91604e-11, 
    1.923458e-11, 1.918469e-11, 1.927303e-11, 1.922267e-11, 1.923054e-11, 
    1.918304e-11, 1.890092e-11, 1.895398e-11, 1.889778e-11, 1.890535e-11, 
    1.890195e-11, 1.886066e-11, 1.883984e-11, 1.879626e-11, 1.880418e-11, 
    1.883619e-11, 1.890875e-11, 1.888413e-11, 1.894619e-11, 1.894479e-11, 
    1.901386e-11, 1.898272e-11, 1.909878e-11, 1.906581e-11, 1.916109e-11, 
    1.913713e-11, 1.915997e-11, 1.915304e-11, 1.916006e-11, 1.912492e-11, 
    1.913997e-11, 1.910905e-11, 1.898855e-11, 1.902397e-11, 1.891831e-11, 
    1.885474e-11, 1.881253e-11, 1.878256e-11, 1.87868e-11, 1.879487e-11, 
    1.883638e-11, 1.887539e-11, 1.890512e-11, 1.8925e-11, 1.894459e-11, 
    1.900385e-11, 1.903523e-11, 1.910544e-11, 1.909278e-11, 1.911424e-11, 
    1.913475e-11, 1.916916e-11, 1.91635e-11, 1.917866e-11, 1.911368e-11, 
    1.915687e-11, 1.908557e-11, 1.910507e-11, 1.894989e-11, 1.889077e-11, 
    1.886561e-11, 1.884361e-11, 1.879005e-11, 1.882704e-11, 1.881246e-11, 
    1.884715e-11, 1.886919e-11, 1.885829e-11, 1.892555e-11, 1.88994e-11, 
    1.903708e-11, 1.897779e-11, 1.913236e-11, 1.909538e-11, 1.914122e-11, 
    1.911783e-11, 1.91579e-11, 1.912184e-11, 1.91843e-11, 1.91979e-11, 
    1.918861e-11, 1.922431e-11, 1.911984e-11, 1.915996e-11, 1.885798e-11, 
    1.885976e-11, 1.886804e-11, 1.883163e-11, 1.882941e-11, 1.879604e-11, 
    1.882573e-11, 1.883837e-11, 1.887047e-11, 1.888944e-11, 1.890748e-11, 
    1.894714e-11, 1.899141e-11, 1.905331e-11, 1.909778e-11, 1.912758e-11, 
    1.910931e-11, 1.912544e-11, 1.91074e-11, 1.909896e-11, 1.91928e-11, 
    1.914011e-11, 1.921917e-11, 1.92148e-11, 1.917902e-11, 1.921529e-11, 
    1.886101e-11, 1.885078e-11, 1.881526e-11, 1.884306e-11, 1.879241e-11, 
    1.882076e-11, 1.883706e-11, 1.889994e-11, 1.891376e-11, 1.892657e-11, 
    1.895186e-11, 1.898432e-11, 1.904124e-11, 1.909075e-11, 1.913594e-11, 
    1.913263e-11, 1.91338e-11, 1.914389e-11, 1.911889e-11, 1.914799e-11, 
    1.915288e-11, 1.914011e-11, 1.921421e-11, 1.919304e-11, 1.921471e-11, 
    1.920093e-11, 1.885411e-11, 1.887132e-11, 1.886202e-11, 1.88795e-11, 
    1.886718e-11, 1.892195e-11, 1.893837e-11, 1.901519e-11, 1.898368e-11, 
    1.903384e-11, 1.898877e-11, 1.899676e-11, 1.903546e-11, 1.899121e-11, 
    1.908801e-11, 1.902238e-11, 1.914428e-11, 1.907875e-11, 1.914839e-11, 
    1.913575e-11, 1.915668e-11, 1.917542e-11, 1.919899e-11, 1.924248e-11, 
    1.923242e-11, 1.926878e-11, 1.889697e-11, 1.891929e-11, 1.891733e-11, 
    1.894068e-11, 1.895795e-11, 1.899538e-11, 1.905539e-11, 1.903283e-11, 
    1.907425e-11, 1.908257e-11, 1.901963e-11, 1.905827e-11, 1.893422e-11, 
    1.895427e-11, 1.894234e-11, 1.889873e-11, 1.903802e-11, 1.896655e-11, 
    1.909851e-11, 1.905981e-11, 1.917274e-11, 1.911658e-11, 1.922687e-11, 
    1.927399e-11, 1.931834e-11, 1.937014e-11, 1.893147e-11, 1.891631e-11, 
    1.894346e-11, 1.898101e-11, 1.901586e-11, 1.906217e-11, 1.906691e-11, 
    1.907558e-11, 1.909805e-11, 1.911694e-11, 1.907832e-11, 1.912167e-11, 
    1.89589e-11, 1.904422e-11, 1.891057e-11, 1.895082e-11, 1.89788e-11, 
    1.896653e-11, 1.903025e-11, 1.904526e-11, 1.910626e-11, 1.907473e-11, 
    1.926235e-11, 1.917937e-11, 1.940958e-11, 1.934527e-11, 1.891101e-11, 
    1.893142e-11, 1.900243e-11, 1.896865e-11, 1.906526e-11, 1.908903e-11, 
    1.910836e-11, 1.913305e-11, 1.913573e-11, 1.915035e-11, 1.912638e-11, 
    1.914941e-11, 1.906227e-11, 1.910122e-11, 1.899433e-11, 1.902034e-11, 
    1.900838e-11, 1.899524e-11, 1.903577e-11, 1.907893e-11, 1.907986e-11, 
    1.909369e-11, 1.913266e-11, 1.906566e-11, 1.927304e-11, 1.914498e-11, 
    1.895368e-11, 1.899297e-11, 1.899859e-11, 1.898337e-11, 1.908665e-11, 
    1.904923e-11, 1.915e-11, 1.912277e-11, 1.916738e-11, 1.914522e-11, 
    1.914195e-11, 1.911348e-11, 1.909575e-11, 1.905095e-11, 1.901449e-11, 
    1.898558e-11, 1.89923e-11, 1.902406e-11, 1.908157e-11, 1.913596e-11, 
    1.912405e-11, 1.916399e-11, 1.905826e-11, 1.91026e-11, 1.908546e-11, 
    1.913015e-11, 1.903223e-11, 1.911559e-11, 1.901091e-11, 1.902009e-11, 
    1.904849e-11, 1.91056e-11, 1.911825e-11, 1.913173e-11, 1.912341e-11, 
    1.908303e-11, 1.907642e-11, 1.90478e-11, 1.90399e-11, 1.901809e-11, 
    1.900004e-11, 1.901653e-11, 1.903385e-11, 1.908305e-11, 1.912737e-11, 
    1.917568e-11, 1.918751e-11, 1.924391e-11, 1.919799e-11, 1.927376e-11, 
    1.920932e-11, 1.932086e-11, 1.912043e-11, 1.920744e-11, 1.904979e-11, 
    1.906678e-11, 1.90975e-11, 1.916797e-11, 1.912994e-11, 1.917441e-11, 
    1.907616e-11, 1.902515e-11, 1.901196e-11, 1.898733e-11, 1.901252e-11, 
    1.901048e-11, 1.903458e-11, 1.902683e-11, 1.908468e-11, 1.905361e-11, 
    1.914187e-11, 1.917407e-11, 1.926497e-11, 1.932067e-11, 1.937737e-11, 
    1.940239e-11, 1.941e-11, 1.941318e-11 ;

 SOIL2N_vr =
  1.818739, 1.81874, 1.81874, 1.818741, 1.81874, 1.818741, 1.818739, 1.81874, 
    1.818739, 1.818739, 1.818743, 1.818741, 1.818745, 1.818744, 1.818748, 
    1.818745, 1.818748, 1.818748, 1.818749, 1.818749, 1.818751, 1.818749, 
    1.818752, 1.81875, 1.818751, 1.818749, 1.818742, 1.818743, 1.818741, 
    1.818742, 1.818742, 1.81874, 1.81874, 1.818739, 1.818739, 1.81874, 
    1.818742, 1.818741, 1.818743, 1.818743, 1.818745, 1.818744, 1.818747, 
    1.818746, 1.818749, 1.818748, 1.818749, 1.818748, 1.818749, 1.818748, 
    1.818748, 1.818747, 1.818744, 1.818745, 1.818742, 1.81874, 1.818739, 
    1.818738, 1.818738, 1.818739, 1.81874, 1.818741, 1.818742, 1.818742, 
    1.818743, 1.818744, 1.818745, 1.818747, 1.818747, 1.818747, 1.818748, 
    1.818749, 1.818749, 1.818749, 1.818747, 1.818749, 1.818747, 1.818747, 
    1.818743, 1.818741, 1.81874, 1.81874, 1.818738, 1.818739, 1.818739, 
    1.81874, 1.818741, 1.81874, 1.818742, 1.818741, 1.818745, 1.818744, 
    1.818748, 1.818747, 1.818748, 1.818748, 1.818749, 1.818748, 1.818749, 
    1.81875, 1.818749, 1.818751, 1.818748, 1.818749, 1.81874, 1.81874, 
    1.818741, 1.81874, 1.81874, 1.818739, 1.818739, 1.81874, 1.818741, 
    1.818741, 1.818742, 1.818743, 1.818744, 1.818746, 1.818747, 1.818748, 
    1.818747, 1.818748, 1.818747, 1.818747, 1.81875, 1.818748, 1.81875, 
    1.81875, 1.818749, 1.81875, 1.81874, 1.81874, 1.818739, 1.81874, 
    1.818738, 1.818739, 1.81874, 1.818741, 1.818742, 1.818742, 1.818743, 
    1.818744, 1.818745, 1.818747, 1.818748, 1.818748, 1.818748, 1.818748, 
    1.818748, 1.818748, 1.818748, 1.818748, 1.81875, 1.81875, 1.81875, 
    1.81875, 1.81874, 1.818741, 1.81874, 1.818741, 1.818741, 1.818742, 
    1.818743, 1.818745, 1.818744, 1.818745, 1.818744, 1.818744, 1.818745, 
    1.818744, 1.818747, 1.818745, 1.818748, 1.818746, 1.818748, 1.818748, 
    1.818749, 1.818749, 1.81875, 1.818751, 1.818751, 1.818752, 1.818741, 
    1.818742, 1.818742, 1.818743, 1.818743, 1.818744, 1.818746, 1.818745, 
    1.818746, 1.818747, 1.818745, 1.818746, 1.818742, 1.818743, 1.818743, 
    1.818741, 1.818745, 1.818743, 1.818747, 1.818746, 1.818749, 1.818748, 
    1.818751, 1.818752, 1.818753, 1.818754, 1.818742, 1.818742, 1.818743, 
    1.818744, 1.818745, 1.818746, 1.818746, 1.818746, 1.818747, 1.818748, 
    1.818746, 1.818748, 1.818743, 1.818745, 1.818742, 1.818743, 1.818744, 
    1.818743, 1.818745, 1.818745, 1.818747, 1.818746, 1.818751, 1.818749, 
    1.818756, 1.818754, 1.818742, 1.818742, 1.818744, 1.818743, 1.818746, 
    1.818747, 1.818747, 1.818748, 1.818748, 1.818748, 1.818748, 1.818748, 
    1.818746, 1.818747, 1.818744, 1.818745, 1.818745, 1.818744, 1.818745, 
    1.818746, 1.818746, 1.818747, 1.818748, 1.818746, 1.818752, 1.818748, 
    1.818743, 1.818744, 1.818744, 1.818744, 1.818747, 1.818746, 1.818748, 
    1.818748, 1.818749, 1.818748, 1.818748, 1.818747, 1.818747, 1.818746, 
    1.818745, 1.818744, 1.818744, 1.818745, 1.818746, 1.818748, 1.818748, 
    1.818749, 1.818746, 1.818747, 1.818747, 1.818748, 1.818745, 1.818747, 
    1.818745, 1.818745, 1.818746, 1.818747, 1.818748, 1.818748, 1.818748, 
    1.818747, 1.818746, 1.818746, 1.818745, 1.818745, 1.818744, 1.818745, 
    1.818745, 1.818747, 1.818748, 1.818749, 1.818749, 1.818751, 1.81875, 
    1.818752, 1.81875, 1.818753, 1.818748, 1.81875, 1.818746, 1.818746, 
    1.818747, 1.818749, 1.818748, 1.818749, 1.818746, 1.818745, 1.818745, 
    1.818744, 1.818745, 1.818745, 1.818745, 1.818745, 1.818747, 1.818746, 
    1.818748, 1.818749, 1.818752, 1.818753, 1.818755, 1.818755, 1.818756, 
    1.818756,
  1.818756, 1.818758, 1.818758, 1.818759, 1.818758, 1.818759, 1.818757, 
    1.818758, 1.818757, 1.818756, 1.818761, 1.818759, 1.818764, 1.818762, 
    1.818766, 1.818763, 1.818766, 1.818766, 1.818767, 1.818767, 1.818769, 
    1.818768, 1.81877, 1.818769, 1.818769, 1.818768, 1.818759, 1.818761, 
    1.818759, 1.818759, 1.818759, 1.818758, 1.818758, 1.818756, 1.818756, 
    1.818757, 1.81876, 1.818759, 1.818761, 1.818761, 1.818763, 1.818762, 
    1.818765, 1.818764, 1.818767, 1.818766, 1.818767, 1.818767, 1.818767, 
    1.818766, 1.818766, 1.818765, 1.818762, 1.818763, 1.81876, 1.818758, 
    1.818757, 1.818756, 1.818756, 1.818756, 1.818757, 1.818759, 1.818759, 
    1.81876, 1.818761, 1.818762, 1.818763, 1.818765, 1.818765, 1.818766, 
    1.818766, 1.818767, 1.818767, 1.818767, 1.818766, 1.818767, 1.818765, 
    1.818765, 1.818761, 1.818759, 1.818758, 1.818758, 1.818756, 1.818757, 
    1.818757, 1.818758, 1.818758, 1.818758, 1.81876, 1.818759, 1.818763, 
    1.818762, 1.818766, 1.818765, 1.818766, 1.818766, 1.818767, 1.818766, 
    1.818768, 1.818768, 1.818768, 1.818769, 1.818766, 1.818767, 1.818758, 
    1.818758, 1.818758, 1.818757, 1.818757, 1.818756, 1.818757, 1.818758, 
    1.818758, 1.818759, 1.81876, 1.818761, 1.818762, 1.818764, 1.818765, 
    1.818766, 1.818765, 1.818766, 1.818765, 1.818765, 1.818768, 1.818766, 
    1.818769, 1.818769, 1.818767, 1.818769, 1.818758, 1.818758, 1.818757, 
    1.818758, 1.818756, 1.818757, 1.818757, 1.818759, 1.81876, 1.81876, 
    1.818761, 1.818762, 1.818763, 1.818765, 1.818766, 1.818766, 1.818766, 
    1.818766, 1.818766, 1.818767, 1.818767, 1.818766, 1.818769, 1.818768, 
    1.818769, 1.818768, 1.818758, 1.818758, 1.818758, 1.818759, 1.818758, 
    1.81876, 1.81876, 1.818763, 1.818762, 1.818763, 1.818762, 1.818762, 
    1.818763, 1.818762, 1.818765, 1.818763, 1.818766, 1.818765, 1.818767, 
    1.818766, 1.818767, 1.818767, 1.818768, 1.818769, 1.818769, 1.81877, 
    1.818759, 1.81876, 1.81876, 1.818761, 1.818761, 1.818762, 1.818764, 
    1.818763, 1.818764, 1.818765, 1.818763, 1.818764, 1.81876, 1.818761, 
    1.818761, 1.818759, 1.818763, 1.818761, 1.818765, 1.818764, 1.818767, 
    1.818766, 1.818769, 1.81877, 1.818772, 1.818773, 1.81876, 1.81876, 
    1.818761, 1.818762, 1.818763, 1.818764, 1.818764, 1.818764, 1.818765, 
    1.818766, 1.818765, 1.818766, 1.818761, 1.818763, 1.81876, 1.818761, 
    1.818762, 1.818761, 1.818763, 1.818764, 1.818765, 1.818764, 1.81877, 
    1.818768, 1.818774, 1.818772, 1.81876, 1.81876, 1.818762, 1.818761, 
    1.818764, 1.818765, 1.818765, 1.818766, 1.818766, 1.818767, 1.818766, 
    1.818767, 1.818764, 1.818765, 1.818762, 1.818763, 1.818762, 1.818762, 
    1.818763, 1.818765, 1.818765, 1.818765, 1.818766, 1.818764, 1.81877, 
    1.818766, 1.818761, 1.818762, 1.818762, 1.818762, 1.818765, 1.818764, 
    1.818767, 1.818766, 1.818767, 1.818766, 1.818766, 1.818766, 1.818765, 
    1.818764, 1.818763, 1.818762, 1.818762, 1.818763, 1.818765, 1.818766, 
    1.818766, 1.818767, 1.818764, 1.818765, 1.818765, 1.818766, 1.818763, 
    1.818766, 1.818763, 1.818763, 1.818764, 1.818765, 1.818766, 1.818766, 
    1.818766, 1.818765, 1.818764, 1.818764, 1.818763, 1.818763, 1.818762, 
    1.818763, 1.818763, 1.818765, 1.818766, 1.818767, 1.818768, 1.818769, 
    1.818768, 1.81877, 1.818768, 1.818772, 1.818766, 1.818768, 1.818764, 
    1.818764, 1.818765, 1.818767, 1.818766, 1.818767, 1.818764, 1.818763, 
    1.818763, 1.818762, 1.818763, 1.818763, 1.818763, 1.818763, 1.818765, 
    1.818764, 1.818766, 1.818767, 1.81877, 1.818772, 1.818773, 1.818774, 
    1.818774, 1.818774,
  1.818758, 1.81876, 1.818759, 1.818761, 1.81876, 1.818761, 1.818759, 
    1.81876, 1.818759, 1.818758, 1.818763, 1.818761, 1.818766, 1.818764, 
    1.818768, 1.818765, 1.818768, 1.818768, 1.818769, 1.818769, 1.818771, 
    1.81877, 1.818772, 1.818771, 1.818771, 1.81877, 1.818761, 1.818763, 
    1.818761, 1.818761, 1.818761, 1.81876, 1.818759, 1.818758, 1.818758, 
    1.818759, 1.818761, 1.818761, 1.818763, 1.818763, 1.818765, 1.818764, 
    1.818767, 1.818766, 1.818769, 1.818768, 1.818769, 1.818769, 1.818769, 
    1.818768, 1.818768, 1.818767, 1.818764, 1.818765, 1.818762, 1.81876, 
    1.818759, 1.818758, 1.818758, 1.818758, 1.818759, 1.818761, 1.818761, 
    1.818762, 1.818763, 1.818764, 1.818765, 1.818767, 1.818767, 1.818768, 
    1.818768, 1.818769, 1.818769, 1.81877, 1.818768, 1.818769, 1.818767, 
    1.818767, 1.818763, 1.818761, 1.81876, 1.81876, 1.818758, 1.818759, 
    1.818759, 1.81876, 1.81876, 1.81876, 1.818762, 1.818761, 1.818765, 
    1.818763, 1.818768, 1.818767, 1.818768, 1.818768, 1.818769, 1.818768, 
    1.81877, 1.81877, 1.81877, 1.818771, 1.818768, 1.818769, 1.81876, 
    1.81876, 1.81876, 1.818759, 1.818759, 1.818758, 1.818759, 1.818759, 
    1.81876, 1.818761, 1.818761, 1.818763, 1.818764, 1.818766, 1.818767, 
    1.818768, 1.818767, 1.818768, 1.818767, 1.818767, 1.81877, 1.818768, 
    1.818771, 1.818771, 1.81877, 1.818771, 1.81876, 1.81876, 1.818759, 
    1.81876, 1.818758, 1.818759, 1.818759, 1.818761, 1.818762, 1.818762, 
    1.818763, 1.818764, 1.818765, 1.818767, 1.818768, 1.818768, 1.818768, 
    1.818769, 1.818768, 1.818769, 1.818769, 1.818768, 1.818771, 1.81877, 
    1.818771, 1.81877, 1.81876, 1.81876, 1.81876, 1.818761, 1.81876, 
    1.818762, 1.818762, 1.818765, 1.818764, 1.818765, 1.818764, 1.818764, 
    1.818765, 1.818764, 1.818767, 1.818765, 1.818769, 1.818767, 1.818769, 
    1.818768, 1.818769, 1.818769, 1.81877, 1.818771, 1.818771, 1.818772, 
    1.818761, 1.818762, 1.818762, 1.818762, 1.818763, 1.818764, 1.818766, 
    1.818765, 1.818766, 1.818767, 1.818765, 1.818766, 1.818762, 1.818763, 
    1.818763, 1.818761, 1.818765, 1.818763, 1.818767, 1.818766, 1.818769, 
    1.818768, 1.818771, 1.818772, 1.818774, 1.818775, 1.818762, 1.818762, 
    1.818763, 1.818764, 1.818765, 1.818766, 1.818766, 1.818766, 1.818767, 
    1.818768, 1.818767, 1.818768, 1.818763, 1.818766, 1.818762, 1.818763, 
    1.818764, 1.818763, 1.818765, 1.818766, 1.818767, 1.818766, 1.818772, 
    1.81877, 1.818776, 1.818774, 1.818762, 1.818762, 1.818764, 1.818763, 
    1.818766, 1.818767, 1.818767, 1.818768, 1.818768, 1.818769, 1.818768, 
    1.818769, 1.818766, 1.818767, 1.818764, 1.818765, 1.818764, 1.818764, 
    1.818765, 1.818767, 1.818767, 1.818767, 1.818768, 1.818766, 1.818772, 
    1.818769, 1.818763, 1.818764, 1.818764, 1.818764, 1.818767, 1.818766, 
    1.818769, 1.818768, 1.818769, 1.818769, 1.818768, 1.818768, 1.818767, 
    1.818766, 1.818765, 1.818764, 1.818764, 1.818765, 1.818767, 1.818768, 
    1.818768, 1.818769, 1.818766, 1.818767, 1.818767, 1.818768, 1.818765, 
    1.818768, 1.818765, 1.818765, 1.818766, 1.818767, 1.818768, 1.818768, 
    1.818768, 1.818767, 1.818766, 1.818766, 1.818765, 1.818765, 1.818764, 
    1.818765, 1.818765, 1.818767, 1.818768, 1.818769, 1.81877, 1.818771, 
    1.81877, 1.818772, 1.81877, 1.818774, 1.818768, 1.81877, 1.818766, 
    1.818766, 1.818767, 1.818769, 1.818768, 1.818769, 1.818766, 1.818765, 
    1.818765, 1.818764, 1.818765, 1.818765, 1.818765, 1.818765, 1.818767, 
    1.818766, 1.818768, 1.818769, 1.818772, 1.818774, 1.818775, 1.818776, 
    1.818776, 1.818776,
  1.818741, 1.818742, 1.818742, 1.818743, 1.818742, 1.818743, 1.818741, 
    1.818742, 1.818741, 1.818741, 1.818745, 1.818743, 1.818748, 1.818746, 
    1.81875, 1.818748, 1.818751, 1.81875, 1.818752, 1.818751, 1.818753, 
    1.818752, 1.818755, 1.818753, 1.818753, 1.818752, 1.818744, 1.818745, 
    1.818743, 1.818744, 1.818744, 1.818742, 1.818742, 1.81874, 1.818741, 
    1.818742, 1.818744, 1.818743, 1.818745, 1.818745, 1.818747, 1.818746, 
    1.818749, 1.818748, 1.818751, 1.818751, 1.818751, 1.818751, 1.818751, 
    1.81875, 1.818751, 1.81875, 1.818746, 1.818747, 1.818744, 1.818742, 
    1.818741, 1.81874, 1.81874, 1.81874, 1.818742, 1.818743, 1.818744, 
    1.818744, 1.818745, 1.818747, 1.818748, 1.81875, 1.818749, 1.81875, 
    1.818751, 1.818751, 1.818751, 1.818752, 1.81875, 1.818751, 1.818749, 
    1.81875, 1.818745, 1.818743, 1.818743, 1.818742, 1.81874, 1.818741, 
    1.818741, 1.818742, 1.818743, 1.818742, 1.818744, 1.818744, 1.818748, 
    1.818746, 1.81875, 1.818749, 1.818751, 1.81875, 1.818751, 1.81875, 
    1.818752, 1.818752, 1.818752, 1.818753, 1.81875, 1.818751, 1.818742, 
    1.818742, 1.818743, 1.818742, 1.818742, 1.81874, 1.818741, 1.818742, 
    1.818743, 1.818743, 1.818744, 1.818745, 1.818746, 1.818748, 1.818749, 
    1.81875, 1.81875, 1.81875, 1.81875, 1.818749, 1.818752, 1.818751, 
    1.818753, 1.818753, 1.818752, 1.818753, 1.818742, 1.818742, 1.818741, 
    1.818742, 1.81874, 1.818741, 1.818742, 1.818744, 1.818744, 1.818744, 
    1.818745, 1.818746, 1.818748, 1.818749, 1.818751, 1.81875, 1.818751, 
    1.818751, 1.81875, 1.818751, 1.818751, 1.818751, 1.818753, 1.818752, 
    1.818753, 1.818752, 1.818742, 1.818743, 1.818743, 1.818743, 1.818743, 
    1.818744, 1.818745, 1.818747, 1.818746, 1.818748, 1.818746, 1.818746, 
    1.818748, 1.818746, 1.818749, 1.818747, 1.818751, 1.818749, 1.818751, 
    1.818751, 1.818751, 1.818752, 1.818752, 1.818754, 1.818753, 1.818754, 
    1.818743, 1.818744, 1.818744, 1.818745, 1.818745, 1.818746, 1.818748, 
    1.818748, 1.818749, 1.818749, 1.818747, 1.818748, 1.818745, 1.818745, 
    1.818745, 1.818744, 1.818748, 1.818745, 1.818749, 1.818748, 1.818752, 
    1.81875, 1.818753, 1.818755, 1.818756, 1.818757, 1.818745, 1.818744, 
    1.818745, 1.818746, 1.818747, 1.818748, 1.818748, 1.818749, 1.818749, 
    1.81875, 1.818749, 1.81875, 1.818745, 1.818748, 1.818744, 1.818745, 
    1.818746, 1.818745, 1.818747, 1.818748, 1.81875, 1.818749, 1.818754, 
    1.818752, 1.818759, 1.818757, 1.818744, 1.818745, 1.818747, 1.818746, 
    1.818748, 1.818749, 1.81875, 1.818751, 1.818751, 1.818751, 1.81875, 
    1.818751, 1.818748, 1.81875, 1.818746, 1.818747, 1.818747, 1.818746, 
    1.818748, 1.818749, 1.818749, 1.818749, 1.81875, 1.818748, 1.818755, 
    1.818751, 1.818745, 1.818746, 1.818746, 1.818746, 1.818749, 1.818748, 
    1.818751, 1.81875, 1.818751, 1.818751, 1.818751, 1.81875, 1.818749, 
    1.818748, 1.818747, 1.818746, 1.818746, 1.818747, 1.818749, 1.818751, 
    1.81875, 1.818751, 1.818748, 1.81875, 1.818749, 1.81875, 1.818748, 
    1.81875, 1.818747, 1.818747, 1.818748, 1.81875, 1.81875, 1.81875, 
    1.81875, 1.818749, 1.818749, 1.818748, 1.818748, 1.818747, 1.818747, 
    1.818747, 1.818748, 1.818749, 1.81875, 1.818752, 1.818752, 1.818754, 
    1.818752, 1.818755, 1.818753, 1.818756, 1.81875, 1.818753, 1.818748, 
    1.818748, 1.818749, 1.818751, 1.81875, 1.818752, 1.818749, 1.818747, 
    1.818747, 1.818746, 1.818747, 1.818747, 1.818748, 1.818747, 1.818749, 
    1.818748, 1.818751, 1.818752, 1.818754, 1.818756, 1.818758, 1.818758, 
    1.818759, 1.818759,
  1.81866, 1.818661, 1.818661, 1.818662, 1.818662, 1.818662, 1.81866, 
    1.818662, 1.818661, 1.81866, 1.818664, 1.818662, 1.818667, 1.818665, 
    1.818669, 1.818666, 1.818669, 1.818668, 1.81867, 1.81867, 1.818672, 
    1.81867, 1.818673, 1.818671, 1.818671, 1.81867, 1.818663, 1.818664, 
    1.818663, 1.818663, 1.818663, 1.818662, 1.818661, 1.81866, 1.81866, 
    1.818661, 1.818663, 1.818662, 1.818664, 1.818664, 1.818666, 1.818665, 
    1.818668, 1.818667, 1.81867, 1.818669, 1.81867, 1.818669, 1.81867, 
    1.818669, 1.818669, 1.818668, 1.818665, 1.818666, 1.818663, 1.818662, 
    1.81866, 1.81866, 1.81866, 1.81866, 1.818661, 1.818662, 1.818663, 
    1.818663, 1.818664, 1.818666, 1.818666, 1.818668, 1.818668, 1.818668, 
    1.818669, 1.81867, 1.81867, 1.81867, 1.818668, 1.818669, 1.818668, 
    1.818668, 1.818664, 1.818663, 1.818662, 1.818661, 1.81866, 1.818661, 
    1.81866, 1.818661, 1.818662, 1.818662, 1.818663, 1.818663, 1.818666, 
    1.818665, 1.818669, 1.818668, 1.818669, 1.818668, 1.81867, 1.818669, 
    1.81867, 1.818671, 1.81867, 1.818671, 1.818668, 1.81867, 1.818662, 
    1.818662, 1.818662, 1.818661, 1.818661, 1.81866, 1.818661, 1.818661, 
    1.818662, 1.818663, 1.818663, 1.818664, 1.818665, 1.818667, 1.818668, 
    1.818669, 1.818668, 1.818669, 1.818668, 1.818668, 1.81867, 1.818669, 
    1.818671, 1.818671, 1.81867, 1.818671, 1.818662, 1.818661, 1.81866, 
    1.818661, 1.81866, 1.818661, 1.818661, 1.818663, 1.818663, 1.818663, 
    1.818664, 1.818665, 1.818666, 1.818668, 1.818669, 1.818669, 1.818669, 
    1.818669, 1.818668, 1.818669, 1.818669, 1.818669, 1.818671, 1.81867, 
    1.818671, 1.818671, 1.818662, 1.818662, 1.818662, 1.818662, 1.818662, 
    1.818663, 1.818664, 1.818666, 1.818665, 1.818666, 1.818665, 1.818665, 
    1.818666, 1.818665, 1.818668, 1.818666, 1.818669, 1.818667, 1.818669, 
    1.818669, 1.818669, 1.81867, 1.818671, 1.818672, 1.818671, 1.818672, 
    1.818663, 1.818663, 1.818663, 1.818664, 1.818664, 1.818665, 1.818667, 
    1.818666, 1.818667, 1.818668, 1.818666, 1.818667, 1.818664, 1.818664, 
    1.818664, 1.818663, 1.818666, 1.818665, 1.818668, 1.818667, 1.81867, 
    1.818668, 1.818671, 1.818673, 1.818674, 1.818675, 1.818664, 1.818663, 
    1.818664, 1.818665, 1.818666, 1.818667, 1.818667, 1.818667, 1.818668, 
    1.818668, 1.818667, 1.818669, 1.818664, 1.818667, 1.818663, 1.818664, 
    1.818665, 1.818665, 1.818666, 1.818667, 1.818668, 1.818667, 1.818672, 
    1.81867, 1.818676, 1.818674, 1.818663, 1.818664, 1.818666, 1.818665, 
    1.818667, 1.818668, 1.818668, 1.818669, 1.818669, 1.818669, 1.818669, 
    1.818669, 1.818667, 1.818668, 1.818665, 1.818666, 1.818666, 1.818665, 
    1.818666, 1.818667, 1.818668, 1.818668, 1.818669, 1.818667, 1.818673, 
    1.818669, 1.818664, 1.818665, 1.818665, 1.818665, 1.818668, 1.818667, 
    1.818669, 1.818669, 1.81867, 1.818669, 1.818669, 1.818668, 1.818668, 
    1.818667, 1.818666, 1.818665, 1.818665, 1.818666, 1.818668, 1.818669, 
    1.818669, 1.81867, 1.818667, 1.818668, 1.818668, 1.818669, 1.818666, 
    1.818668, 1.818666, 1.818666, 1.818667, 1.818668, 1.818668, 1.818669, 
    1.818669, 1.818668, 1.818667, 1.818667, 1.818666, 1.818666, 1.818665, 
    1.818666, 1.818666, 1.818668, 1.818669, 1.81867, 1.81867, 1.818672, 
    1.818671, 1.818673, 1.818671, 1.818674, 1.818668, 1.818671, 1.818667, 
    1.818667, 1.818668, 1.81867, 1.818669, 1.81867, 1.818667, 1.818666, 
    1.818666, 1.818665, 1.818666, 1.818666, 1.818666, 1.818666, 1.818668, 
    1.818667, 1.818669, 1.81867, 1.818672, 1.818674, 1.818675, 1.818676, 
    1.818676, 1.818676,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2_HR_S1 =
  1.592376e-09, 1.596739e-09, 1.595891e-09, 1.599409e-09, 1.597458e-09, 
    1.599761e-09, 1.593261e-09, 1.596912e-09, 1.594582e-09, 1.59277e-09, 
    1.606232e-09, 1.599566e-09, 1.613157e-09, 1.608907e-09, 1.619583e-09, 
    1.612496e-09, 1.621011e-09, 1.619379e-09, 1.624293e-09, 1.622886e-09, 
    1.629168e-09, 1.624943e-09, 1.632426e-09, 1.62816e-09, 1.628827e-09, 
    1.624804e-09, 1.600908e-09, 1.605402e-09, 1.600642e-09, 1.601283e-09, 
    1.600995e-09, 1.597498e-09, 1.595735e-09, 1.592043e-09, 1.592714e-09, 
    1.595425e-09, 1.601571e-09, 1.599485e-09, 1.604742e-09, 1.604624e-09, 
    1.610474e-09, 1.607837e-09, 1.617667e-09, 1.614874e-09, 1.622944e-09, 
    1.620915e-09, 1.622849e-09, 1.622263e-09, 1.622857e-09, 1.61988e-09, 
    1.621155e-09, 1.618536e-09, 1.60833e-09, 1.61133e-09, 1.602381e-09, 
    1.596997e-09, 1.593421e-09, 1.590883e-09, 1.591242e-09, 1.591926e-09, 
    1.595441e-09, 1.598746e-09, 1.601264e-09, 1.602948e-09, 1.604607e-09, 
    1.609626e-09, 1.612284e-09, 1.618231e-09, 1.617159e-09, 1.618976e-09, 
    1.620713e-09, 1.623628e-09, 1.623149e-09, 1.624432e-09, 1.618929e-09, 
    1.622587e-09, 1.616548e-09, 1.618199e-09, 1.605055e-09, 1.600048e-09, 
    1.597917e-09, 1.596054e-09, 1.591518e-09, 1.59465e-09, 1.593415e-09, 
    1.596354e-09, 1.59822e-09, 1.597297e-09, 1.602994e-09, 1.600779e-09, 
    1.612441e-09, 1.607419e-09, 1.620511e-09, 1.617379e-09, 1.621261e-09, 
    1.61928e-09, 1.622674e-09, 1.61962e-09, 1.624911e-09, 1.626062e-09, 
    1.625275e-09, 1.628299e-09, 1.61945e-09, 1.622849e-09, 1.597271e-09, 
    1.597422e-09, 1.598123e-09, 1.595039e-09, 1.594851e-09, 1.592025e-09, 
    1.59454e-09, 1.59561e-09, 1.598328e-09, 1.599936e-09, 1.601464e-09, 
    1.604822e-09, 1.608573e-09, 1.613816e-09, 1.617582e-09, 1.620106e-09, 
    1.618558e-09, 1.619925e-09, 1.618397e-09, 1.617681e-09, 1.62563e-09, 
    1.621167e-09, 1.627864e-09, 1.627494e-09, 1.624463e-09, 1.627535e-09, 
    1.597527e-09, 1.596661e-09, 1.593652e-09, 1.596007e-09, 1.591717e-09, 
    1.594118e-09, 1.595499e-09, 1.600825e-09, 1.601996e-09, 1.60308e-09, 
    1.605223e-09, 1.607972e-09, 1.612793e-09, 1.616986e-09, 1.620814e-09, 
    1.620534e-09, 1.620633e-09, 1.621487e-09, 1.61937e-09, 1.621835e-09, 
    1.622249e-09, 1.621167e-09, 1.627444e-09, 1.625651e-09, 1.627486e-09, 
    1.626318e-09, 1.596943e-09, 1.598401e-09, 1.597613e-09, 1.599094e-09, 
    1.59805e-09, 1.60269e-09, 1.60408e-09, 1.610587e-09, 1.607917e-09, 
    1.612166e-09, 1.608349e-09, 1.609025e-09, 1.612304e-09, 1.608556e-09, 
    1.616755e-09, 1.611196e-09, 1.62152e-09, 1.61597e-09, 1.621868e-09, 
    1.620798e-09, 1.622571e-09, 1.624158e-09, 1.626155e-09, 1.629838e-09, 
    1.628986e-09, 1.632066e-09, 1.600574e-09, 1.602464e-09, 1.602298e-09, 
    1.604276e-09, 1.605738e-09, 1.608909e-09, 1.613992e-09, 1.612081e-09, 
    1.615589e-09, 1.616293e-09, 1.610963e-09, 1.614236e-09, 1.603729e-09, 
    1.605426e-09, 1.604416e-09, 1.600723e-09, 1.61252e-09, 1.606467e-09, 
    1.617644e-09, 1.614366e-09, 1.623931e-09, 1.619175e-09, 1.628516e-09, 
    1.632507e-09, 1.636264e-09, 1.640651e-09, 1.603496e-09, 1.602211e-09, 
    1.604511e-09, 1.607692e-09, 1.610643e-09, 1.614566e-09, 1.614967e-09, 
    1.615702e-09, 1.617605e-09, 1.619205e-09, 1.615934e-09, 1.619606e-09, 
    1.605819e-09, 1.613046e-09, 1.601726e-09, 1.605134e-09, 1.607504e-09, 
    1.606465e-09, 1.611862e-09, 1.613134e-09, 1.6183e-09, 1.61563e-09, 
    1.631521e-09, 1.624492e-09, 1.643991e-09, 1.638544e-09, 1.601763e-09, 
    1.603491e-09, 1.609506e-09, 1.606645e-09, 1.614828e-09, 1.616841e-09, 
    1.618478e-09, 1.62057e-09, 1.620796e-09, 1.622035e-09, 1.620004e-09, 
    1.621955e-09, 1.614574e-09, 1.617873e-09, 1.608819e-09, 1.611023e-09, 
    1.610009e-09, 1.608897e-09, 1.61233e-09, 1.615985e-09, 1.616064e-09, 
    1.617236e-09, 1.620536e-09, 1.614861e-09, 1.632427e-09, 1.62158e-09, 
    1.605376e-09, 1.608704e-09, 1.609181e-09, 1.607891e-09, 1.616639e-09, 
    1.61347e-09, 1.622005e-09, 1.619699e-09, 1.623477e-09, 1.6216e-09, 
    1.621324e-09, 1.618912e-09, 1.61741e-09, 1.613615e-09, 1.610527e-09, 
    1.608078e-09, 1.608648e-09, 1.611338e-09, 1.616209e-09, 1.620816e-09, 
    1.619807e-09, 1.62319e-09, 1.614235e-09, 1.61799e-09, 1.616539e-09, 
    1.620323e-09, 1.61203e-09, 1.61909e-09, 1.610224e-09, 1.611002e-09, 
    1.613407e-09, 1.618244e-09, 1.619315e-09, 1.620458e-09, 1.619753e-09, 
    1.616333e-09, 1.615773e-09, 1.613349e-09, 1.612679e-09, 1.610832e-09, 
    1.609303e-09, 1.6107e-09, 1.612167e-09, 1.616334e-09, 1.620088e-09, 
    1.62418e-09, 1.625182e-09, 1.629959e-09, 1.626069e-09, 1.632487e-09, 
    1.62703e-09, 1.636477e-09, 1.619501e-09, 1.62687e-09, 1.613517e-09, 
    1.614956e-09, 1.617558e-09, 1.623527e-09, 1.620306e-09, 1.624073e-09, 
    1.615751e-09, 1.61143e-09, 1.610313e-09, 1.608227e-09, 1.610361e-09, 
    1.610187e-09, 1.612229e-09, 1.611573e-09, 1.616473e-09, 1.613841e-09, 
    1.621316e-09, 1.624043e-09, 1.631743e-09, 1.636461e-09, 1.641263e-09, 
    1.643382e-09, 1.644027e-09, 1.644297e-09 ;

 SOIL2_HR_S3 =
  1.137412e-10, 1.140528e-10, 1.139922e-10, 1.142435e-10, 1.141041e-10, 
    1.142686e-10, 1.138044e-10, 1.140651e-10, 1.138987e-10, 1.137693e-10, 
    1.147309e-10, 1.142547e-10, 1.152255e-10, 1.14922e-10, 1.156845e-10, 
    1.151783e-10, 1.157865e-10, 1.156699e-10, 1.16021e-10, 1.159204e-10, 
    1.163692e-10, 1.160674e-10, 1.166018e-10, 1.162971e-10, 1.163448e-10, 
    1.160574e-10, 1.143506e-10, 1.146716e-10, 1.143316e-10, 1.143773e-10, 
    1.143568e-10, 1.14107e-10, 1.13981e-10, 1.137174e-10, 1.137653e-10, 
    1.139589e-10, 1.143979e-10, 1.14249e-10, 1.146245e-10, 1.14616e-10, 
    1.150339e-10, 1.148455e-10, 1.155476e-10, 1.153481e-10, 1.159246e-10, 
    1.157796e-10, 1.159178e-10, 1.158759e-10, 1.159183e-10, 1.157057e-10, 
    1.157968e-10, 1.156097e-10, 1.148807e-10, 1.15095e-10, 1.144558e-10, 
    1.140712e-10, 1.138158e-10, 1.136345e-10, 1.136601e-10, 1.13709e-10, 
    1.139601e-10, 1.141961e-10, 1.14376e-10, 1.144963e-10, 1.146148e-10, 
    1.149733e-10, 1.151631e-10, 1.155879e-10, 1.155113e-10, 1.156412e-10, 
    1.157652e-10, 1.159734e-10, 1.159392e-10, 1.160309e-10, 1.156378e-10, 
    1.15899e-10, 1.154677e-10, 1.155857e-10, 1.146468e-10, 1.142892e-10, 
    1.14137e-10, 1.140039e-10, 1.136798e-10, 1.139036e-10, 1.138154e-10, 
    1.140253e-10, 1.141586e-10, 1.140927e-10, 1.144995e-10, 1.143414e-10, 
    1.151744e-10, 1.148156e-10, 1.157507e-10, 1.155271e-10, 1.158044e-10, 
    1.156629e-10, 1.159053e-10, 1.156871e-10, 1.16065e-10, 1.161473e-10, 
    1.160911e-10, 1.163071e-10, 1.15675e-10, 1.159178e-10, 1.140908e-10, 
    1.141016e-10, 1.141517e-10, 1.139314e-10, 1.139179e-10, 1.137161e-10, 
    1.138957e-10, 1.139722e-10, 1.141663e-10, 1.142811e-10, 1.143903e-10, 
    1.146302e-10, 1.14898e-10, 1.152725e-10, 1.155416e-10, 1.157218e-10, 
    1.156113e-10, 1.157089e-10, 1.155998e-10, 1.155487e-10, 1.161165e-10, 
    1.157977e-10, 1.16276e-10, 1.162495e-10, 1.160331e-10, 1.162525e-10, 
    1.141091e-10, 1.140472e-10, 1.138323e-10, 1.140005e-10, 1.136941e-10, 
    1.138656e-10, 1.139642e-10, 1.143446e-10, 1.144283e-10, 1.145057e-10, 
    1.146588e-10, 1.148551e-10, 1.151995e-10, 1.15499e-10, 1.157724e-10, 
    1.157524e-10, 1.157595e-10, 1.158205e-10, 1.156693e-10, 1.158454e-10, 
    1.158749e-10, 1.157976e-10, 1.16246e-10, 1.161179e-10, 1.16249e-10, 
    1.161656e-10, 1.140673e-10, 1.141715e-10, 1.141152e-10, 1.14221e-10, 
    1.141465e-10, 1.144778e-10, 1.145772e-10, 1.150419e-10, 1.148512e-10, 
    1.151547e-10, 1.148821e-10, 1.149304e-10, 1.151645e-10, 1.148968e-10, 
    1.154825e-10, 1.150854e-10, 1.158229e-10, 1.154264e-10, 1.158477e-10, 
    1.157713e-10, 1.158979e-10, 1.160113e-10, 1.161539e-10, 1.16417e-10, 
    1.163561e-10, 1.165761e-10, 1.143267e-10, 1.144617e-10, 1.144498e-10, 
    1.145911e-10, 1.146956e-10, 1.149221e-10, 1.152851e-10, 1.151486e-10, 
    1.153992e-10, 1.154495e-10, 1.150688e-10, 1.153025e-10, 1.145521e-10, 
    1.146733e-10, 1.146011e-10, 1.143373e-10, 1.1518e-10, 1.147476e-10, 
    1.15546e-10, 1.153119e-10, 1.159951e-10, 1.156553e-10, 1.163226e-10, 
    1.166076e-10, 1.16876e-10, 1.171893e-10, 1.145354e-10, 1.144437e-10, 
    1.146079e-10, 1.148351e-10, 1.150459e-10, 1.153261e-10, 1.153548e-10, 
    1.154073e-10, 1.155432e-10, 1.156575e-10, 1.154238e-10, 1.156861e-10, 
    1.147014e-10, 1.152176e-10, 1.14409e-10, 1.146525e-10, 1.148217e-10, 
    1.147475e-10, 1.15133e-10, 1.152238e-10, 1.155928e-10, 1.154021e-10, 
    1.165372e-10, 1.160352e-10, 1.17428e-10, 1.170389e-10, 1.144116e-10, 
    1.145351e-10, 1.149647e-10, 1.147603e-10, 1.153448e-10, 1.154887e-10, 
    1.156056e-10, 1.15755e-10, 1.157711e-10, 1.158596e-10, 1.157146e-10, 
    1.158539e-10, 1.153267e-10, 1.155624e-10, 1.149157e-10, 1.150731e-10, 
    1.150007e-10, 1.149212e-10, 1.151664e-10, 1.154275e-10, 1.154331e-10, 
    1.155168e-10, 1.157526e-10, 1.153472e-10, 1.166019e-10, 1.158271e-10, 
    1.146697e-10, 1.149075e-10, 1.149415e-10, 1.148494e-10, 1.154742e-10, 
    1.152479e-10, 1.158575e-10, 1.156928e-10, 1.159627e-10, 1.158286e-10, 
    1.158088e-10, 1.156366e-10, 1.155293e-10, 1.152582e-10, 1.150377e-10, 
    1.148627e-10, 1.149034e-10, 1.150956e-10, 1.154435e-10, 1.157726e-10, 
    1.157005e-10, 1.159422e-10, 1.153025e-10, 1.155707e-10, 1.15467e-10, 
    1.157374e-10, 1.15145e-10, 1.156493e-10, 1.15016e-10, 1.150716e-10, 
    1.152434e-10, 1.155889e-10, 1.156654e-10, 1.15747e-10, 1.156966e-10, 
    1.154523e-10, 1.154123e-10, 1.152392e-10, 1.151914e-10, 1.150595e-10, 
    1.149502e-10, 1.1505e-10, 1.151548e-10, 1.154524e-10, 1.157206e-10, 
    1.160129e-10, 1.160844e-10, 1.164257e-10, 1.161478e-10, 1.166062e-10, 
    1.162164e-10, 1.168912e-10, 1.156786e-10, 1.16205e-10, 1.152512e-10, 
    1.15354e-10, 1.155399e-10, 1.159662e-10, 1.157361e-10, 1.160052e-10, 
    1.154108e-10, 1.151022e-10, 1.150224e-10, 1.148734e-10, 1.150258e-10, 
    1.150134e-10, 1.151592e-10, 1.151123e-10, 1.154623e-10, 1.152743e-10, 
    1.158083e-10, 1.160031e-10, 1.165531e-10, 1.168901e-10, 1.172331e-10, 
    1.173844e-10, 1.174305e-10, 1.174498e-10 ;

 SOIL3C =
  5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782616, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782616, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 
    5.782615, 5.782615, 5.782615, 5.782615, 5.782615, 5.782616, 5.782616, 
    5.782616, 5.782616 ;

 SOIL3C_TO_SOIL1C =
  3.139971e-11, 3.148571e-11, 3.1469e-11, 3.153834e-11, 3.149989e-11, 
    3.154528e-11, 3.141715e-11, 3.148912e-11, 3.144318e-11, 3.140746e-11, 
    3.167286e-11, 3.154144e-11, 3.180938e-11, 3.172559e-11, 3.193604e-11, 
    3.179634e-11, 3.196421e-11, 3.193203e-11, 3.202891e-11, 3.200116e-11, 
    3.212501e-11, 3.204171e-11, 3.218922e-11, 3.210513e-11, 3.211828e-11, 
    3.203897e-11, 3.15679e-11, 3.16565e-11, 3.156265e-11, 3.157529e-11, 
    3.156962e-11, 3.150067e-11, 3.146591e-11, 3.139315e-11, 3.140636e-11, 
    3.145981e-11, 3.158097e-11, 3.153986e-11, 3.164349e-11, 3.164115e-11, 
    3.175648e-11, 3.170449e-11, 3.189828e-11, 3.184321e-11, 3.200231e-11, 
    3.196231e-11, 3.200043e-11, 3.198887e-11, 3.200058e-11, 3.194191e-11, 
    3.196705e-11, 3.191541e-11, 3.171422e-11, 3.177336e-11, 3.159694e-11, 
    3.14908e-11, 3.142031e-11, 3.137027e-11, 3.137735e-11, 3.139083e-11, 
    3.146012e-11, 3.152527e-11, 3.157491e-11, 3.160811e-11, 3.164081e-11, 
    3.173976e-11, 3.179215e-11, 3.19094e-11, 3.188826e-11, 3.192408e-11, 
    3.195833e-11, 3.201579e-11, 3.200634e-11, 3.203165e-11, 3.192315e-11, 
    3.199526e-11, 3.187621e-11, 3.190877e-11, 3.164966e-11, 3.155095e-11, 
    3.150894e-11, 3.147221e-11, 3.138278e-11, 3.144454e-11, 3.14202e-11, 
    3.147812e-11, 3.151491e-11, 3.149672e-11, 3.160901e-11, 3.156536e-11, 
    3.179525e-11, 3.169625e-11, 3.195433e-11, 3.18926e-11, 3.196913e-11, 
    3.193008e-11, 3.199698e-11, 3.193677e-11, 3.204107e-11, 3.206377e-11, 
    3.204826e-11, 3.210786e-11, 3.193344e-11, 3.200043e-11, 3.14962e-11, 
    3.149917e-11, 3.1513e-11, 3.145221e-11, 3.144849e-11, 3.139278e-11, 
    3.144236e-11, 3.146346e-11, 3.151705e-11, 3.154873e-11, 3.157885e-11, 
    3.164507e-11, 3.1719e-11, 3.182235e-11, 3.18966e-11, 3.194635e-11, 
    3.191585e-11, 3.194278e-11, 3.191267e-11, 3.189856e-11, 3.205526e-11, 
    3.196728e-11, 3.209929e-11, 3.209199e-11, 3.203225e-11, 3.209281e-11, 
    3.150126e-11, 3.148418e-11, 3.142487e-11, 3.147128e-11, 3.138671e-11, 
    3.143405e-11, 3.146126e-11, 3.156626e-11, 3.158934e-11, 3.161072e-11, 
    3.165295e-11, 3.170714e-11, 3.180219e-11, 3.188486e-11, 3.196032e-11, 
    3.195479e-11, 3.195674e-11, 3.197359e-11, 3.193184e-11, 3.198044e-11, 
    3.19886e-11, 3.196727e-11, 3.209101e-11, 3.205567e-11, 3.209184e-11, 
    3.206882e-11, 3.148973e-11, 3.151847e-11, 3.150294e-11, 3.153214e-11, 
    3.151156e-11, 3.160302e-11, 3.163044e-11, 3.17587e-11, 3.170608e-11, 
    3.178983e-11, 3.171459e-11, 3.172792e-11, 3.179255e-11, 3.171866e-11, 
    3.188029e-11, 3.17707e-11, 3.197424e-11, 3.186482e-11, 3.19811e-11, 
    3.195999e-11, 3.199494e-11, 3.202623e-11, 3.20656e-11, 3.213822e-11, 
    3.21214e-11, 3.218213e-11, 3.156131e-11, 3.159857e-11, 3.15953e-11, 
    3.163429e-11, 3.166312e-11, 3.172562e-11, 3.182582e-11, 3.178815e-11, 
    3.185732e-11, 3.18712e-11, 3.176612e-11, 3.183063e-11, 3.162351e-11, 
    3.165697e-11, 3.163705e-11, 3.156424e-11, 3.179682e-11, 3.167748e-11, 
    3.189782e-11, 3.18332e-11, 3.202177e-11, 3.192799e-11, 3.211215e-11, 
    3.219082e-11, 3.226488e-11, 3.235136e-11, 3.161891e-11, 3.159359e-11, 
    3.163893e-11, 3.170162e-11, 3.175981e-11, 3.183714e-11, 3.184506e-11, 
    3.185954e-11, 3.189705e-11, 3.192859e-11, 3.186411e-11, 3.19365e-11, 
    3.166472e-11, 3.180718e-11, 3.158402e-11, 3.165122e-11, 3.169794e-11, 
    3.167745e-11, 3.178385e-11, 3.180891e-11, 3.191075e-11, 3.185812e-11, 
    3.217139e-11, 3.203283e-11, 3.241722e-11, 3.230984e-11, 3.158475e-11, 
    3.161883e-11, 3.17374e-11, 3.168099e-11, 3.184231e-11, 3.1882e-11, 
    3.191427e-11, 3.19555e-11, 3.195996e-11, 3.198439e-11, 3.194435e-11, 
    3.198281e-11, 3.183731e-11, 3.190233e-11, 3.172386e-11, 3.17673e-11, 
    3.174732e-11, 3.172539e-11, 3.179306e-11, 3.186512e-11, 3.186668e-11, 
    3.188978e-11, 3.195483e-11, 3.184296e-11, 3.218924e-11, 3.197541e-11, 
    3.165598e-11, 3.172159e-11, 3.173098e-11, 3.170557e-11, 3.187802e-11, 
    3.181554e-11, 3.198379e-11, 3.193833e-11, 3.201282e-11, 3.197581e-11, 
    3.197036e-11, 3.192282e-11, 3.189321e-11, 3.181841e-11, 3.175753e-11, 
    3.170925e-11, 3.172048e-11, 3.177351e-11, 3.186953e-11, 3.196035e-11, 
    3.194046e-11, 3.200716e-11, 3.183061e-11, 3.190465e-11, 3.187603e-11, 
    3.195064e-11, 3.178715e-11, 3.192634e-11, 3.175155e-11, 3.176688e-11, 
    3.18143e-11, 3.190966e-11, 3.193077e-11, 3.195329e-11, 3.19394e-11, 
    3.187197e-11, 3.186093e-11, 3.181315e-11, 3.179995e-11, 3.176355e-11, 
    3.173339e-11, 3.176094e-11, 3.178986e-11, 3.187201e-11, 3.194601e-11, 
    3.202667e-11, 3.204642e-11, 3.21406e-11, 3.206392e-11, 3.219043e-11, 
    3.208285e-11, 3.226908e-11, 3.193442e-11, 3.20797e-11, 3.181646e-11, 
    3.184484e-11, 3.189614e-11, 3.201379e-11, 3.195029e-11, 3.202456e-11, 
    3.18605e-11, 3.177533e-11, 3.17533e-11, 3.171218e-11, 3.175425e-11, 
    3.175083e-11, 3.179107e-11, 3.177814e-11, 3.187473e-11, 3.182285e-11, 
    3.197022e-11, 3.202398e-11, 3.217576e-11, 3.226876e-11, 3.236343e-11, 
    3.240521e-11, 3.241792e-11, 3.242324e-11 ;

 SOIL3C_vr =
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 20.00008, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00009, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 20.00008, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 
    20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00009, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00009, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00009, 20.00008, 
    20.00008, 20.00008, 20.00009, 20.00008, 20.00009, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009,
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00009, 20.00008, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 
    20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00008, 20.00009, 20.00008, 20.00008, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009,
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00009, 20.00008, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00008, 20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00009, 20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00008, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 20.00009, 
    20.00009, 20.00009,
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00008, 20.00008, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00008, 20.00008, 
    20.00008, 20.00008,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N =
  0.5256922, 0.5256923, 0.5256922, 0.5256923, 0.5256923, 0.5256923, 
    0.5256922, 0.5256923, 0.5256922, 0.5256922, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256922, 0.5256922, 0.5256922, 0.5256922, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256922, 0.5256922, 0.5256922, 0.5256922, 
    0.5256922, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256922, 0.5256922, 0.5256922, 
    0.5256922, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256922, 
    0.5256922, 0.5256922, 0.5256922, 0.5256922, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256922, 0.5256922, 0.5256922, 0.5256922, 0.5256922, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 0.5256923, 
    0.5256923, 0.5256923 ;

 SOIL3N_TNDNCY_VERT_TRANS =
  1.027984e-20, 2.569961e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, 
    -2.569961e-21, 7.709882e-21, -5.139921e-21, -2.569961e-21, 7.709882e-21, 
    7.709882e-21, -1.798972e-20, -2.055969e-20, 0, -7.709882e-21, 
    -2.826957e-20, -2.569961e-21, -2.826957e-20, 5.139921e-21, 1.28498e-20, 
    -2.569961e-21, -5.139921e-21, -7.709882e-21, 1.027984e-20, -5.139921e-21, 
    -1.027984e-20, 1.28498e-20, 0, -2.569961e-21, -7.709882e-21, 
    5.139921e-21, 5.139921e-21, 1.003089e-36, -1.28498e-20, -7.709882e-21, 
    1.541976e-20, -1.798972e-20, -5.139921e-21, -2.569961e-21, 7.709882e-21, 
    -2.569961e-21, -1.798972e-20, 1.798972e-20, -2.569961e-21, -1.541976e-20, 
    -1.003089e-36, 7.709882e-21, 5.139921e-21, -2.055969e-20, -7.709882e-21, 
    -1.798972e-20, -5.139921e-21, 2.569961e-21, -2.569961e-21, -2.569961e-21, 
    7.709882e-21, 0, 2.569961e-21, -1.28498e-20, -5.139921e-21, 
    -7.709882e-21, 0, 7.709882e-21, -1.28498e-20, -1.003089e-36, 
    -1.28498e-20, 2.569961e-21, 2.569961e-21, 2.055969e-20, -1.798972e-20, 
    -7.709882e-21, -5.139921e-21, 1.003089e-36, 1.027984e-20, 2.312965e-20, 
    -5.139921e-21, -2.569961e-20, -5.139921e-21, -2.569961e-21, 1.28498e-20, 
    5.139921e-21, 5.139921e-21, -2.569961e-21, 2.569961e-21, -7.709882e-21, 
    2.569961e-21, 1.027984e-20, -2.569961e-21, 5.139921e-21, 2.569961e-21, 
    -2.569961e-20, 5.139921e-21, 5.139921e-21, 5.139921e-21, 1.28498e-20, 
    2.569961e-21, 2.569961e-21, -1.798972e-20, -2.569961e-21, -1.003089e-36, 
    -7.709882e-21, 2.569961e-21, 7.709882e-21, -1.541976e-20, -5.139921e-21, 
    1.003089e-36, -2.569961e-21, 1.541976e-20, -2.569961e-21, 0, 
    -1.28498e-20, 1.027984e-20, -2.569961e-21, -5.139921e-21, 7.709882e-21, 
    -1.28498e-20, -2.312965e-20, 1.541976e-20, -1.798972e-20, 5.139921e-21, 
    5.139921e-21, -5.139921e-21, 0, -1.027984e-20, -2.569961e-21, 
    7.709882e-21, 1.541976e-20, -5.139921e-21, -1.003089e-36, -1.541976e-20, 
    5.139921e-21, -7.709882e-21, -1.28498e-20, -7.709882e-21, 5.139921e-21, 
    -1.28498e-20, -2.569961e-21, -5.139921e-21, 2.569961e-21, -2.569961e-21, 
    5.139921e-21, -2.569961e-21, -2.569961e-21, -5.139921e-21, -1.027984e-20, 
    7.709882e-21, 7.709882e-21, -2.055969e-20, 2.569961e-21, -7.709882e-21, 
    -5.139921e-21, 0, 1.541976e-20, -1.28498e-20, 5.139921e-21, 
    -5.139921e-21, 2.569961e-21, -5.139921e-21, 1.003089e-36, 1.027984e-20, 
    -2.569961e-21, 2.569961e-21, 2.569961e-21, 0, -2.569961e-21, 
    5.139921e-21, -5.139921e-21, 0, 2.569961e-21, -5.139921e-21, 
    1.541976e-20, 2.569961e-21, -1.027984e-20, -7.709882e-21, -2.055969e-20, 
    2.569961e-21, 1.28498e-20, -7.709882e-21, -2.569961e-21, 2.569961e-21, 
    2.569961e-21, -2.569961e-21, -2.569961e-21, -1.003089e-36, -5.139921e-21, 
    -1.027984e-20, -5.139921e-21, -1.541976e-20, 7.709882e-21, 5.139921e-21, 
    5.139921e-21, 1.027984e-20, 1.003089e-36, -1.027984e-20, -5.139921e-21, 
    2.569961e-21, -5.139921e-21, 5.139921e-21, -1.003089e-36, -2.055969e-20, 
    7.709882e-21, -1.28498e-20, 0, 2.569961e-21, -7.709882e-21, 2.569961e-21, 
    -1.027984e-20, -7.709882e-21, -2.569961e-21, -1.28498e-20, -1.027984e-20, 
    -5.139921e-21, 1.541976e-20, -2.569961e-21, -1.541976e-20, -7.709882e-21, 
    5.139921e-21, -1.541976e-20, -5.139921e-21, -2.569961e-21, 2.569961e-21, 
    -2.569961e-20, 1.027984e-20, 1.28498e-20, 5.139921e-21, -2.569961e-21, 
    -2.569961e-21, 5.139921e-21, -5.139921e-21, 2.569961e-21, -2.569961e-21, 
    -2.569961e-21, -1.003089e-36, 0, -1.027984e-20, 5.139921e-21, 
    1.027984e-20, 5.139921e-21, -1.541976e-20, 1.003089e-36, -5.139921e-21, 
    -1.541976e-20, -7.709882e-21, 5.139921e-21, -2.569961e-21, -5.139921e-21, 
    1.28498e-20, 1.027984e-20, 1.027984e-20, -1.798972e-20, 1.027984e-20, 
    -5.139921e-21, -1.027984e-20, 1.798972e-20, 7.709882e-21, 1.28498e-20, 
    1.027984e-20, 7.709882e-21, -1.541976e-20, -5.139921e-21, 5.139921e-21, 
    1.541976e-20, -2.569961e-21, -2.569961e-21, 0, -2.569961e-21, 
    7.709882e-21, 0, 2.826957e-20, 5.139921e-21, 7.709882e-21, 2.569961e-21, 
    -2.569961e-21, 1.003089e-36, -2.569961e-21, 5.139921e-21, 2.569961e-21, 
    -5.139921e-21, -7.709882e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, 
    2.569961e-21, -2.569961e-21, -1.541976e-20, -1.003089e-36, -2.569961e-21, 
    7.709882e-21, -7.709882e-21, -5.139921e-21, 0, -2.569961e-21, 
    -2.569961e-21, 1.798972e-20, 1.027984e-20, -1.027984e-20, 2.569961e-21, 
    -2.569961e-21, -1.541976e-20, -5.139921e-21, -5.139921e-21, 2.569961e-21, 
    -2.569961e-21, 1.027984e-20, 1.003089e-36, -2.569961e-21, 1.798972e-20, 
    -7.709882e-21, 1.027984e-20, 1.798972e-20, -1.28498e-20, 1.28498e-20, 
    -2.569961e-21, -7.709882e-21, 5.139921e-21, -1.027984e-20, -2.569961e-21, 
    1.798972e-20, 2.569961e-21, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    2.569961e-21, 5.139921e-21, -1.28498e-20, -7.709882e-21, 2.569961e-21, 
    -7.709882e-21, 5.139921e-21, 7.709882e-21, 1.027984e-20, 1.28498e-20, 
    1.027984e-20, -2.569961e-21, -1.003089e-36, 7.709882e-21, -1.003089e-36, 
    5.139921e-21,
  0, 1.541976e-20, 0, -1.027984e-20, -5.139921e-21, 5.139921e-21, 
    -1.541976e-20, 2.569961e-21, 0, 2.569961e-21, 1.28498e-20, -2.569961e-21, 
    -1.027984e-20, 1.027984e-20, -2.569961e-21, -7.709882e-21, 2.569961e-21, 
    5.139921e-21, -2.569961e-21, -1.027984e-20, 2.569961e-21, 5.139921e-21, 
    -5.139921e-21, -7.709882e-21, -2.569961e-21, 1.798972e-20, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, -1.798972e-20, -1.027984e-20, 1.798972e-20, 
    7.709882e-21, 7.709882e-21, -2.569961e-21, -2.569961e-21, 7.709882e-21, 
    2.569961e-21, -5.139921e-21, 5.139921e-21, 2.569961e-21, -2.569961e-21, 
    7.709882e-21, -1.003089e-36, -2.569961e-21, -5.139921e-21, 0, 0, 0, 
    -2.569961e-21, -1.003089e-36, -2.569961e-21, 0, -1.027984e-20, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, 5.139921e-21, -5.139921e-21, 
    -2.569961e-21, -7.709882e-21, -2.569961e-21, -5.139921e-21, 
    -5.139921e-21, -2.569961e-21, -7.709882e-21, 7.709882e-21, 1.28498e-20, 
    2.569961e-21, 1.027984e-20, -5.139921e-21, -1.003089e-36, -7.709882e-21, 
    -1.28498e-20, 0, -2.569961e-21, -5.139921e-21, 0, -7.709882e-21, 
    7.709882e-21, 2.569961e-21, -2.569961e-21, 1.798972e-20, 2.055969e-20, 
    -2.569961e-21, 2.569961e-21, 0, -5.139921e-21, -7.709882e-21, 
    -2.569961e-21, 7.709882e-21, -7.709882e-21, -1.28498e-20, 1.28498e-20, 
    2.569961e-21, 2.569961e-21, 5.139921e-21, 5.139921e-21, -2.569961e-21, 
    2.569961e-21, 1.541976e-20, 7.709882e-21, -5.139921e-21, 0, 
    -1.798972e-20, 1.541976e-20, 2.569961e-21, 7.709882e-21, -2.569961e-21, 
    -2.569961e-21, -7.709882e-21, -1.28498e-20, 5.139921e-21, -2.569961e-21, 
    1.027984e-20, -2.569961e-21, -2.569961e-21, 7.709882e-21, -5.139921e-21, 
    5.139921e-21, 7.709882e-21, 2.569961e-21, -1.003089e-36, 5.139921e-21, 0, 
    7.709882e-21, 7.709882e-21, 7.709882e-21, 2.569961e-21, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, 1.003089e-36, -1.027984e-20, -2.569961e-21, 
    -1.28498e-20, 2.569961e-21, 2.569961e-21, 1.027984e-20, -2.569961e-21, 
    5.139921e-21, -1.027984e-20, -7.709882e-21, 2.569961e-21, 5.139921e-21, 
    1.027984e-20, 5.139921e-21, 2.569961e-21, -1.541976e-20, -5.139921e-21, 
    -1.541976e-20, 0, 1.027984e-20, 5.139921e-21, 2.569961e-21, 
    -2.569961e-21, -2.569961e-21, 1.027984e-20, 1.28498e-20, 7.709882e-21, 
    -5.139921e-21, 2.569961e-21, -1.28498e-20, 0, 1.798972e-20, 
    -1.541976e-20, -7.709882e-21, -5.139921e-21, 2.569961e-21, -7.709882e-21, 
    -1.003089e-36, 5.139921e-21, 7.709882e-21, 5.139921e-21, 1.027984e-20, 
    -2.569961e-21, -5.139921e-21, 1.027984e-20, 7.709882e-21, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -7.709882e-21, 0, -2.569961e-21, 
    -2.569961e-21, 2.055969e-20, -5.139921e-21, -2.569961e-21, 1.28498e-20, 
    2.569961e-21, -1.003089e-36, 2.569961e-21, -5.139921e-21, 7.709882e-21, 
    -5.139921e-21, -2.569961e-21, 0, 2.569961e-21, -1.541976e-20, 
    2.569961e-21, 2.569961e-21, -5.139921e-21, 2.569961e-21, 1.027984e-20, 
    -5.139921e-21, -7.709882e-21, 2.569961e-21, -1.28498e-20, 5.139921e-21, 
    -1.027984e-20, -1.798972e-20, 2.569961e-21, 0, 0, 7.709882e-21, 
    5.139921e-21, 2.569961e-21, -1.027984e-20, 7.709882e-21, -7.709882e-21, 
    5.139921e-21, -5.139921e-21, 5.139921e-21, -5.139921e-21, -2.569961e-21, 
    -2.569961e-21, 0, -2.569961e-21, 1.003089e-36, 5.139921e-21, 1.28498e-20, 
    -7.709882e-21, -1.003089e-36, 0, -5.139921e-21, 2.569961e-21, 
    7.709882e-21, -2.569961e-21, -1.003089e-36, 2.569961e-21, -7.709882e-21, 
    1.027984e-20, 5.139921e-21, -1.027984e-20, -2.569961e-21, -2.569961e-21, 
    1.541976e-20, -7.709882e-21, 0, -1.541976e-20, 0, 7.709882e-21, 
    -1.541976e-20, -1.28498e-20, 7.709882e-21, -2.569961e-21, -1.027984e-20, 
    7.709882e-21, 2.569961e-21, -7.709882e-21, -7.709882e-21, -5.139921e-21, 
    0, 1.003089e-36, -1.027984e-20, 1.027984e-20, 5.139921e-21, 7.709882e-21, 
    -2.569961e-21, 7.709882e-21, 2.569961e-21, -1.28498e-20, -7.709882e-21, 
    7.709882e-21, -2.569961e-21, 5.139921e-21, -7.709882e-21, 2.569961e-21, 
    -1.027984e-20, -5.139921e-21, 1.027984e-20, -1.28498e-20, 0, 
    -5.139921e-21, -1.027984e-20, 1.28498e-20, -1.541976e-20, -5.139921e-21, 
    -2.569961e-21, -7.709882e-21, 7.709882e-21, -7.709882e-21, 2.569961e-21, 
    -7.709882e-21, 5.139921e-21, -2.569961e-21, 1.027984e-20, -2.569961e-21, 
    1.003089e-36, 1.027984e-20, 1.28498e-20, 7.709882e-21, 7.709882e-21, 
    -5.139921e-21, -2.569961e-21, -1.003089e-36, 1.28498e-20, -1.027984e-20, 
    1.003089e-36, -1.28498e-20, -7.709882e-21, 5.139921e-21, -2.569961e-21, 
    -2.569961e-21, 1.027984e-20, 1.28498e-20, 2.569961e-21, 1.28498e-20, 
    1.027984e-20, 7.709882e-21, 7.709882e-21, 0, 5.139921e-21, 0, 
    5.139921e-21, 1.541976e-20, 7.709882e-21, -5.139921e-21, 2.569961e-21, 
    -5.139921e-21, -1.027984e-20, 2.569961e-21, 5.139921e-21, 1.027984e-20, 
    1.28498e-20, -2.569961e-21, 1.027984e-20,
  0, -1.28498e-20, 7.709882e-21, 2.055969e-20, -1.027984e-20, -1.027984e-20, 
    2.569961e-21, 1.003089e-36, -1.027984e-20, -2.569961e-21, 0, 
    1.027984e-20, -5.139921e-21, -7.709882e-21, -7.709882e-21, -7.709882e-21, 
    -1.027984e-20, -5.139921e-21, -5.139921e-21, -7.709882e-21, 
    -7.709882e-21, 0, -7.709882e-21, 2.569961e-21, -1.027984e-20, 
    -1.003089e-36, -5.139921e-21, -1.027984e-20, 7.709882e-21, 1.003089e-36, 
    -1.027984e-20, 5.139921e-21, -1.003089e-36, -1.003089e-36, 7.709882e-21, 
    -1.003089e-36, -5.139921e-21, 5.139921e-21, -2.569961e-21, -1.541976e-20, 
    -1.027984e-20, -1.28498e-20, 2.569961e-21, -7.709882e-21, -2.569961e-21, 
    0, 7.709882e-21, -5.139921e-21, -5.139921e-21, -2.569961e-21, 
    -2.312965e-20, 1.003089e-36, 7.709882e-21, 7.709882e-21, 0, 
    -5.139921e-21, 1.28498e-20, -5.139921e-21, -1.28498e-20, 1.027984e-20, 
    2.569961e-21, 2.569961e-21, -5.139921e-21, -7.709882e-21, -2.569961e-21, 
    -5.139921e-21, 7.709882e-21, -1.28498e-20, -2.569961e-21, -1.003089e-36, 
    2.569961e-21, 1.28498e-20, 2.569961e-21, -7.709882e-21, 1.027984e-20, 
    2.569961e-21, -5.139921e-21, -7.709882e-21, 2.569961e-21, -7.709882e-21, 
    1.541976e-20, 2.569961e-21, -1.28498e-20, 0, 1.027984e-20, -5.139921e-21, 
    0, -2.569961e-21, 2.569961e-21, -2.569961e-21, 5.139921e-21, 
    -1.003089e-36, 2.569961e-21, -7.709882e-21, 7.709882e-21, -5.139921e-21, 
    5.139921e-21, 0, 0, 7.709882e-21, 0, -2.569961e-21, -7.709882e-21, 
    1.027984e-20, 1.28498e-20, -7.709882e-21, 1.28498e-20, -1.003089e-36, 0, 
    1.027984e-20, -2.569961e-21, -2.055969e-20, -2.569961e-21, 0, 
    2.569961e-21, 1.003089e-36, -2.569961e-21, -2.569961e-21, -5.139921e-21, 
    2.569961e-21, 2.569961e-21, -2.569961e-21, 2.569961e-21, 5.139921e-21, 0, 
    5.139921e-21, -2.569961e-21, 1.027984e-20, 2.569961e-21, -5.139921e-21, 
    -5.139921e-21, 2.569961e-21, -1.027984e-20, 0, -7.709882e-21, 
    -1.027984e-20, -1.027984e-20, 5.139921e-21, -2.569961e-21, -5.139921e-21, 
    2.569961e-21, -1.027984e-20, 1.003089e-36, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, 2.569961e-21, 2.569961e-21, -1.541976e-20, 1.28498e-20, 
    -7.709882e-21, -1.28498e-20, -5.139921e-21, -5.139921e-21, 1.541976e-20, 
    -7.709882e-21, 2.569961e-21, -1.003089e-36, -5.139921e-21, 1.027984e-20, 
    0, 1.28498e-20, 5.139921e-21, -5.139921e-21, -1.541976e-20, 
    -5.139921e-21, 5.139921e-21, 0, -5.139921e-21, 5.139921e-21, 
    -5.139921e-21, 7.709882e-21, 5.139921e-21, 7.709882e-21, 2.569961e-21, 
    -1.027984e-20, 5.139921e-21, -5.139921e-21, 1.027984e-20, 1.003089e-36, 
    1.027984e-20, 5.139921e-21, -5.139921e-21, -2.569961e-21, 1.541976e-20, 
    1.027984e-20, -5.139921e-21, 1.027984e-20, -1.027984e-20, 7.709882e-21, 
    -5.139921e-21, 0, -7.709882e-21, 2.569961e-21, -1.003089e-36, 
    5.139921e-21, 0, -5.139921e-21, -2.312965e-20, 1.28498e-20, 
    -1.027984e-20, -2.569961e-21, 1.027984e-20, -5.139921e-21, -1.003089e-36, 
    7.709882e-21, -7.709882e-21, 1.027984e-20, -2.569961e-21, 1.541976e-20, 
    2.569961e-21, 5.139921e-21, 7.709882e-21, -1.027984e-20, 5.139921e-21, 
    1.541976e-20, -1.027984e-20, 2.569961e-21, -2.569961e-21, 2.569961e-21, 
    -2.569961e-21, -7.709882e-21, 1.003089e-36, -5.139921e-21, -5.139921e-21, 
    1.003089e-36, 5.139921e-21, -1.003089e-36, -1.798972e-20, 7.709882e-21, 
    0, 7.709882e-21, 1.027984e-20, 7.709882e-21, 2.569961e-21, 0, 
    1.798972e-20, 1.28498e-20, 5.139921e-21, -1.28498e-20, 1.28498e-20, 
    -1.027984e-20, -1.027984e-20, -5.139921e-21, 5.139921e-21, -1.541976e-20, 
    2.569961e-21, -5.139921e-21, -1.027984e-20, 1.798972e-20, 1.541976e-20, 
    1.027984e-20, 1.28498e-20, -2.569961e-21, -1.027984e-20, 0, 0, 
    -1.027984e-20, 1.003089e-36, -1.28498e-20, -2.569961e-21, 0, 0, 
    2.569961e-21, 0, 7.709882e-21, -2.569961e-21, 1.027984e-20, 
    -2.569961e-21, -7.709882e-21, 7.709882e-21, -5.139921e-21, -5.139921e-21, 
    1.027984e-20, 7.709882e-21, 0, 2.569961e-21, 7.709882e-21, 7.709882e-21, 
    -2.055969e-20, -2.569961e-21, 0, -7.709882e-21, -2.569961e-21, 
    1.798972e-20, -1.027984e-20, -1.003089e-36, 2.569961e-21, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, 7.709882e-21, 0, 2.055969e-20, 1.027984e-20, 
    5.139921e-21, -2.569961e-21, -2.569961e-21, 2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, 5.139921e-21, 
    7.709882e-21, -7.709882e-21, -1.027984e-20, 2.569961e-21, 1.541976e-20, 
    1.003089e-36, 1.027984e-20, 1.541976e-20, 1.027984e-20, -7.709882e-21, 
    -1.28498e-20, 5.139921e-21, 2.569961e-21, 5.139921e-21, -5.139921e-21, 
    1.027984e-20, 5.139921e-21, -1.027984e-20, 5.139921e-21, 2.055969e-20, 
    -1.798972e-20, 1.541976e-20, 1.798972e-20, 2.569961e-21, 2.569961e-21, 
    1.003089e-36, 7.709882e-21, -2.569961e-21, -2.569961e-21, -1.003089e-36, 
    2.569961e-21, -7.709882e-21, 5.139921e-21,
  2.569961e-21, 2.569961e-21, -1.003089e-36, 2.569961e-21, 1.027984e-20, 
    1.027984e-20, -1.28498e-20, -1.541976e-20, 1.027984e-20, -1.003089e-36, 
    -5.139921e-21, -1.541976e-20, -2.569961e-21, -1.027984e-20, 2.569961e-21, 
    -1.027984e-20, 7.709882e-21, 1.28498e-20, 7.709882e-21, 2.055969e-20, 
    1.003089e-36, 1.798972e-20, 5.139921e-21, 1.003089e-36, 1.28498e-20, 
    -2.569961e-21, -5.139921e-21, -1.798972e-20, -7.709882e-21, 
    -7.709882e-21, 5.139921e-21, 2.569961e-21, 2.569961e-21, -1.541976e-20, 
    -5.139921e-21, -2.569961e-21, -2.055969e-20, -1.541976e-20, 2.569961e-21, 
    -2.055969e-20, -1.28498e-20, -1.541976e-20, -5.139921e-21, 5.139921e-21, 
    -7.709882e-21, -1.003089e-36, -2.569961e-21, -1.027984e-20, 
    -2.569961e-21, -5.139921e-21, -1.28498e-20, -5.139921e-21, 0, 
    7.709882e-21, 0, 2.569961e-21, 1.027984e-20, -7.709882e-21, 1.28498e-20, 
    -5.139921e-21, 1.541976e-20, -1.798972e-20, -7.709882e-21, -7.709882e-21, 
    -1.027984e-20, -1.28498e-20, -1.003089e-36, 0, -1.027984e-20, 
    -1.003089e-36, -7.709882e-21, -2.569961e-21, 0, -1.798972e-20, 
    1.541976e-20, 1.28498e-20, -5.139921e-21, 1.027984e-20, 5.139921e-21, 
    -5.139921e-21, 1.027984e-20, -2.569961e-21, 1.541976e-20, -5.139921e-21, 
    -7.709882e-21, 1.003089e-36, 1.541976e-20, -7.709882e-21, -1.798972e-20, 
    2.569961e-21, -5.139921e-21, -2.569961e-21, 5.139921e-21, -1.027984e-20, 
    -2.569961e-21, -2.569961e-21, -1.28498e-20, -5.139921e-21, -2.569961e-21, 
    1.28498e-20, -7.709882e-21, 1.003089e-36, 1.003089e-36, -7.709882e-21, 
    -1.003089e-36, 1.541976e-20, 5.139921e-21, -1.027984e-20, 5.139921e-21, 
    5.139921e-21, 5.139921e-21, -5.139921e-21, -1.541976e-20, -1.027984e-20, 
    7.709882e-21, -1.003089e-36, 2.569961e-21, 2.569961e-21, 1.027984e-20, 
    2.312965e-20, 1.28498e-20, 2.569961e-21, -1.027984e-20, -7.709882e-21, 
    5.139921e-21, 7.709882e-21, 5.139921e-21, -1.28498e-20, 1.003089e-36, 
    -2.055969e-20, -1.027984e-20, 1.027984e-20, -7.709882e-21, -5.139921e-21, 
    -1.027984e-20, -7.709882e-21, -1.027984e-20, -7.709882e-21, 2.569961e-21, 
    -7.709882e-21, 0, 7.709882e-21, 5.139921e-21, -1.28498e-20, 0, 
    -7.709882e-21, 2.569961e-21, -2.569961e-21, -7.709882e-21, -1.003089e-36, 
    5.139921e-21, -7.709882e-21, -1.798972e-20, 1.003089e-36, 2.055969e-20, 
    -7.709882e-21, 2.569961e-21, 0, 7.709882e-21, -2.569961e-21, 
    -2.569961e-21, 3.009266e-36, -1.28498e-20, -1.541976e-20, -2.569961e-21, 
    -5.139921e-21, 5.139921e-21, 5.139921e-21, 2.055969e-20, 1.28498e-20, 
    5.139921e-21, -7.709882e-21, -7.709882e-21, 1.027984e-20, 1.541976e-20, 
    -5.139921e-21, -1.541976e-20, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    2.569961e-21, -1.027984e-20, 1.541976e-20, 2.569961e-21, 2.569961e-21, 
    7.709882e-21, 2.569961e-21, -2.569961e-21, 7.709882e-21, -5.139921e-21, 
    -1.003089e-36, 2.569961e-21, -1.541976e-20, -2.312965e-20, -2.569961e-21, 
    1.28498e-20, -2.569961e-21, 7.709882e-21, -1.28498e-20, 0, -2.569961e-21, 
    -7.709882e-21, -5.139921e-21, -1.027984e-20, 5.139921e-21, -7.709882e-21, 
    5.139921e-21, -5.139921e-21, 2.569961e-21, 7.709882e-21, 1.003089e-36, 
    1.027984e-20, -5.139921e-21, 1.027984e-20, 1.003089e-36, 1.798972e-20, 
    2.055969e-20, -7.709882e-21, 1.541976e-20, 1.027984e-20, -1.027984e-20, 
    -2.569961e-21, 1.027984e-20, 0, -2.569961e-21, -5.139921e-21, 
    2.312965e-20, -2.569961e-21, 2.569961e-21, 1.027984e-20, 1.541976e-20, 
    -2.569961e-21, -1.027984e-20, 1.003089e-36, -5.139921e-21, 1.003089e-36, 
    7.709882e-21, 0, -5.139921e-21, -1.027984e-20, -5.139921e-21, 
    1.003089e-36, -5.139921e-21, -1.027984e-20, 2.569961e-21, -7.709882e-21, 
    -7.709882e-21, 2.569961e-21, -1.003089e-36, 0, 2.569961e-21, 
    -2.569961e-21, -1.28498e-20, 7.709882e-21, -2.569961e-21, -1.798972e-20, 
    1.027984e-20, -1.027984e-20, -1.798972e-20, 7.709882e-21, 1.28498e-20, 
    -7.709882e-21, -7.709882e-21, 5.139921e-21, 0, -1.027984e-20, 
    -2.312965e-20, 2.569961e-21, 7.709882e-21, -7.709882e-21, -7.709882e-21, 
    -2.569961e-21, -2.569961e-21, 2.569961e-20, 7.709882e-21, 7.709882e-21, 
    2.569961e-21, 2.569961e-21, -5.139921e-21, -1.027984e-20, -2.569961e-21, 
    2.569961e-21, -1.28498e-20, 1.003089e-36, -5.139921e-21, -1.003089e-36, 
    -1.28498e-20, -1.027984e-20, -5.139921e-21, 1.003089e-36, 7.709882e-21, 
    -5.139921e-21, -2.569961e-21, -7.709882e-21, -1.003089e-36, 1.28498e-20, 
    5.139921e-21, 0, -1.003089e-36, -2.569961e-21, -1.28498e-20, 
    2.569961e-21, -1.027984e-20, -7.709882e-21, 5.139921e-21, 7.709882e-21, 
    5.139921e-21, -5.139921e-21, -1.28498e-20, 5.139921e-21, 1.027984e-20, 
    2.569961e-21, 1.003089e-36, 5.139921e-21, 1.28498e-20, -1.027984e-20, 
    -5.139921e-21, 0, 1.28498e-20, -2.569961e-21, 1.027984e-20, 1.027984e-20, 
    2.569961e-21, 0, 1.003089e-36, 5.139921e-21, 1.28498e-20, -1.003089e-36, 
    2.569961e-21, 2.569961e-21, 5.139921e-21, 2.569961e-21, 5.139921e-21, 
    1.027984e-20, 1.541976e-20, -1.027984e-20, -2.569961e-21, -7.709882e-21,
  -5.139921e-21, 5.139921e-21, 1.003089e-36, -1.027984e-20, 2.569961e-21, 
    1.28498e-20, 2.569961e-21, 1.027984e-20, -1.027984e-20, 5.139921e-21, 
    -5.139921e-21, 1.541976e-20, -5.139921e-21, 2.569961e-21, -2.569961e-21, 
    -1.541976e-20, 1.798972e-20, -1.027984e-20, -1.027984e-20, -7.709882e-21, 
    7.709882e-21, -1.541976e-20, -2.569961e-21, -1.798972e-20, -2.569961e-21, 
    -1.28498e-20, -1.28498e-20, -2.569961e-21, -1.28498e-20, -2.569961e-21, 
    1.003089e-36, -5.139921e-21, 2.569961e-21, 2.569961e-21, 0, 
    -3.009266e-36, 1.027984e-20, -5.139921e-21, 2.569961e-21, 2.569961e-21, 
    2.569961e-21, -1.027984e-20, -1.541976e-20, -1.28498e-20, 1.541976e-20, 
    -7.709882e-21, 2.569961e-21, -1.027984e-20, -5.139921e-21, 1.027984e-20, 
    -1.027984e-20, -1.28498e-20, 5.139921e-21, -1.003089e-36, 2.569961e-21, 
    -1.003089e-36, 1.541976e-20, -2.055969e-20, 5.139921e-21, 7.709882e-21, 
    -2.569961e-20, -1.027984e-20, -1.003089e-36, -1.28498e-20, -5.139921e-21, 
    7.709882e-21, -1.003089e-36, 2.569961e-21, -1.027984e-20, 2.055969e-20, 
    -1.003089e-36, 0, -1.003089e-36, -1.541976e-20, 1.541976e-20, 
    -2.569961e-21, -5.139921e-21, 0, 5.139921e-21, -1.003089e-36, 
    1.027984e-20, -7.709882e-21, -2.569961e-21, 2.826957e-20, 1.798972e-20, 
    2.569961e-21, 7.709882e-21, -1.027984e-20, -1.541976e-20, 5.139921e-21, 
    -7.709882e-21, 1.003089e-36, -1.027984e-20, 1.798972e-20, -1.541976e-20, 
    7.709882e-21, -1.027984e-20, 2.569961e-21, -2.569961e-21, 5.139921e-21, 
    2.569961e-21, -7.709882e-21, 1.541976e-20, -5.139921e-21, 1.798972e-20, 
    -7.709882e-21, -1.798972e-20, 1.28498e-20, 1.027984e-20, -2.569961e-21, 
    -5.139921e-21, 1.003089e-36, -2.569961e-20, -2.569961e-21, 2.569961e-21, 
    1.798972e-20, -2.569961e-21, -2.569961e-21, 2.569961e-21, -1.027984e-20, 
    2.569961e-21, 7.709882e-21, -2.569961e-21, 1.003089e-36, -1.003089e-36, 
    -5.139921e-21, -2.569961e-20, -5.139921e-21, -1.027984e-20, 
    -7.709882e-21, -5.139921e-21, -2.569961e-21, 5.139921e-21, -2.569961e-21, 
    3.340949e-20, -1.28498e-20, -5.139921e-21, -2.569961e-21, 1.28498e-20, 
    5.139921e-21, 1.541976e-20, -2.569961e-21, -7.709882e-21, -1.027984e-20, 
    -1.027984e-20, 7.709882e-21, -2.569961e-21, 7.709882e-21, -1.003089e-36, 
    -1.027984e-20, -1.003089e-36, 3.009266e-36, 1.027984e-20, -2.312965e-20, 
    2.569961e-21, 2.569961e-21, 5.139921e-21, 7.709882e-21, 1.027984e-20, 
    -1.027984e-20, 2.569961e-21, -1.28498e-20, 1.541976e-20, -1.541976e-20, 
    -5.139921e-21, 1.541976e-20, -2.569961e-21, 2.055969e-20, 7.709882e-21, 
    1.541976e-20, 1.541976e-20, 7.709882e-21, 2.569961e-21, 1.28498e-20, 
    5.139921e-21, 1.027984e-20, -1.28498e-20, 2.569961e-21, -2.569961e-21, 
    2.569961e-21, -2.569961e-21, 1.28498e-20, -1.798972e-20, 7.709882e-21, 
    -2.569961e-21, 2.569961e-21, -1.027984e-20, 1.541976e-20, -1.798972e-20, 
    -2.055969e-20, 5.139921e-21, -1.28498e-20, -1.28498e-20, -2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 1.541976e-20, -1.027984e-20, 1.541976e-20, 
    2.569961e-21, 1.541976e-20, -5.139921e-21, -7.709882e-21, -2.569961e-21, 
    -1.28498e-20, 7.709882e-21, -1.027984e-20, -2.569961e-21, -1.28498e-20, 
    -2.569961e-21, -7.709882e-21, -2.569961e-21, -1.003089e-36, 
    -7.709882e-21, 0, 2.312965e-20, -1.28498e-20, -5.139921e-21, 
    2.312965e-20, -5.139921e-21, -1.027984e-20, 5.139921e-21, -5.139921e-21, 
    2.569961e-21, -1.28498e-20, 3.340949e-20, -5.139921e-21, 1.798972e-20, 
    7.709882e-21, -5.139921e-21, 2.569961e-21, -1.541976e-20, -2.569961e-21, 
    -1.28498e-20, -1.541976e-20, -7.709882e-21, -7.709882e-21, -1.027984e-20, 
    0, -7.709882e-21, -7.709882e-21, 5.139921e-21, -5.139921e-21, 0, 
    1.003089e-36, 2.569961e-21, 5.139921e-21, -1.798972e-20, 5.139921e-21, 
    -1.003089e-36, -1.003089e-36, 2.569961e-21, 2.569961e-21, 1.003089e-36, 
    -2.055969e-20, -1.027984e-20, -1.027984e-20, -1.798972e-20, 7.709882e-21, 
    1.027984e-20, 5.139921e-21, -7.709882e-21, -5.139921e-21, -1.28498e-20, 
    7.709882e-21, 1.541976e-20, 3.340949e-20, -5.139921e-21, -1.027984e-20, 
    -1.28498e-20, 2.312965e-20, -5.139921e-21, 1.027984e-20, 1.541976e-20, 
    7.709882e-21, -5.139921e-21, -1.003089e-36, -5.139921e-21, -1.003089e-36, 
    -1.027984e-20, 1.027984e-20, -1.28498e-20, -2.569961e-21, -2.569961e-21, 
    -7.709882e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, 1.003089e-36, 
    -2.569961e-21, 1.541976e-20, 7.709882e-21, -5.139921e-21, 1.798972e-20, 
    1.798972e-20, 7.709882e-21, -5.139921e-21, -5.139921e-21, 7.709882e-21, 
    -7.709882e-21, -1.027984e-20, -1.541976e-20, 7.709882e-21, 0, 
    -1.027984e-20, 2.569961e-21, 1.003089e-36, -1.541976e-20, -1.027984e-20, 
    1.28498e-20, 1.003089e-36, -2.569961e-21, 5.139921e-21, -2.569961e-20, 
    -2.569961e-21, -7.709882e-21, 1.798972e-20, 2.569961e-20, 1.027984e-20, 
    1.28498e-20, -5.139921e-21, -1.798972e-20, 1.003089e-36, -1.541976e-20, 
    -1.798972e-20, 1.027984e-20, 2.569961e-21, -7.709882e-21, -5.139921e-21, 
    1.28498e-20, -7.709882e-21, 1.027984e-20, -1.027984e-20, 5.139921e-21, 
    -5.139921e-21, -2.055969e-20, -1.798972e-20, -7.709882e-21,
  6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.25807e-29, 6.258069e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.258069e-29, 6.25807e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.25807e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.25807e-29, 6.258069e-29, 6.258069e-29, 6.25807e-29, 6.258069e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.25807e-29, 6.258069e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.258069e-29, 6.25807e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.258069e-29, 6.25807e-29, 
    6.258069e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.258069e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.258069e-29, 
    6.258069e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.258069e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.258069e-29, 6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.258069e-29, 6.258069e-29, 6.258069e-29, 
    6.258069e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 6.25807e-29, 
    6.25807e-29, 6.25807e-29, 6.25807e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N_TO_SOIL1N =
  6.343376e-12, 6.36075e-12, 6.357374e-12, 6.371383e-12, 6.363613e-12, 
    6.372785e-12, 6.3469e-12, 6.361438e-12, 6.352158e-12, 6.344942e-12, 
    6.398558e-12, 6.372008e-12, 6.426137e-12, 6.409211e-12, 6.451725e-12, 
    6.423502e-12, 6.457415e-12, 6.450914e-12, 6.470486e-12, 6.46488e-12, 
    6.489901e-12, 6.473074e-12, 6.502872e-12, 6.485884e-12, 6.488541e-12, 
    6.472518e-12, 6.377355e-12, 6.395252e-12, 6.376294e-12, 6.378846e-12, 
    6.377701e-12, 6.363772e-12, 6.35675e-12, 6.34205e-12, 6.344719e-12, 
    6.355517e-12, 6.379994e-12, 6.371688e-12, 6.392624e-12, 6.392152e-12, 
    6.415451e-12, 6.404946e-12, 6.444096e-12, 6.432972e-12, 6.465114e-12, 
    6.457032e-12, 6.464734e-12, 6.462399e-12, 6.464764e-12, 6.452911e-12, 
    6.457989e-12, 6.447559e-12, 6.406913e-12, 6.41886e-12, 6.38322e-12, 
    6.361777e-12, 6.347537e-12, 6.337428e-12, 6.338857e-12, 6.341581e-12, 
    6.355581e-12, 6.368742e-12, 6.378769e-12, 6.385476e-12, 6.392084e-12, 
    6.412073e-12, 6.422657e-12, 6.446343e-12, 6.442072e-12, 6.44931e-12, 
    6.456228e-12, 6.467837e-12, 6.465926e-12, 6.47104e-12, 6.449121e-12, 
    6.463689e-12, 6.439638e-12, 6.446216e-12, 6.393871e-12, 6.37393e-12, 
    6.365444e-12, 6.358022e-12, 6.339956e-12, 6.352432e-12, 6.347514e-12, 
    6.359216e-12, 6.366649e-12, 6.362973e-12, 6.385659e-12, 6.37684e-12, 
    6.423284e-12, 6.403283e-12, 6.455421e-12, 6.442949e-12, 6.45841e-12, 
    6.450522e-12, 6.464037e-12, 6.451874e-12, 6.472944e-12, 6.47753e-12, 
    6.474396e-12, 6.486437e-12, 6.451199e-12, 6.464733e-12, 6.36287e-12, 
    6.363469e-12, 6.366263e-12, 6.353981e-12, 6.35323e-12, 6.341976e-12, 
    6.351991e-12, 6.356254e-12, 6.36708e-12, 6.373482e-12, 6.379567e-12, 
    6.392943e-12, 6.407878e-12, 6.428759e-12, 6.443757e-12, 6.453809e-12, 
    6.447646e-12, 6.453087e-12, 6.447004e-12, 6.444154e-12, 6.475811e-12, 
    6.458036e-12, 6.484706e-12, 6.483231e-12, 6.471161e-12, 6.483397e-12, 
    6.36389e-12, 6.36044e-12, 6.348458e-12, 6.357835e-12, 6.34075e-12, 
    6.350313e-12, 6.35581e-12, 6.377022e-12, 6.381684e-12, 6.386004e-12, 
    6.394536e-12, 6.405484e-12, 6.424684e-12, 6.441386e-12, 6.45663e-12, 
    6.455514e-12, 6.455907e-12, 6.459311e-12, 6.450877e-12, 6.460695e-12, 
    6.462342e-12, 6.458035e-12, 6.483033e-12, 6.475892e-12, 6.483199e-12, 
    6.47855e-12, 6.361562e-12, 6.367367e-12, 6.36423e-12, 6.370129e-12, 
    6.365973e-12, 6.384449e-12, 6.389987e-12, 6.415899e-12, 6.405268e-12, 
    6.422189e-12, 6.406988e-12, 6.409681e-12, 6.422737e-12, 6.40781e-12, 
    6.440463e-12, 6.418324e-12, 6.459443e-12, 6.437338e-12, 6.460828e-12, 
    6.456564e-12, 6.463624e-12, 6.469946e-12, 6.477899e-12, 6.492569e-12, 
    6.489172e-12, 6.50144e-12, 6.376022e-12, 6.383549e-12, 6.382888e-12, 
    6.390766e-12, 6.396591e-12, 6.409216e-12, 6.429459e-12, 6.421848e-12, 
    6.435821e-12, 6.438626e-12, 6.417397e-12, 6.43043e-12, 6.388588e-12, 
    6.395348e-12, 6.391324e-12, 6.376615e-12, 6.423599e-12, 6.39949e-12, 
    6.444005e-12, 6.43095e-12, 6.469044e-12, 6.4501e-12, 6.487302e-12, 
    6.503195e-12, 6.518157e-12, 6.535628e-12, 6.387658e-12, 6.382544e-12, 
    6.391703e-12, 6.404369e-12, 6.416124e-12, 6.431745e-12, 6.433345e-12, 
    6.43627e-12, 6.44385e-12, 6.450221e-12, 6.437194e-12, 6.451818e-12, 
    6.396913e-12, 6.425692e-12, 6.380609e-12, 6.394186e-12, 6.403623e-12, 
    6.399485e-12, 6.420979e-12, 6.426043e-12, 6.446617e-12, 6.435983e-12, 
    6.499271e-12, 6.471278e-12, 6.548933e-12, 6.527241e-12, 6.380757e-12, 
    6.387642e-12, 6.411596e-12, 6.4002e-12, 6.432789e-12, 6.440808e-12, 
    6.447327e-12, 6.455657e-12, 6.456558e-12, 6.461492e-12, 6.453405e-12, 
    6.461173e-12, 6.431779e-12, 6.444917e-12, 6.40886e-12, 6.417637e-12, 
    6.4136e-12, 6.409171e-12, 6.422841e-12, 6.437398e-12, 6.437712e-12, 
    6.442379e-12, 6.455522e-12, 6.432921e-12, 6.502878e-12, 6.459679e-12, 
    6.395148e-12, 6.408402e-12, 6.410299e-12, 6.405165e-12, 6.440003e-12, 
    6.427382e-12, 6.461372e-12, 6.452189e-12, 6.467236e-12, 6.459759e-12, 
    6.458659e-12, 6.449054e-12, 6.443073e-12, 6.427961e-12, 6.415662e-12, 
    6.40591e-12, 6.408178e-12, 6.41889e-12, 6.438289e-12, 6.456637e-12, 
    6.452618e-12, 6.466092e-12, 6.430427e-12, 6.445383e-12, 6.439602e-12, 
    6.454675e-12, 6.421646e-12, 6.449765e-12, 6.414455e-12, 6.417552e-12, 
    6.427132e-12, 6.446396e-12, 6.450661e-12, 6.45521e-12, 6.452403e-12, 
    6.438782e-12, 6.436551e-12, 6.426899e-12, 6.424233e-12, 6.416878e-12, 
    6.410787e-12, 6.416351e-12, 6.422194e-12, 6.438789e-12, 6.453739e-12, 
    6.470035e-12, 6.474024e-12, 6.493051e-12, 6.477559e-12, 6.503118e-12, 
    6.481383e-12, 6.519006e-12, 6.451398e-12, 6.480749e-12, 6.427569e-12, 
    6.433301e-12, 6.443664e-12, 6.467432e-12, 6.454605e-12, 6.469608e-12, 
    6.436464e-12, 6.419258e-12, 6.414809e-12, 6.406502e-12, 6.414999e-12, 
    6.414308e-12, 6.422438e-12, 6.419826e-12, 6.43934e-12, 6.428859e-12, 
    6.458631e-12, 6.46949e-12, 6.500154e-12, 6.518942e-12, 6.538067e-12, 
    6.546506e-12, 6.549075e-12, 6.550149e-12 ;

 SOIL3N_vr =
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.81819, 1.818189, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.818189, 1.81819, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.81819, 1.818189, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.818189, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.818189, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.818189, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.818189, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819,
  1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819,
  1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819,
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.81819, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.81819, 1.81819, 1.81819, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.81819, 1.81819, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.81819, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.81819, 1.818189, 1.81819, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.81819, 1.81819, 1.81819, 1.81819, 
    1.81819, 1.81819,
  1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 
    1.818189, 1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 
    1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818188, 
    1.818189, 1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3_HR =
  3.837742e-11, 3.848254e-11, 3.846211e-11, 3.854686e-11, 3.849986e-11, 
    3.855535e-11, 3.839875e-11, 3.84867e-11, 3.843056e-11, 3.83869e-11, 
    3.871127e-11, 3.855065e-11, 3.887813e-11, 3.877573e-11, 3.903294e-11, 
    3.886219e-11, 3.906736e-11, 3.902803e-11, 3.914644e-11, 3.911252e-11, 
    3.92639e-11, 3.916209e-11, 3.934238e-11, 3.92396e-11, 3.925567e-11, 
    3.915873e-11, 3.858299e-11, 3.869128e-11, 3.857658e-11, 3.859202e-11, 
    3.858509e-11, 3.850082e-11, 3.845834e-11, 3.83694e-11, 3.838555e-11, 
    3.845088e-11, 3.859896e-11, 3.854871e-11, 3.867538e-11, 3.867252e-11, 
    3.881348e-11, 3.874993e-11, 3.898678e-11, 3.891948e-11, 3.911394e-11, 
    3.906504e-11, 3.911164e-11, 3.909751e-11, 3.911182e-11, 3.904011e-11, 
    3.907083e-11, 3.900773e-11, 3.876182e-11, 3.88341e-11, 3.861848e-11, 
    3.848875e-11, 3.84026e-11, 3.834144e-11, 3.835009e-11, 3.836657e-11, 
    3.845126e-11, 3.853089e-11, 3.859156e-11, 3.863213e-11, 3.867211e-11, 
    3.879304e-11, 3.885707e-11, 3.900038e-11, 3.897454e-11, 3.901833e-11, 
    3.906018e-11, 3.913041e-11, 3.911885e-11, 3.914979e-11, 3.901718e-11, 
    3.910531e-11, 3.895981e-11, 3.899961e-11, 3.868292e-11, 3.856227e-11, 
    3.851093e-11, 3.846604e-11, 3.835673e-11, 3.843221e-11, 3.840246e-11, 
    3.847326e-11, 3.851823e-11, 3.849599e-11, 3.863324e-11, 3.857988e-11, 
    3.886087e-11, 3.873987e-11, 3.905529e-11, 3.897984e-11, 3.907338e-11, 
    3.902566e-11, 3.910742e-11, 3.903384e-11, 3.916131e-11, 3.918905e-11, 
    3.917009e-11, 3.924295e-11, 3.902976e-11, 3.911163e-11, 3.849536e-11, 
    3.849899e-11, 3.851589e-11, 3.844159e-11, 3.843704e-11, 3.836895e-11, 
    3.842954e-11, 3.845534e-11, 3.852084e-11, 3.855956e-11, 3.859638e-11, 
    3.86773e-11, 3.876766e-11, 3.889399e-11, 3.898473e-11, 3.904554e-11, 
    3.900826e-11, 3.904118e-11, 3.900438e-11, 3.898713e-11, 3.917866e-11, 
    3.907112e-11, 3.923247e-11, 3.922354e-11, 3.915053e-11, 3.922455e-11, 
    3.850154e-11, 3.848066e-11, 3.840817e-11, 3.84649e-11, 3.836154e-11, 
    3.841939e-11, 3.845265e-11, 3.858099e-11, 3.860919e-11, 3.863532e-11, 
    3.868695e-11, 3.875318e-11, 3.886934e-11, 3.897038e-11, 3.906261e-11, 
    3.905586e-11, 3.905824e-11, 3.907883e-11, 3.902781e-11, 3.908721e-11, 
    3.909717e-11, 3.907111e-11, 3.922235e-11, 3.917915e-11, 3.922335e-11, 
    3.919523e-11, 3.848745e-11, 3.852257e-11, 3.850359e-11, 3.853928e-11, 
    3.851414e-11, 3.862591e-11, 3.865942e-11, 3.881619e-11, 3.875187e-11, 
    3.885424e-11, 3.876227e-11, 3.877857e-11, 3.885756e-11, 3.876725e-11, 
    3.89648e-11, 3.883086e-11, 3.907963e-11, 3.894589e-11, 3.908801e-11, 
    3.906222e-11, 3.910493e-11, 3.914317e-11, 3.919129e-11, 3.928004e-11, 
    3.925949e-11, 3.933371e-11, 3.857493e-11, 3.862047e-11, 3.861647e-11, 
    3.866413e-11, 3.869937e-11, 3.877576e-11, 3.889822e-11, 3.885218e-11, 
    3.893672e-11, 3.895369e-11, 3.882526e-11, 3.890411e-11, 3.865095e-11, 
    3.869185e-11, 3.866751e-11, 3.857852e-11, 3.886278e-11, 3.871692e-11, 
    3.898623e-11, 3.890725e-11, 3.913772e-11, 3.902311e-11, 3.924818e-11, 
    3.934433e-11, 3.943485e-11, 3.954055e-11, 3.864533e-11, 3.861439e-11, 
    3.86698e-11, 3.874643e-11, 3.881755e-11, 3.891206e-11, 3.892173e-11, 
    3.893944e-11, 3.898529e-11, 3.902384e-11, 3.894502e-11, 3.90335e-11, 
    3.870132e-11, 3.887544e-11, 3.860268e-11, 3.868482e-11, 3.874192e-11, 
    3.871688e-11, 3.884692e-11, 3.887756e-11, 3.900203e-11, 3.89377e-11, 
    3.932059e-11, 3.915123e-11, 3.962105e-11, 3.94898e-11, 3.860358e-11, 
    3.864523e-11, 3.879016e-11, 3.872121e-11, 3.891838e-11, 3.896689e-11, 
    3.900633e-11, 3.905672e-11, 3.906217e-11, 3.909203e-11, 3.90431e-11, 
    3.90901e-11, 3.891226e-11, 3.899174e-11, 3.877361e-11, 3.88267e-11, 
    3.880228e-11, 3.877548e-11, 3.885819e-11, 3.894626e-11, 3.894816e-11, 
    3.897639e-11, 3.905591e-11, 3.891918e-11, 3.934241e-11, 3.908106e-11, 
    3.869065e-11, 3.877084e-11, 3.878231e-11, 3.875125e-11, 3.896202e-11, 
    3.888566e-11, 3.90913e-11, 3.903574e-11, 3.912678e-11, 3.908154e-11, 
    3.907488e-11, 3.901678e-11, 3.898059e-11, 3.888916e-11, 3.881476e-11, 
    3.875575e-11, 3.876948e-11, 3.883429e-11, 3.895165e-11, 3.906266e-11, 
    3.903834e-11, 3.911986e-11, 3.890408e-11, 3.899457e-11, 3.895959e-11, 
    3.905079e-11, 3.885096e-11, 3.902108e-11, 3.880745e-11, 3.882619e-11, 
    3.888415e-11, 3.900069e-11, 3.90265e-11, 3.905402e-11, 3.903704e-11, 
    3.895463e-11, 3.894114e-11, 3.888274e-11, 3.886661e-11, 3.882211e-11, 
    3.878526e-11, 3.881893e-11, 3.885427e-11, 3.895467e-11, 3.904512e-11, 
    3.914371e-11, 3.916785e-11, 3.928296e-11, 3.918923e-11, 3.934386e-11, 
    3.921237e-11, 3.943999e-11, 3.903096e-11, 3.920853e-11, 3.888679e-11, 
    3.892147e-11, 3.898417e-11, 3.912796e-11, 3.905036e-11, 3.914113e-11, 
    3.894061e-11, 3.883651e-11, 3.88096e-11, 3.875934e-11, 3.881075e-11, 
    3.880657e-11, 3.885575e-11, 3.883995e-11, 3.895801e-11, 3.88946e-11, 
    3.907471e-11, 3.914042e-11, 3.932593e-11, 3.94396e-11, 3.95553e-11, 
    3.960636e-11, 3.962191e-11, 3.96284e-11 ;

 SOILC =
  17.34412, 17.34411, 17.34411, 17.3441, 17.34411, 17.3441, 17.34412, 
    17.34411, 17.34411, 17.34412, 17.34409, 17.3441, 17.34407, 17.34408, 
    17.34406, 17.34407, 17.34406, 17.34406, 17.34405, 17.34405, 17.34404, 
    17.34405, 17.34403, 17.34404, 17.34404, 17.34405, 17.3441, 17.34409, 
    17.3441, 17.3441, 17.3441, 17.34411, 17.34411, 17.34412, 17.34412, 
    17.34411, 17.3441, 17.3441, 17.34409, 17.34409, 17.34408, 17.34408, 
    17.34406, 17.34407, 17.34405, 17.34406, 17.34405, 17.34405, 17.34405, 
    17.34406, 17.34405, 17.34406, 17.34408, 17.34408, 17.3441, 17.34411, 
    17.34412, 17.34412, 17.34412, 17.34412, 17.34411, 17.3441, 17.3441, 
    17.3441, 17.34409, 17.34408, 17.34407, 17.34406, 17.34406, 17.34406, 
    17.34406, 17.34405, 17.34405, 17.34405, 17.34406, 17.34405, 17.34406, 
    17.34406, 17.34409, 17.3441, 17.34411, 17.34411, 17.34412, 17.34411, 
    17.34412, 17.34411, 17.34411, 17.34411, 17.3441, 17.3441, 17.34407, 
    17.34409, 17.34406, 17.34406, 17.34405, 17.34406, 17.34405, 17.34406, 
    17.34405, 17.34404, 17.34405, 17.34404, 17.34406, 17.34405, 17.34411, 
    17.34411, 17.34411, 17.34411, 17.34411, 17.34412, 17.34411, 17.34411, 
    17.34411, 17.3441, 17.3441, 17.34409, 17.34408, 17.34407, 17.34406, 
    17.34406, 17.34406, 17.34406, 17.34406, 17.34406, 17.34404, 17.34405, 
    17.34404, 17.34404, 17.34405, 17.34404, 17.34411, 17.34411, 17.34412, 
    17.34411, 17.34412, 17.34412, 17.34411, 17.3441, 17.3441, 17.3441, 
    17.34409, 17.34408, 17.34407, 17.34406, 17.34406, 17.34406, 17.34406, 
    17.34405, 17.34406, 17.34405, 17.34405, 17.34405, 17.34404, 17.34404, 
    17.34404, 17.34404, 17.34411, 17.34411, 17.34411, 17.3441, 17.34411, 
    17.3441, 17.34409, 17.34408, 17.34408, 17.34407, 17.34408, 17.34408, 
    17.34407, 17.34408, 17.34406, 17.34408, 17.34405, 17.34407, 17.34405, 
    17.34406, 17.34405, 17.34405, 17.34404, 17.34403, 17.34404, 17.34403, 
    17.3441, 17.3441, 17.3441, 17.34409, 17.34409, 17.34408, 17.34407, 
    17.34407, 17.34407, 17.34406, 17.34408, 17.34407, 17.34409, 17.34409, 
    17.34409, 17.3441, 17.34407, 17.34409, 17.34406, 17.34407, 17.34405, 
    17.34406, 17.34404, 17.34403, 17.34402, 17.34401, 17.3441, 17.3441, 
    17.34409, 17.34409, 17.34408, 17.34407, 17.34407, 17.34407, 17.34406, 
    17.34406, 17.34407, 17.34406, 17.34409, 17.34407, 17.3441, 17.34409, 
    17.34409, 17.34409, 17.34408, 17.34407, 17.34406, 17.34407, 17.34403, 
    17.34405, 17.344, 17.34402, 17.3441, 17.3441, 17.34408, 17.34409, 
    17.34407, 17.34406, 17.34406, 17.34406, 17.34406, 17.34405, 17.34406, 
    17.34405, 17.34407, 17.34406, 17.34408, 17.34408, 17.34408, 17.34408, 
    17.34407, 17.34407, 17.34407, 17.34406, 17.34406, 17.34407, 17.34403, 
    17.34405, 17.34409, 17.34408, 17.34408, 17.34408, 17.34406, 17.34407, 
    17.34405, 17.34406, 17.34405, 17.34405, 17.34405, 17.34406, 17.34406, 
    17.34407, 17.34408, 17.34408, 17.34408, 17.34408, 17.34406, 17.34406, 
    17.34406, 17.34405, 17.34407, 17.34406, 17.34406, 17.34406, 17.34407, 
    17.34406, 17.34408, 17.34408, 17.34407, 17.34406, 17.34406, 17.34406, 
    17.34406, 17.34406, 17.34407, 17.34407, 17.34407, 17.34408, 17.34408, 
    17.34408, 17.34407, 17.34406, 17.34406, 17.34405, 17.34405, 17.34403, 
    17.34404, 17.34403, 17.34404, 17.34402, 17.34406, 17.34404, 17.34407, 
    17.34407, 17.34406, 17.34405, 17.34406, 17.34405, 17.34407, 17.34408, 
    17.34408, 17.34408, 17.34408, 17.34408, 17.34407, 17.34408, 17.34406, 
    17.34407, 17.34405, 17.34405, 17.34403, 17.34402, 17.34401, 17.344, 
    17.344, 17.344 ;

 SOILC_HR =
  7.62417e-08, 7.645039e-08, 7.640983e-08, 7.657811e-08, 7.648478e-08, 
    7.659495e-08, 7.628402e-08, 7.645866e-08, 7.634719e-08, 7.626051e-08, 
    7.690453e-08, 7.658562e-08, 7.72358e-08, 7.70325e-08, 7.754317e-08, 
    7.720416e-08, 7.761152e-08, 7.753343e-08, 7.776852e-08, 7.770118e-08, 
    7.800173e-08, 7.77996e-08, 7.815754e-08, 7.795349e-08, 7.79854e-08, 
    7.779293e-08, 7.664984e-08, 7.686482e-08, 7.663709e-08, 7.666775e-08, 
    7.6654e-08, 7.648669e-08, 7.640234e-08, 7.622577e-08, 7.625783e-08, 
    7.638754e-08, 7.668154e-08, 7.658178e-08, 7.683326e-08, 7.682758e-08, 
    7.710744e-08, 7.698127e-08, 7.745152e-08, 7.731791e-08, 7.770399e-08, 
    7.760691e-08, 7.769943e-08, 7.767138e-08, 7.769979e-08, 7.755741e-08, 
    7.761841e-08, 7.749312e-08, 7.700489e-08, 7.71484e-08, 7.67203e-08, 
    7.646273e-08, 7.629168e-08, 7.617025e-08, 7.618742e-08, 7.622014e-08, 
    7.63883e-08, 7.654639e-08, 7.666684e-08, 7.674739e-08, 7.682677e-08, 
    7.706688e-08, 7.719401e-08, 7.747852e-08, 7.742722e-08, 7.751416e-08, 
    7.759725e-08, 7.773669e-08, 7.771375e-08, 7.777518e-08, 7.751189e-08, 
    7.768687e-08, 7.739798e-08, 7.7477e-08, 7.684823e-08, 7.66087e-08, 
    7.650677e-08, 7.641763e-08, 7.620062e-08, 7.635047e-08, 7.62914e-08, 
    7.643196e-08, 7.652125e-08, 7.647709e-08, 7.674959e-08, 7.664367e-08, 
    7.720153e-08, 7.696129e-08, 7.758756e-08, 7.743775e-08, 7.762347e-08, 
    7.752871e-08, 7.769106e-08, 7.754495e-08, 7.779804e-08, 7.785313e-08, 
    7.781549e-08, 7.796012e-08, 7.753685e-08, 7.769941e-08, 7.647585e-08, 
    7.648305e-08, 7.651661e-08, 7.636908e-08, 7.636006e-08, 7.622488e-08, 
    7.634518e-08, 7.639639e-08, 7.652643e-08, 7.660332e-08, 7.667641e-08, 
    7.683709e-08, 7.701648e-08, 7.726729e-08, 7.744746e-08, 7.75682e-08, 
    7.749417e-08, 7.755953e-08, 7.748646e-08, 7.745222e-08, 7.783248e-08, 
    7.761898e-08, 7.793933e-08, 7.792161e-08, 7.777663e-08, 7.79236e-08, 
    7.648811e-08, 7.644667e-08, 7.630274e-08, 7.641538e-08, 7.621016e-08, 
    7.632502e-08, 7.639106e-08, 7.664585e-08, 7.670185e-08, 7.675374e-08, 
    7.685622e-08, 7.698772e-08, 7.721835e-08, 7.741897e-08, 7.760209e-08, 
    7.758867e-08, 7.75934e-08, 7.763429e-08, 7.753298e-08, 7.765092e-08, 
    7.76707e-08, 7.761896e-08, 7.791923e-08, 7.783346e-08, 7.792123e-08, 
    7.786539e-08, 7.646015e-08, 7.652987e-08, 7.649219e-08, 7.656304e-08, 
    7.651312e-08, 7.673505e-08, 7.680158e-08, 7.711283e-08, 7.698513e-08, 
    7.718838e-08, 7.700579e-08, 7.703814e-08, 7.719496e-08, 7.701567e-08, 
    7.740789e-08, 7.714196e-08, 7.763587e-08, 7.737035e-08, 7.765251e-08, 
    7.76013e-08, 7.76861e-08, 7.776203e-08, 7.785756e-08, 7.803377e-08, 
    7.799298e-08, 7.814034e-08, 7.663383e-08, 7.672424e-08, 7.67163e-08, 
    7.681093e-08, 7.68809e-08, 7.703256e-08, 7.727571e-08, 7.718429e-08, 
    7.735214e-08, 7.738582e-08, 7.713083e-08, 7.728738e-08, 7.678477e-08, 
    7.686597e-08, 7.681763e-08, 7.664095e-08, 7.720533e-08, 7.691573e-08, 
    7.745043e-08, 7.729361e-08, 7.77512e-08, 7.752365e-08, 7.797052e-08, 
    7.816141e-08, 7.834114e-08, 7.8551e-08, 7.677361e-08, 7.671218e-08, 
    7.682219e-08, 7.697433e-08, 7.711554e-08, 7.730318e-08, 7.732238e-08, 
    7.735753e-08, 7.744857e-08, 7.75251e-08, 7.736862e-08, 7.754428e-08, 
    7.688477e-08, 7.723047e-08, 7.668893e-08, 7.685201e-08, 7.696537e-08, 
    7.691567e-08, 7.717384e-08, 7.723467e-08, 7.748181e-08, 7.735408e-08, 
    7.811428e-08, 7.777804e-08, 7.871082e-08, 7.845025e-08, 7.669071e-08, 
    7.677341e-08, 7.706114e-08, 7.692425e-08, 7.731571e-08, 7.741203e-08, 
    7.749034e-08, 7.759039e-08, 7.760121e-08, 7.766049e-08, 7.756335e-08, 
    7.765666e-08, 7.730358e-08, 7.746139e-08, 7.702828e-08, 7.713371e-08, 
    7.708522e-08, 7.703201e-08, 7.719621e-08, 7.737107e-08, 7.737484e-08, 
    7.74309e-08, 7.758878e-08, 7.73173e-08, 7.815761e-08, 7.763871e-08, 
    7.686358e-08, 7.702278e-08, 7.704556e-08, 7.698389e-08, 7.740237e-08, 
    7.725077e-08, 7.765905e-08, 7.754873e-08, 7.772948e-08, 7.763967e-08, 
    7.762645e-08, 7.751108e-08, 7.743924e-08, 7.725771e-08, 7.710998e-08, 
    7.699284e-08, 7.702008e-08, 7.714876e-08, 7.738178e-08, 7.760217e-08, 
    7.75539e-08, 7.771575e-08, 7.728734e-08, 7.746699e-08, 7.739755e-08, 
    7.75786e-08, 7.718186e-08, 7.751962e-08, 7.709549e-08, 7.713269e-08, 
    7.724775e-08, 7.747915e-08, 7.753039e-08, 7.758502e-08, 7.755131e-08, 
    7.73877e-08, 7.73609e-08, 7.724496e-08, 7.721293e-08, 7.712459e-08, 
    7.705142e-08, 7.711827e-08, 7.718845e-08, 7.738778e-08, 7.756736e-08, 
    7.77631e-08, 7.781102e-08, 7.803957e-08, 7.785348e-08, 7.81605e-08, 
    7.789941e-08, 7.835134e-08, 7.753925e-08, 7.789179e-08, 7.7253e-08, 
    7.732185e-08, 7.744634e-08, 7.773184e-08, 7.757776e-08, 7.775797e-08, 
    7.735986e-08, 7.715318e-08, 7.709974e-08, 7.699995e-08, 7.710202e-08, 
    7.709372e-08, 7.719137e-08, 7.716e-08, 7.73944e-08, 7.72685e-08, 
    7.762611e-08, 7.775656e-08, 7.812488e-08, 7.835057e-08, 7.858029e-08, 
    7.868167e-08, 7.871252e-08, 7.872543e-08 ;

 SOILC_LOSS =
  7.62417e-08, 7.645039e-08, 7.640983e-08, 7.657811e-08, 7.648478e-08, 
    7.659495e-08, 7.628402e-08, 7.645866e-08, 7.634719e-08, 7.626051e-08, 
    7.690453e-08, 7.658562e-08, 7.72358e-08, 7.70325e-08, 7.754317e-08, 
    7.720416e-08, 7.761152e-08, 7.753343e-08, 7.776852e-08, 7.770118e-08, 
    7.800173e-08, 7.77996e-08, 7.815754e-08, 7.795349e-08, 7.79854e-08, 
    7.779293e-08, 7.664984e-08, 7.686482e-08, 7.663709e-08, 7.666775e-08, 
    7.6654e-08, 7.648669e-08, 7.640234e-08, 7.622577e-08, 7.625783e-08, 
    7.638754e-08, 7.668154e-08, 7.658178e-08, 7.683326e-08, 7.682758e-08, 
    7.710744e-08, 7.698127e-08, 7.745152e-08, 7.731791e-08, 7.770399e-08, 
    7.760691e-08, 7.769943e-08, 7.767138e-08, 7.769979e-08, 7.755741e-08, 
    7.761841e-08, 7.749312e-08, 7.700489e-08, 7.71484e-08, 7.67203e-08, 
    7.646273e-08, 7.629168e-08, 7.617025e-08, 7.618742e-08, 7.622014e-08, 
    7.63883e-08, 7.654639e-08, 7.666684e-08, 7.674739e-08, 7.682677e-08, 
    7.706688e-08, 7.719401e-08, 7.747852e-08, 7.742722e-08, 7.751416e-08, 
    7.759725e-08, 7.773669e-08, 7.771375e-08, 7.777518e-08, 7.751189e-08, 
    7.768687e-08, 7.739798e-08, 7.7477e-08, 7.684823e-08, 7.66087e-08, 
    7.650677e-08, 7.641763e-08, 7.620062e-08, 7.635047e-08, 7.62914e-08, 
    7.643196e-08, 7.652125e-08, 7.647709e-08, 7.674959e-08, 7.664367e-08, 
    7.720153e-08, 7.696129e-08, 7.758756e-08, 7.743775e-08, 7.762347e-08, 
    7.752871e-08, 7.769106e-08, 7.754495e-08, 7.779804e-08, 7.785313e-08, 
    7.781549e-08, 7.796012e-08, 7.753685e-08, 7.769941e-08, 7.647585e-08, 
    7.648305e-08, 7.651661e-08, 7.636908e-08, 7.636006e-08, 7.622488e-08, 
    7.634518e-08, 7.639639e-08, 7.652643e-08, 7.660332e-08, 7.667641e-08, 
    7.683709e-08, 7.701648e-08, 7.726729e-08, 7.744746e-08, 7.75682e-08, 
    7.749417e-08, 7.755953e-08, 7.748646e-08, 7.745222e-08, 7.783248e-08, 
    7.761898e-08, 7.793933e-08, 7.792161e-08, 7.777663e-08, 7.79236e-08, 
    7.648811e-08, 7.644667e-08, 7.630274e-08, 7.641538e-08, 7.621016e-08, 
    7.632502e-08, 7.639106e-08, 7.664585e-08, 7.670185e-08, 7.675374e-08, 
    7.685622e-08, 7.698772e-08, 7.721835e-08, 7.741897e-08, 7.760209e-08, 
    7.758867e-08, 7.75934e-08, 7.763429e-08, 7.753298e-08, 7.765092e-08, 
    7.76707e-08, 7.761896e-08, 7.791923e-08, 7.783346e-08, 7.792123e-08, 
    7.786539e-08, 7.646015e-08, 7.652987e-08, 7.649219e-08, 7.656304e-08, 
    7.651312e-08, 7.673505e-08, 7.680158e-08, 7.711283e-08, 7.698513e-08, 
    7.718838e-08, 7.700579e-08, 7.703814e-08, 7.719496e-08, 7.701567e-08, 
    7.740789e-08, 7.714196e-08, 7.763587e-08, 7.737035e-08, 7.765251e-08, 
    7.76013e-08, 7.76861e-08, 7.776203e-08, 7.785756e-08, 7.803377e-08, 
    7.799298e-08, 7.814034e-08, 7.663383e-08, 7.672424e-08, 7.67163e-08, 
    7.681093e-08, 7.68809e-08, 7.703256e-08, 7.727571e-08, 7.718429e-08, 
    7.735214e-08, 7.738582e-08, 7.713083e-08, 7.728738e-08, 7.678477e-08, 
    7.686597e-08, 7.681763e-08, 7.664095e-08, 7.720533e-08, 7.691573e-08, 
    7.745043e-08, 7.729361e-08, 7.77512e-08, 7.752365e-08, 7.797052e-08, 
    7.816141e-08, 7.834114e-08, 7.8551e-08, 7.677361e-08, 7.671218e-08, 
    7.682219e-08, 7.697433e-08, 7.711554e-08, 7.730318e-08, 7.732238e-08, 
    7.735753e-08, 7.744857e-08, 7.75251e-08, 7.736862e-08, 7.754428e-08, 
    7.688477e-08, 7.723047e-08, 7.668893e-08, 7.685201e-08, 7.696537e-08, 
    7.691567e-08, 7.717384e-08, 7.723467e-08, 7.748181e-08, 7.735408e-08, 
    7.811428e-08, 7.777804e-08, 7.871082e-08, 7.845025e-08, 7.669071e-08, 
    7.677341e-08, 7.706114e-08, 7.692425e-08, 7.731571e-08, 7.741203e-08, 
    7.749034e-08, 7.759039e-08, 7.760121e-08, 7.766049e-08, 7.756335e-08, 
    7.765666e-08, 7.730358e-08, 7.746139e-08, 7.702828e-08, 7.713371e-08, 
    7.708522e-08, 7.703201e-08, 7.719621e-08, 7.737107e-08, 7.737484e-08, 
    7.74309e-08, 7.758878e-08, 7.73173e-08, 7.815761e-08, 7.763871e-08, 
    7.686358e-08, 7.702278e-08, 7.704556e-08, 7.698389e-08, 7.740237e-08, 
    7.725077e-08, 7.765905e-08, 7.754873e-08, 7.772948e-08, 7.763967e-08, 
    7.762645e-08, 7.751108e-08, 7.743924e-08, 7.725771e-08, 7.710998e-08, 
    7.699284e-08, 7.702008e-08, 7.714876e-08, 7.738178e-08, 7.760217e-08, 
    7.75539e-08, 7.771575e-08, 7.728734e-08, 7.746699e-08, 7.739755e-08, 
    7.75786e-08, 7.718186e-08, 7.751962e-08, 7.709549e-08, 7.713269e-08, 
    7.724775e-08, 7.747915e-08, 7.753039e-08, 7.758502e-08, 7.755131e-08, 
    7.73877e-08, 7.73609e-08, 7.724496e-08, 7.721293e-08, 7.712459e-08, 
    7.705142e-08, 7.711827e-08, 7.718845e-08, 7.738778e-08, 7.756736e-08, 
    7.77631e-08, 7.781102e-08, 7.803957e-08, 7.785348e-08, 7.81605e-08, 
    7.789941e-08, 7.835134e-08, 7.753925e-08, 7.789179e-08, 7.7253e-08, 
    7.732185e-08, 7.744634e-08, 7.773184e-08, 7.757776e-08, 7.775797e-08, 
    7.735986e-08, 7.715318e-08, 7.709974e-08, 7.699995e-08, 7.710202e-08, 
    7.709372e-08, 7.719137e-08, 7.716e-08, 7.73944e-08, 7.72685e-08, 
    7.762611e-08, 7.775656e-08, 7.812488e-08, 7.835057e-08, 7.858029e-08, 
    7.868167e-08, 7.871252e-08, 7.872543e-08 ;

 SOILICE =
  98.96801, 99.40324, 99.31853, 99.67024, 99.47503, 99.70547, 99.05614, 
    99.42056, 99.18781, 99.00712, 100.355, 99.68594, 101.0525, 100.6238, 
    101.7027, 100.9857, 101.8476, 101.6819, 102.1809, 102.0378, 102.6777, 
    102.2469, 103.0101, 102.5747, 102.6427, 102.2328, 99.82032, 100.2716, 
    99.79363, 99.85789, 99.82905, 99.47907, 99.30302, 98.93476, 99.00155, 
    99.27203, 99.8868, 99.67783, 100.2049, 100.193, 100.7816, 100.516, 
    101.5084, 101.2257, 102.0437, 101.8377, 102.0341, 101.9745, 102.0348, 
    101.7327, 101.8621, 101.5965, 100.5657, 100.868, 99.96798, 99.42916, 
    99.07211, 98.81924, 98.85497, 98.9231, 99.27362, 99.60381, 99.85588, 
    100.0247, 100.1912, 100.6964, 100.9643, 101.5656, 101.4569, 101.6411, 
    101.8172, 102.1133, 102.0645, 102.1951, 101.6362, 102.0074, 101.395, 
    101.5623, 100.2367, 99.73417, 99.52116, 99.33482, 98.88245, 99.19472, 
    99.07156, 99.36469, 99.55124, 99.45894, 100.0293, 99.80737, 100.9802, 
    100.474, 101.7966, 101.4792, 101.8728, 101.6718, 102.0163, 101.7063, 
    102.2437, 102.3609, 102.2808, 102.5887, 101.6891, 102.0341, 99.45636, 
    99.47141, 99.54153, 99.23354, 99.21471, 98.93294, 99.18362, 99.2905, 
    99.56205, 99.72292, 99.87596, 100.213, 100.5901, 101.1189, 101.4998, 
    101.7555, 101.5987, 101.7372, 101.5823, 101.5098, 102.317, 101.8633, 
    102.5444, 102.5067, 102.1982, 102.5109, 99.48198, 99.39539, 99.09515, 
    99.33006, 98.90228, 99.14162, 99.27941, 99.81204, 99.92924, 100.0381, 
    100.2531, 100.5296, 101.0156, 101.4395, 101.8274, 101.799, 101.809, 
    101.8958, 101.6809, 101.9311, 101.9731, 101.8632, 102.5016, 102.319, 
    102.5059, 102.3869, 99.42352, 99.56927, 99.4905, 99.63866, 99.53429, 
    99.99897, 100.1385, 100.7931, 100.5241, 100.9524, 100.5676, 100.6357, 
    100.9664, 100.5883, 101.4162, 100.8546, 101.8991, 101.3368, 101.9344, 
    101.8257, 102.0057, 102.1671, 102.3703, 102.7459, 102.6588, 102.9733, 
    99.78677, 99.97626, 99.95953, 100.158, 100.305, 100.6239, 101.1366, 
    100.9436, 101.2981, 101.3693, 100.8309, 101.1613, 100.1032, 100.2737, 
    100.1721, 99.80173, 100.9881, 100.3783, 101.5061, 101.1744, 102.1441, 
    101.6612, 102.6109, 103.0185, 103.4028, 103.8531, 100.0797, 99.95088, 
    100.1816, 100.5015, 100.7987, 101.1947, 101.2352, 101.3095, 101.5021, 
    101.6642, 101.333, 101.7048, 100.3134, 101.0412, 99.90222, 100.2444, 
    100.4826, 100.378, 100.9216, 101.0499, 101.5726, 101.3022, 102.9179, 
    102.2013, 104.1966, 103.6369, 99.90589, 100.0793, 100.6841, 100.3961, 
    101.2211, 101.4248, 101.5905, 101.8027, 101.8256, 101.9514, 101.7453, 
    101.9432, 101.1955, 101.5293, 100.6149, 100.837, 100.7348, 100.6227, 
    100.9688, 101.3383, 101.3461, 101.4648, 101.7997, 101.2244, 103.0107, 
    101.9055, 100.2685, 100.6035, 100.6513, 100.5214, 101.4044, 101.0839, 
    101.9483, 101.7143, 102.0979, 101.9072, 101.8791, 101.6345, 101.4824, 
    101.0986, 100.787, 100.5403, 100.5976, 100.8688, 101.3609, 101.8277, 
    101.7253, 102.0687, 101.1611, 101.5412, 101.3942, 101.7776, 100.9385, 
    101.653, 100.7564, 100.8348, 101.0776, 101.567, 101.6754, 101.7913, 
    101.7198, 101.3734, 101.3167, 101.0717, 101.0041, 100.8177, 100.6636, 
    100.8044, 100.9525, 101.3735, 101.7538, 102.1694, 102.2712, 102.7585, 
    102.3618, 103.0169, 102.4599, 103.4251, 101.6944, 102.4435, 101.0886, 
    101.2341, 101.4975, 102.1031, 101.7758, 102.1586, 101.3144, 100.8781, 
    100.7654, 100.5553, 100.7702, 100.7527, 100.9586, 100.8924, 101.3875, 
    101.1214, 101.8784, 102.1556, 102.9404, 103.4232, 103.9159, 104.1338, 
    104.2002, 104.228,
  115.3993, 115.8093, 115.7295, 116.0607, 115.8768, 116.0938, 115.4823, 
    115.8256, 115.6063, 115.4361, 116.705, 116.0754, 117.3605, 116.9576, 
    117.9709, 117.2978, 118.1068, 117.9513, 118.4194, 118.2852, 118.8852, 
    118.4814, 119.1967, 118.7886, 118.8525, 118.4681, 116.2019, 116.6266, 
    116.1768, 116.2373, 116.2101, 115.8807, 115.7149, 115.3679, 115.4308, 
    115.6857, 116.2645, 116.0677, 116.5636, 116.5524, 117.1059, 116.8562, 
    117.7885, 117.5231, 118.2908, 118.0975, 118.2817, 118.2258, 118.2824, 
    117.999, 118.1204, 117.8711, 116.903, 117.1871, 116.3408, 115.8338, 
    115.4974, 115.259, 115.2927, 115.357, 115.6872, 115.9981, 116.2353, 
    116.3942, 116.5508, 117.026, 117.2776, 117.8423, 117.7401, 117.9131, 
    118.0783, 118.356, 118.3102, 118.4327, 117.9084, 118.2568, 117.682, 
    117.8391, 116.5938, 116.1208, 115.9204, 115.7448, 115.3186, 115.6129, 
    115.4968, 115.7729, 115.9486, 115.8617, 116.3985, 116.1897, 117.2925, 
    116.8168, 118.059, 117.7611, 118.1304, 117.9419, 118.2651, 117.9742, 
    118.4783, 118.5883, 118.5131, 118.8018, 117.9581, 118.2818, 115.8593, 
    115.8734, 115.9394, 115.6494, 115.6317, 115.3662, 115.6024, 115.7031, 
    115.9587, 116.1102, 116.2542, 116.5713, 116.926, 117.4228, 117.7804, 
    118.0204, 117.8732, 118.0032, 117.8579, 117.7898, 118.5471, 118.1216, 
    118.7602, 118.7248, 118.4357, 118.7288, 115.8834, 115.8018, 115.5191, 
    115.7403, 115.3373, 115.5628, 115.6927, 116.1941, 116.3044, 116.4068, 
    116.609, 116.869, 117.3257, 117.7239, 118.0879, 118.0612, 118.0706, 
    118.152, 117.9504, 118.1851, 118.2246, 118.1215, 118.7201, 118.5489, 
    118.7241, 118.6126, 115.8283, 115.9656, 115.8914, 116.0309, 115.9326, 
    116.37, 116.5014, 117.1167, 116.8639, 117.2663, 116.9047, 116.9688, 
    117.2797, 116.9242, 117.702, 117.1745, 118.1552, 117.6275, 118.1883, 
    118.0863, 118.2551, 118.4065, 118.597, 118.9491, 118.8675, 119.1621, 
    116.1703, 116.3486, 116.3329, 116.5196, 116.6578, 116.9576, 117.4394, 
    117.2581, 117.591, 117.6579, 117.1521, 117.4626, 116.468, 116.6285, 
    116.5329, 116.1844, 117.3, 116.7268, 117.7863, 117.4749, 118.3849, 
    117.932, 118.8226, 119.2046, 119.5643, 119.9858, 116.446, 116.3247, 
    116.5418, 116.8426, 117.1219, 117.4939, 117.532, 117.6017, 117.7825, 
    117.9347, 117.6239, 117.9728, 116.6659, 117.3498, 116.279, 116.601, 
    116.8249, 116.7265, 117.2374, 117.358, 117.8487, 117.5949, 119.1103, 
    118.4386, 120.307, 119.7834, 116.2824, 116.4455, 117.0143, 116.7435, 
    117.5187, 117.71, 117.8655, 118.0647, 118.0861, 118.2042, 118.0108, 
    118.1965, 117.4947, 117.808, 116.9491, 117.1579, 117.0618, 116.9565, 
    117.2817, 117.6288, 117.6361, 117.7475, 118.0621, 117.5219, 119.1974, 
    118.1614, 116.6235, 116.9385, 116.9834, 116.8613, 117.6908, 117.3899, 
    118.2013, 117.9817, 118.3416, 118.1627, 118.1364, 117.9068, 117.764, 
    117.4037, 117.111, 116.879, 116.9329, 117.1878, 117.65, 118.0881, 
    117.9921, 118.3142, 117.4624, 117.8193, 117.6813, 118.0412, 117.2533, 
    117.9244, 117.0821, 117.1558, 117.3839, 117.8436, 117.9452, 118.054, 
    117.9868, 117.6618, 117.6085, 117.3784, 117.3149, 117.1398, 116.9949, 
    117.1273, 117.2664, 117.6618, 118.0188, 118.4087, 118.5041, 118.961, 
    118.5892, 119.2032, 118.6814, 119.5853, 117.9632, 118.6658, 117.3943, 
    117.5309, 117.7783, 118.3466, 118.0395, 118.3986, 117.6064, 117.1966, 
    117.0906, 116.8931, 117.0951, 117.0787, 117.2721, 117.2099, 117.675, 
    117.425, 118.1358, 118.3957, 119.1313, 119.5835, 120.0444, 120.2483, 
    120.3103, 120.3363,
  168.5663, 169.1457, 169.0329, 169.501, 169.2412, 169.5479, 168.6836, 
    169.1688, 168.8589, 168.6183, 170.4117, 169.5219, 171.3382, 170.7687, 
    172.2011, 171.2496, 172.3932, 172.1734, 172.8351, 172.6454, 173.4937, 
    172.9227, 173.934, 173.3571, 173.4474, 172.9039, 169.7006, 170.3009, 
    169.6651, 169.7506, 169.7122, 169.2466, 169.0124, 168.5219, 168.6109, 
    168.9711, 169.7891, 169.511, 170.2119, 170.1961, 170.9784, 170.6254, 
    171.9432, 171.5681, 172.6533, 172.3801, 172.6405, 172.5615, 172.6415, 
    172.2408, 172.4125, 172.0601, 170.6915, 171.0931, 169.897, 169.1803, 
    168.7049, 168.3681, 168.4157, 168.5065, 168.9732, 169.4126, 169.7479, 
    169.9724, 170.1938, 170.8653, 171.221, 172.0192, 171.8749, 172.1194, 
    172.3529, 172.7455, 172.6808, 172.854, 172.1128, 172.6052, 171.7927, 
    172.0148, 170.2546, 169.586, 169.3027, 169.0546, 168.4523, 168.8681, 
    168.7041, 169.0943, 169.3426, 169.2198, 169.9786, 169.6833, 171.2421, 
    170.5697, 172.3256, 171.9045, 172.4266, 172.16, 172.617, 172.2057, 
    172.9184, 173.0739, 172.9676, 173.3757, 172.183, 172.6405, 169.2164, 
    169.2364, 169.3297, 168.9198, 168.8947, 168.5195, 168.8533, 168.9956, 
    169.357, 169.571, 169.7746, 170.2227, 170.724, 171.4263, 171.9318, 
    172.2711, 172.063, 172.2467, 172.0413, 171.9451, 173.0157, 172.4141, 
    173.317, 173.267, 172.8581, 173.2726, 169.2505, 169.1352, 168.7355, 
    169.0482, 168.4787, 168.7974, 168.9809, 169.6896, 169.8454, 169.9902, 
    170.2761, 170.6435, 171.2891, 171.8519, 172.3664, 172.3287, 172.342, 
    172.4571, 172.1721, 172.5039, 172.5597, 172.414, 173.2603, 173.0182, 
    173.2659, 173.1083, 169.1726, 169.3666, 169.2618, 169.459, 169.3201, 
    169.9383, 170.1239, 170.9937, 170.6363, 171.2052, 170.694, 170.7845, 
    171.224, 170.7215, 171.8209, 171.0753, 172.4616, 171.7157, 172.5084, 
    172.3642, 172.6029, 172.8169, 173.0862, 173.584, 173.4686, 173.8852, 
    169.656, 169.908, 169.8857, 170.1497, 170.345, 170.7688, 171.4498, 
    171.1935, 171.6641, 171.7587, 171.0437, 171.4826, 170.0768, 170.3036, 
    170.1684, 169.6759, 171.2527, 170.4425, 171.9402, 171.5, 172.7864, 
    172.1461, 173.4052, 173.9453, 174.4539, 175.0499, 170.0456, 169.8742, 
    170.181, 170.6062, 171.001, 171.5268, 171.5806, 171.6793, 171.9348, 
    172.1499, 171.7106, 172.2038, 170.3564, 171.3231, 169.8095, 170.2646, 
    170.5811, 170.4421, 171.1642, 171.3347, 172.0284, 171.6695, 173.812, 
    172.8623, 175.5041, 174.7637, 169.8144, 170.0449, 170.8489, 170.4661, 
    171.5619, 171.8323, 172.0522, 172.3337, 172.364, 172.5309, 172.2574, 
    172.5201, 171.5279, 171.9709, 170.7568, 171.0519, 170.916, 170.7672, 
    171.2269, 171.7175, 171.7278, 171.8854, 172.33, 171.5663, 173.9351, 
    172.4704, 170.2966, 170.7418, 170.8052, 170.6327, 171.8052, 171.3798, 
    172.5268, 172.2164, 172.7251, 172.4722, 172.435, 172.1105, 171.9087, 
    171.3994, 170.9855, 170.6577, 170.7338, 171.0941, 171.7475, 172.3668, 
    172.2311, 172.6864, 171.4823, 171.9867, 171.7917, 172.3004, 171.1867, 
    172.1354, 170.9448, 171.0489, 171.3714, 172.0211, 172.1648, 172.3186, 
    172.2236, 171.7641, 171.6888, 171.3635, 171.2738, 171.0262, 170.8215, 
    171.0086, 171.2053, 171.7642, 172.2689, 172.82, 172.9549, 173.6008, 
    173.0752, 173.9433, 173.2054, 174.4836, 172.1902, 173.1834, 171.386, 
    171.5791, 171.9288, 172.7321, 172.298, 172.8057, 171.6858, 171.1066, 
    170.9567, 170.6776, 170.9631, 170.9399, 171.2133, 171.1254, 171.7828, 
    171.4295, 172.4342, 172.8017, 173.8416, 174.4809, 175.1328, 175.421, 
    175.5088, 175.5455,
  257.5365, 258.4081, 258.2411, 258.9342, 258.5495, 259.0037, 257.7162, 
    258.4422, 257.9834, 257.6162, 260.2836, 258.9652, 261.6576, 260.813, 
    262.9382, 261.5261, 263.2235, 262.8972, 263.8799, 263.5981, 264.8584, 
    264.01, 265.5131, 264.6555, 264.7896, 263.9821, 259.2299, 260.1193, 
    259.1773, 259.304, 259.2471, 258.5575, 258.2106, 257.4687, 257.6049, 
    258.1495, 259.361, 258.9491, 259.9876, 259.9641, 261.1239, 260.6006, 
    262.5555, 261.9987, 263.6098, 263.204, 263.5908, 263.4734, 263.5923, 
    262.9973, 263.2521, 262.7289, 260.6985, 261.2941, 259.5209, 258.4593, 
    257.7488, 257.2331, 257.3059, 257.4449, 258.1526, 258.8033, 259.3, 
    259.6327, 259.9608, 260.9562, 261.4838, 262.6683, 262.454, 262.8169, 
    263.1636, 263.7468, 263.6507, 263.9079, 262.8072, 263.5384, 262.3321, 
    262.6617, 260.0507, 259.0602, 258.6406, 258.2732, 257.362, 257.9971, 
    257.7477, 258.332, 258.6997, 258.5178, 259.6418, 259.2044, 261.5151, 
    260.5179, 263.1232, 262.498, 263.2732, 262.8774, 263.5558, 262.9452, 
    264.0036, 264.2346, 264.0767, 264.6832, 262.9113, 263.5909, 258.5127, 
    258.5424, 258.6805, 258.0736, 258.0365, 257.465, 257.9752, 258.1858, 
    258.7209, 259.038, 259.3396, 260.0036, 260.7467, 261.7884, 262.5385, 
    263.0422, 262.7332, 263.006, 262.7011, 262.5582, 264.148, 263.2545, 
    264.5959, 264.5215, 263.914, 264.5299, 258.5632, 258.3925, 257.7958, 
    258.2638, 257.4024, 257.8906, 258.164, 259.2137, 259.4445, 259.659, 
    260.0827, 260.6273, 261.5848, 262.4199, 263.1838, 263.1277, 263.1475, 
    263.3184, 262.8953, 263.3879, 263.4708, 263.2544, 264.5115, 264.1519, 
    264.5199, 264.2857, 258.448, 258.7352, 258.58, 258.872, 258.6663, 
    259.582, 259.857, 261.1466, 260.6166, 261.4603, 260.7022, 260.8364, 
    261.4881, 260.743, 262.3739, 261.2677, 263.3251, 262.2177, 263.3946, 
    263.1805, 263.535, 263.8528, 264.253, 264.9926, 264.8212, 265.4405, 
    259.1638, 259.5372, 259.5042, 259.8953, 260.1849, 260.8131, 261.8232, 
    261.443, 262.1412, 262.2816, 261.2209, 261.8719, 259.7873, 260.1234, 
    259.9232, 259.1933, 261.5308, 260.3293, 262.5509, 261.8977, 263.8075, 
    262.8566, 264.7269, 265.5297, 266.2863, 267.1732, 259.7411, 259.4872, 
    259.9418, 260.5721, 261.1575, 261.9375, 262.0173, 262.1637, 262.543, 
    262.8623, 262.2101, 262.9424, 260.2016, 261.6352, 259.3913, 260.0657, 
    260.5349, 260.3288, 261.3995, 261.6524, 262.6819, 262.1493, 265.3315, 
    263.9202, 267.8495, 266.7472, 259.3985, 259.7401, 260.9319, 260.3643, 
    261.9896, 262.3908, 262.7172, 263.1351, 263.1801, 263.428, 263.022, 
    263.4119, 261.9392, 262.5965, 260.7953, 261.233, 261.0315, 260.8108, 
    261.4925, 262.2204, 262.2358, 262.4696, 263.1295, 261.9962, 265.5145, 
    263.338, 260.1131, 260.773, 260.8671, 260.6113, 262.3506, 261.7194, 
    263.4219, 262.961, 263.7165, 263.3409, 263.2856, 262.8038, 262.5042, 
    261.7484, 261.1345, 260.6484, 260.7613, 261.2955, 262.265, 263.1843, 
    262.9828, 263.659, 261.8715, 262.6201, 262.3306, 263.0858, 261.433, 
    262.8406, 261.0741, 261.2286, 261.7069, 262.671, 262.8844, 263.1127, 
    262.9717, 262.2896, 262.1778, 261.6952, 261.5622, 261.1949, 260.8913, 
    261.1688, 261.4604, 262.2898, 263.0389, 263.8574, 264.0579, 265.0176, 
    264.2364, 265.5266, 264.4298, 266.3304, 262.922, 264.3972, 261.7286, 
    262.0151, 262.5341, 263.7268, 263.0822, 263.8361, 262.1735, 261.3141, 
    261.0918, 260.6779, 261.1013, 261.0668, 261.4724, 261.342, 262.3174, 
    261.7931, 263.2843, 263.8301, 265.3756, 266.3265, 267.2966, 267.7258, 
    267.8565, 267.9112,
  404.2754, 405.7091, 405.43, 406.5895, 405.9458, 406.7057, 404.5656, 
    405.7663, 404.9993, 404.4041, 408.8498, 406.6413, 411.0924, 409.722, 
    413.1736, 410.8789, 413.6379, 413.107, 414.7066, 414.2477, 416.3015, 
    414.9186, 417.3701, 415.9707, 416.1893, 414.8731, 407.0846, 408.5742, 
    406.9965, 407.2085, 407.1133, 405.9591, 405.3789, 404.1659, 404.3858, 
    405.2768, 407.3039, 406.6145, 408.3539, 408.3146, 410.2264, 409.3776, 
    412.5513, 411.6465, 414.2668, 413.6062, 414.2357, 414.0447, 414.2383, 
    413.2698, 413.6844, 412.8333, 409.5364, 410.5025, 407.5718, 405.7946, 
    404.6182, 403.7856, 403.9032, 404.1275, 405.282, 406.3704, 407.2019, 
    407.7591, 408.3089, 409.9541, 410.8102, 412.7346, 412.3864, 412.9763, 
    413.5405, 414.4898, 414.3333, 414.7522, 412.9606, 414.1504, 412.1883, 
    412.724, 408.4592, 406.8003, 406.0979, 405.4836, 403.9937, 405.022, 
    404.6163, 405.5821, 406.1971, 405.8927, 407.7744, 407.0418, 410.8611, 
    409.2431, 413.4746, 412.4579, 413.7188, 413.0748, 414.1789, 413.1851, 
    414.9081, 415.2844, 415.0273, 416.0159, 413.1301, 414.2358, 405.8842, 
    405.9339, 406.165, 405.1499, 405.0879, 404.1599, 404.9854, 405.3376, 
    406.2327, 406.7632, 407.2682, 408.3806, 409.6145, 411.3048, 412.5237, 
    413.343, 412.8404, 413.2841, 412.7881, 412.5558, 415.1434, 413.6884, 
    415.8735, 415.7523, 414.7622, 415.7659, 405.9687, 405.6833, 404.694, 
    405.468, 404.0589, 404.8471, 405.3011, 407.0573, 407.444, 407.8031, 
    408.5133, 409.421, 410.9743, 412.3308, 413.5733, 413.4821, 413.5142, 
    413.7924, 413.1039, 413.9055, 414.0403, 413.6881, 415.736, 415.1498, 
    415.7497, 415.3679, 405.776, 406.2565, 405.9968, 406.4854, 406.1411, 
    407.6741, 408.1349, 410.2631, 409.4036, 410.7721, 409.5424, 409.76, 
    410.8171, 409.6086, 412.256, 410.4594, 413.8032, 412.0021, 413.9164, 
    413.5679, 414.1449, 414.6625, 415.3145, 416.5206, 416.241, 417.2517, 
    406.9738, 407.5992, 407.5439, 408.1992, 408.6846, 409.7223, 411.3615, 
    410.7442, 411.8781, 412.1061, 410.3837, 411.4405, 408.0181, 408.5814, 
    408.2458, 407.0232, 410.8865, 408.9267, 412.5439, 411.4824, 414.5887, 
    413.0408, 416.0871, 417.3972, 418.6336, 420.0843, 407.9407, 407.5154, 
    408.2772, 409.3313, 410.2809, 411.5471, 411.6768, 411.9146, 412.5311, 
    413.0503, 411.99, 413.1805, 408.7124, 411.0561, 407.3548, 408.4846, 
    409.271, 408.926, 410.6737, 411.0842, 412.7568, 411.8911, 417.0735, 
    414.7721, 421.1922, 419.3873, 407.3669, 407.9392, 409.9148, 408.9855, 
    411.6317, 412.2836, 412.8143, 413.494, 413.5674, 413.9707, 413.31, 
    413.9445, 411.5498, 412.6181, 409.6934, 410.4033, 410.0765, 409.7185, 
    410.8246, 412.0067, 412.0317, 412.4116, 413.4846, 411.6424, 417.372, 
    413.8238, 408.5642, 409.6571, 409.8098, 409.3951, 412.2182, 411.1929, 
    413.9608, 413.2108, 414.4405, 413.8289, 413.739, 412.9552, 412.468, 
    411.2399, 410.2435, 409.4552, 409.6383, 410.5048, 412.079, 413.5741, 
    413.2462, 414.3469, 411.4399, 412.6563, 412.1857, 413.4138, 410.7278, 
    413.0146, 410.1456, 410.3962, 411.1726, 412.7391, 413.0862, 413.4576, 
    413.2283, 412.119, 411.9375, 411.1536, 410.9376, 410.3416, 409.8491, 
    410.2992, 410.7724, 412.1194, 413.3375, 414.6699, 414.9966, 416.5611, 
    415.2873, 417.3919, 415.6024, 418.7053, 413.1472, 415.5494, 411.2079, 
    411.6732, 412.5164, 414.4572, 413.408, 414.6352, 411.9304, 410.5349, 
    410.1743, 409.5031, 410.1897, 410.1338, 410.7919, 410.5803, 412.1642, 
    411.3126, 413.7368, 414.6254, 417.1458, 418.6992, 420.2865, 420.9895, 
    421.2038, 421.2933,
  676.3469, 678.8848, 678.3902, 680.4385, 679.3041, 680.6378, 676.8602, 
    678.9859, 677.6277, 676.5746, 684.3205, 680.5273, 688.2945, 685.8498, 
    692.0167, 687.9133, 692.8488, 691.8975, 694.7661, 693.9424, 697.6327, 
    695.1468, 699.5576, 697.0376, 697.431, 695.0651, 681.2878, 683.8466, 
    681.1367, 681.5005, 681.3372, 679.3277, 678.2997, 676.1533, 676.5422, 
    678.1189, 681.6642, 680.4814, 683.468, 683.4004, 686.7491, 685.236, 
    690.9028, 689.2847, 693.9767, 692.792, 693.921, 693.5784, 693.9255, 
    692.1893, 692.9324, 691.4076, 685.519, 687.2416, 682.1242, 679.0361, 
    676.9532, 675.4811, 675.689, 676.0854, 678.1282, 680.0568, 681.4892, 
    682.4459, 683.3906, 686.2633, 687.7908, 691.2308, 690.6078, 691.6636, 
    692.6743, 694.3768, 694.0961, 694.8478, 691.6356, 693.7679, 690.2533, 
    691.2119, 683.6487, 680.8002, 679.5737, 678.4852, 675.8488, 677.6679, 
    676.95, 678.6597, 679.7495, 679.2101, 682.4721, 681.2144, 687.8815, 
    684.9974, 692.5563, 690.7355, 692.9938, 691.84, 693.819, 692.0375, 
    695.1279, 695.8038, 695.3419, 697.119, 691.939, 693.9211, 679.1951, 
    679.283, 679.6927, 677.8943, 677.7845, 676.1427, 677.6032, 678.2266, 
    679.8127, 680.7365, 681.6029, 683.5139, 685.6582, 688.674, 690.8534, 
    692.3204, 691.4202, 692.2148, 691.3267, 690.9109, 695.5505, 692.9393, 
    696.8629, 696.6448, 694.8658, 696.6694, 679.3447, 678.8389, 677.0875, 
    678.4576, 675.9643, 677.3583, 678.1619, 681.2409, 681.9048, 682.5215, 
    683.742, 685.3134, 688.0837, 690.5082, 692.7332, 692.5697, 692.6273, 
    693.1259, 691.892, 693.3287, 693.5704, 692.9389, 696.6157, 695.5621, 
    696.6402, 695.9539, 679.0032, 679.8549, 679.3945, 680.2599, 679.6503, 
    682.2999, 683.0915, 686.8144, 685.2824, 687.7228, 685.5297, 685.9175, 
    687.803, 685.6478, 690.3743, 687.1647, 693.1452, 689.9202, 693.3481, 
    692.7235, 693.7581, 694.6868, 695.8579, 698.0273, 697.5239, 699.3442, 
    681.0978, 682.1712, 682.0764, 683.2021, 684.0365, 685.8503, 688.7753, 
    687.673, 689.6985, 690.1063, 687.0298, 688.9163, 682.8909, 683.8589, 
    683.2822, 681.1826, 687.927, 684.4529, 690.8895, 688.9913, 694.5543, 
    691.7791, 697.2471, 699.6063, 701.8374, 704.4604, 682.7579, 682.0273, 
    683.3361, 685.1536, 686.8462, 689.1069, 689.3387, 689.7639, 690.8666, 
    691.7961, 689.8985, 692.0294, 684.0842, 688.2297, 681.7516, 683.6926, 
    685.0462, 684.4517, 687.5471, 688.28, 691.2706, 689.7219, 699.0229, 
    694.8835, 706.4677, 703.1993, 681.7725, 682.7553, 686.1935, 684.5542, 
    689.2581, 690.4238, 691.3736, 692.591, 692.7225, 693.4456, 692.2614, 
    693.3987, 689.1117, 691.0223, 685.7989, 687.0646, 686.4818, 685.8436, 
    687.8164, 689.9283, 689.9733, 690.6528, 692.5737, 689.2773, 699.5607, 
    693.1819, 683.8296, 685.7339, 686.0063, 685.2672, 690.3068, 688.4741, 
    693.4279, 692.0835, 694.2884, 693.1914, 693.0302, 691.6257, 690.7537, 
    688.558, 686.7796, 685.3743, 685.7006, 687.2457, 690.0578, 692.7346, 
    692.1469, 694.1204, 688.9153, 691.0906, 690.2487, 692.4473, 687.6438, 
    691.7318, 686.605, 687.0521, 688.4379, 691.2387, 691.8604, 692.5256, 
    692.1149, 690.1294, 689.8048, 688.4041, 688.0182, 686.9547, 686.0764, 
    686.8789, 687.7233, 690.1301, 692.3105, 694.7001, 695.2868, 698.1, 
    695.809, 699.5966, 696.3749, 701.9666, 691.9694, 696.2799, 688.5009, 
    689.3323, 690.8403, 694.3182, 692.4369, 694.6378, 689.7921, 687.2993, 
    686.6562, 685.4597, 686.6837, 686.584, 687.7582, 687.3805, 690.2102, 
    688.6879, 693.0262, 694.6203, 699.1532, 701.9557, 704.8267, 706.1004, 
    706.4888, 706.6513,
  1152.655, 1157.944, 1156.911, 1161.209, 1158.82, 1161.641, 1153.723, 
    1158.155, 1155.321, 1153.129, 1169.655, 1161.401, 1178.194, 1172.999, 
    1186.157, 1177.383, 1187.946, 1185.901, 1192.079, 1190.301, 1198.292, 
    1192.902, 1202.486, 1196.999, 1197.854, 1192.726, 1163.051, 1168.62, 
    1162.723, 1163.513, 1163.158, 1158.87, 1156.722, 1152.253, 1153.061, 
    1156.345, 1163.868, 1161.302, 1167.794, 1167.647, 1174.907, 1171.656, 
    1183.768, 1180.307, 1190.375, 1187.824, 1190.255, 1189.517, 1190.265, 
    1186.528, 1188.126, 1184.85, 1172.276, 1175.953, 1164.868, 1158.26, 
    1153.917, 1150.857, 1151.288, 1152.112, 1156.365, 1160.395, 1163.488, 
    1165.568, 1167.625, 1173.875, 1177.122, 1184.471, 1183.136, 1185.399, 
    1187.57, 1191.239, 1190.633, 1192.256, 1185.339, 1189.925, 1182.377, 
    1184.43, 1168.188, 1161.993, 1159.384, 1157.11, 1151.62, 1155.405, 
    1153.91, 1157.474, 1159.752, 1158.624, 1165.625, 1162.892, 1177.315, 
    1171.134, 1187.317, 1183.409, 1188.258, 1185.778, 1190.035, 1186.202, 
    1192.861, 1194.324, 1193.324, 1197.176, 1185.99, 1190.256, 1158.592, 
    1158.776, 1159.633, 1155.877, 1155.648, 1152.231, 1155.27, 1156.57, 
    1159.884, 1161.855, 1163.735, 1167.894, 1172.58, 1179.004, 1183.662, 
    1186.81, 1184.877, 1186.583, 1184.676, 1183.785, 1193.776, 1188.141, 
    1196.62, 1196.147, 1192.295, 1196.2, 1158.905, 1157.848, 1154.196, 
    1157.052, 1151.86, 1154.76, 1156.435, 1162.949, 1164.391, 1165.732, 
    1168.392, 1171.825, 1177.745, 1182.922, 1187.697, 1187.346, 1187.469, 
    1188.542, 1185.889, 1188.979, 1189.5, 1188.14, 1196.083, 1193.801, 
    1196.137, 1194.649, 1158.191, 1159.972, 1159.009, 1160.822, 1159.544, 
    1165.25, 1166.974, 1175.045, 1171.758, 1176.977, 1172.299, 1173.142, 
    1177.148, 1172.558, 1182.636, 1175.79, 1188.584, 1181.664, 1189.021, 
    1187.676, 1189.904, 1191.908, 1194.441, 1199.15, 1198.056, 1202.02, 
    1162.639, 1164.97, 1164.764, 1167.215, 1169.035, 1173, 1179.219, 
    1176.871, 1181.191, 1182.063, 1175.503, 1179.52, 1166.536, 1168.647, 
    1167.389, 1162.822, 1177.412, 1169.944, 1183.739, 1179.68, 1191.622, 
    1185.647, 1197.454, 1202.592, 1207.477, 1213.251, 1166.247, 1164.658, 
    1167.507, 1171.476, 1175.113, 1179.927, 1180.422, 1181.33, 1183.69, 
    1185.683, 1181.618, 1186.184, 1169.138, 1178.057, 1164.058, 1168.284, 
    1171.241, 1169.941, 1176.603, 1178.164, 1184.556, 1181.241, 1201.319, 
    1192.333, 1217.693, 1210.47, 1164.104, 1166.241, 1173.727, 1170.165, 
    1180.25, 1182.742, 1184.777, 1187.391, 1187.674, 1189.231, 1186.683, 
    1189.13, 1179.937, 1184.024, 1172.889, 1175.577, 1174.339, 1172.985, 
    1177.176, 1181.682, 1181.778, 1183.232, 1187.354, 1180.291, 1202.493, 
    1188.663, 1168.583, 1172.746, 1173.33, 1171.724, 1182.492, 1178.577, 
    1189.193, 1186.301, 1191.048, 1188.683, 1188.336, 1185.318, 1183.448, 
    1178.756, 1174.972, 1171.959, 1172.673, 1175.962, 1181.959, 1187.7, 
    1186.437, 1190.686, 1179.518, 1184.17, 1182.367, 1187.082, 1176.809, 
    1185.545, 1174.601, 1175.551, 1178.5, 1184.488, 1185.821, 1187.251, 
    1186.368, 1182.112, 1181.418, 1178.428, 1177.606, 1175.344, 1173.479, 
    1175.183, 1176.978, 1182.113, 1186.788, 1191.937, 1193.205, 1199.309, 
    1194.335, 1202.571, 1195.561, 1207.76, 1186.056, 1195.355, 1178.634, 
    1180.408, 1183.634, 1191.112, 1187.06, 1191.802, 1181.391, 1176.076, 
    1174.71, 1172.146, 1174.768, 1174.556, 1177.052, 1176.249, 1182.285, 
    1179.033, 1188.328, 1191.765, 1201.604, 1207.736, 1214.06, 1216.879, 
    1217.74, 1218.1,
  2105.699, 2120.385, 2117.501, 2129.56, 2122.839, 2130.781, 2108.646, 
    2120.976, 2113.075, 2107.006, 2153.699, 2130.104, 2179.253, 2163.429, 
    2204.022, 2176.763, 2209.558, 2203.216, 2222.352, 2216.827, 2241.925, 
    2224.92, 2255.381, 2237.816, 2240.529, 2224.368, 2134.775, 2150.71, 
    2133.845, 2136.087, 2135.08, 2122.978, 2116.974, 2104.591, 2106.819, 
    2115.923, 2137.098, 2129.823, 2148.331, 2147.907, 2169.21, 2159.509, 
    2196.521, 2185.761, 2217.056, 2209.183, 2216.684, 2214.399, 2216.714, 
    2205.191, 2210.111, 2199.911, 2161.314, 2172.396, 2139.947, 2121.27, 
    2109.182, 2100.754, 2101.938, 2104.203, 2115.977, 2127.265, 2136.017, 
    2141.945, 2147.846, 2166.082, 2175.965, 2198.722, 2194.547, 2201.636, 
    2208.406, 2219.735, 2217.855, 2222.903, 2201.447, 2215.662, 2192.183, 
    2198.594, 2149.466, 2131.776, 2124.421, 2118.054, 2102.851, 2113.308, 
    2109.163, 2119.071, 2125.455, 2122.289, 2142.108, 2134.323, 2176.556, 
    2157.99, 2207.627, 2195.402, 2210.518, 2202.827, 2216.003, 2204.163, 
    2224.792, 2229.375, 2226.239, 2238.376, 2203.496, 2216.685, 2122.2, 
    2122.716, 2125.121, 2114.62, 2113.983, 2104.53, 2112.933, 2116.549, 
    2125.827, 2131.386, 2136.719, 2148.619, 2162.203, 2181.74, 2196.19, 
    2206.073, 2199.995, 2205.364, 2199.366, 2196.576, 2227.654, 2210.157, 
    2236.615, 2235.118, 2223.023, 2235.286, 2123.078, 2120.117, 2109.955, 
    2117.893, 2103.51, 2111.518, 2116.173, 2134.486, 2138.586, 2142.416, 
    2150.052, 2160.001, 2177.875, 2193.883, 2208.794, 2207.716, 2208.095, 
    2211.393, 2203.178, 2212.739, 2214.346, 2210.155, 2234.917, 2227.732, 
    2235.086, 2230.396, 2121.078, 2126.075, 2123.37, 2128.469, 2124.872, 
    2141.037, 2145.972, 2169.632, 2159.804, 2175.522, 2161.381, 2163.863, 
    2176.044, 2162.136, 2192.99, 2171.898, 2211.521, 2189.968, 2212.868, 
    2208.73, 2215.597, 2221.818, 2229.742, 2244.662, 2241.172, 2253.877, 
    2133.606, 2140.238, 2139.65, 2146.665, 2151.907, 2163.432, 2182.406, 
    2175.198, 2188.498, 2191.205, 2171.024, 2183.333, 2144.718, 2150.788, 
    2147.166, 2134.127, 2176.853, 2154.537, 2196.432, 2183.827, 2220.927, 
    2202.415, 2239.26, 2255.725, 2271.663, 2290.879, 2143.889, 2139.346, 
    2147.504, 2158.984, 2169.838, 2184.588, 2186.118, 2188.931, 2196.279, 
    2202.53, 2189.824, 2204.108, 2152.207, 2178.83, 2137.638, 2149.741, 
    2158.3, 2154.529, 2174.379, 2179.158, 2198.989, 2188.653, 2251.618, 
    2223.143, 2305.953, 2281.574, 2137.767, 2143.872, 2165.633, 2155.178, 
    2185.585, 2193.32, 2199.682, 2207.856, 2208.724, 2213.516, 2205.679, 
    2213.204, 2184.62, 2197.322, 2163.103, 2171.25, 2167.487, 2163.389, 
    2176.132, 2190.022, 2190.321, 2194.848, 2207.741, 2185.712, 2255.403, 
    2211.764, 2150.603, 2162.687, 2164.432, 2159.708, 2192.54, 2180.429, 
    2213.398, 2204.474, 2219.143, 2211.827, 2210.759, 2201.38, 2195.523, 
    2180.98, 2169.407, 2160.39, 2162.474, 2172.423, 2190.882, 2208.803, 
    2204.903, 2218.018, 2183.327, 2197.78, 2192.152, 2206.908, 2175.008, 
    2202.095, 2168.281, 2171.169, 2180.192, 2198.775, 2202.964, 2207.425, 
    2204.687, 2191.358, 2189.202, 2179.97, 2177.448, 2170.539, 2164.881, 
    2170.049, 2175.526, 2191.363, 2206.008, 2221.908, 2225.867, 2245.167, 
    2229.409, 2255.656, 2233.269, 2272.596, 2203.702, 2232.62, 2180.605, 
    2186.075, 2196.103, 2219.343, 2206.84, 2221.488, 2189.118, 2172.77, 
    2168.612, 2160.935, 2168.788, 2168.146, 2175.752, 2173.297, 2191.896, 
    2181.832, 2210.733, 2221.371, 2252.533, 2272.518, 2293.605, 2303.17, 
    2306.114, 2307.349,
  5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 5230.692, 
    5230.692, 5230.692,
  8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 8623.953, 
    8623.953, 8623.953,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILLIQ =
  4.706965, 4.72543, 4.721836, 4.736757, 4.728476, 4.738252, 4.710704, 
    4.726165, 4.71629, 4.708624, 4.765807, 4.737423, 4.795399, 4.777212, 
    4.822982, 4.792567, 4.82913, 4.822101, 4.84327, 4.8372, 4.864346, 
    4.846074, 4.878452, 4.859977, 4.862865, 4.845472, 4.743124, 4.762268, 
    4.741992, 4.744719, 4.743495, 4.728647, 4.721178, 4.705555, 4.708388, 
    4.719863, 4.745944, 4.737079, 4.759439, 4.758934, 4.783909, 4.772637, 
    4.814741, 4.80275, 4.837453, 4.828711, 4.837042, 4.834515, 4.837075, 
    4.824258, 4.829747, 4.818477, 4.774747, 4.787573, 4.749389, 4.72653, 
    4.711382, 4.700654, 4.70217, 4.70506, 4.719931, 4.733939, 4.744634, 
    4.751797, 4.758861, 4.780293, 4.791656, 4.817169, 4.812557, 4.820371, 
    4.827841, 4.840402, 4.838333, 4.843873, 4.820163, 4.835913, 4.809931, 
    4.817029, 4.76079, 4.73947, 4.730433, 4.722527, 4.703335, 4.716583, 
    4.711358, 4.723794, 4.731709, 4.727793, 4.751993, 4.742575, 4.792331, 
    4.770857, 4.82697, 4.813503, 4.830201, 4.821675, 4.836289, 4.823135, 
    4.845935, 4.850909, 4.84751, 4.860575, 4.822407, 4.837043, 4.727684, 
    4.728323, 4.731297, 4.71823, 4.717432, 4.705478, 4.716113, 4.720647, 
    4.732168, 4.738992, 4.745485, 4.759782, 4.775784, 4.798218, 4.814375, 
    4.825226, 4.818571, 4.824447, 4.817878, 4.814802, 4.849045, 4.829798, 
    4.858694, 4.857092, 4.844005, 4.857273, 4.728771, 4.725097, 4.712359, 
    4.722326, 4.704177, 4.714331, 4.720176, 4.742773, 4.747746, 4.752362, 
    4.761487, 4.773214, 4.793833, 4.81182, 4.828276, 4.827069, 4.827494, 
    4.831175, 4.82206, 4.832673, 4.834456, 4.829795, 4.856877, 4.84913, 
    4.857058, 4.852013, 4.726291, 4.732474, 4.729132, 4.735418, 4.730989, 
    4.750704, 4.756625, 4.784395, 4.772983, 4.791151, 4.774826, 4.777717, 
    4.791748, 4.775707, 4.810828, 4.787001, 4.831318, 4.807462, 4.832816, 
    4.828205, 4.83584, 4.842687, 4.851307, 4.86724, 4.863547, 4.87689, 
    4.741701, 4.749741, 4.749031, 4.757452, 4.763686, 4.777215, 4.798969, 
    4.790781, 4.805819, 4.808842, 4.785998, 4.800016, 4.755125, 4.76236, 
    4.75805, 4.742336, 4.792669, 4.766795, 4.814643, 4.800573, 4.84171, 
    4.821225, 4.861516, 4.878808, 4.895112, 4.914216, 4.75413, 4.748664, 
    4.758453, 4.772023, 4.784632, 4.801431, 4.803151, 4.806303, 4.814474, 
    4.821351, 4.807302, 4.823076, 4.764042, 4.794919, 4.746599, 4.761117, 
    4.771222, 4.766786, 4.789845, 4.795291, 4.817463, 4.805993, 4.874538, 
    4.844135, 4.928788, 4.90504, 4.746755, 4.754111, 4.779772, 4.767551, 
    4.802553, 4.811194, 4.818226, 4.827226, 4.828197, 4.833535, 4.82479, 
    4.833189, 4.801466, 4.815626, 4.776833, 4.786257, 4.781919, 4.777166, 
    4.791847, 4.807523, 4.807856, 4.81289, 4.827098, 4.802695, 4.878475, 
    4.831589, 4.762141, 4.776349, 4.778378, 4.77287, 4.810328, 4.796733, 
    4.833405, 4.823476, 4.839751, 4.831659, 4.83047, 4.820091, 4.813637, 
    4.797357, 4.784136, 4.773668, 4.776101, 4.787604, 4.808482, 4.828286, 
    4.823944, 4.838512, 4.800009, 4.816132, 4.809896, 4.826164, 4.790564, 
    4.820875, 4.782837, 4.786164, 4.796464, 4.817228, 4.821826, 4.826743, 
    4.823708, 4.809013, 4.806607, 4.796213, 4.793347, 4.785439, 4.7789, 
    4.784875, 4.791155, 4.809018, 4.825153, 4.842784, 4.847105, 4.867774, 
    4.850947, 4.878737, 4.855108, 4.896054, 4.822632, 4.85441, 4.796932, 
    4.803103, 4.814279, 4.839971, 4.826087, 4.842325, 4.806512, 4.788002, 
    4.783218, 4.774304, 4.783422, 4.78268, 4.791414, 4.788606, 4.809612, 
    4.798321, 4.83044, 4.842196, 4.875492, 4.895975, 4.916878, 4.926125, 
    4.928941, 4.930119,
  6.780723, 6.803222, 6.798844, 6.817019, 6.806932, 6.818839, 6.785279, 
    6.804117, 6.792088, 6.782745, 6.852374, 6.81783, 6.888354, 6.866245, 
    6.921859, 6.884912, 6.929322, 6.920789, 6.946483, 6.939116, 6.972045, 
    6.949884, 6.989145, 6.966748, 6.97025, 6.949154, 6.824771, 6.848068, 
    6.823392, 6.826711, 6.825222, 6.807141, 6.798043, 6.779003, 6.782457, 
    6.796441, 6.828204, 6.81741, 6.844627, 6.844012, 6.874388, 6.860682, 
    6.911852, 6.897285, 6.939424, 6.928813, 6.938926, 6.935858, 6.938966, 
    6.923408, 6.930071, 6.916389, 6.863248, 6.878842, 6.832397, 6.804562, 
    6.786105, 6.773028, 6.774876, 6.7784, 6.796523, 6.813586, 6.826608, 
    6.835327, 6.843924, 6.869991, 6.883806, 6.914801, 6.909199, 6.918689, 
    6.927758, 6.943003, 6.940492, 6.947214, 6.918437, 6.937555, 6.90601, 
    6.91463, 6.84627, 6.820321, 6.809316, 6.799686, 6.776298, 6.792444, 
    6.786077, 6.80123, 6.810871, 6.806101, 6.835565, 6.824102, 6.884625, 
    6.858517, 6.9267, 6.910348, 6.930622, 6.920272, 6.938012, 6.922045, 
    6.949716, 6.95575, 6.951626, 6.967473, 6.921161, 6.938927, 6.805968, 
    6.806746, 6.810369, 6.794451, 6.793478, 6.778909, 6.791871, 6.797395, 
    6.811429, 6.819739, 6.827645, 6.845045, 6.864509, 6.891779, 6.911408, 
    6.924583, 6.916502, 6.923637, 6.915662, 6.911925, 6.953489, 6.930134, 
    6.965192, 6.963249, 6.947374, 6.963468, 6.807292, 6.802817, 6.787296, 
    6.799441, 6.777323, 6.789699, 6.796822, 6.824343, 6.830396, 6.836015, 
    6.847118, 6.861383, 6.886451, 6.908303, 6.928286, 6.92682, 6.927336, 
    6.931805, 6.920739, 6.933622, 6.935787, 6.93013, 6.962989, 6.953592, 
    6.963208, 6.957088, 6.804271, 6.811802, 6.807732, 6.815387, 6.809994, 
    6.833997, 6.841203, 6.874979, 6.861103, 6.883191, 6.863344, 6.866859, 
    6.883916, 6.864415, 6.907099, 6.878147, 6.931979, 6.903011, 6.933796, 
    6.928199, 6.937467, 6.945775, 6.956233, 6.975554, 6.971077, 6.987252, 
    6.823038, 6.832824, 6.831961, 6.842209, 6.849794, 6.86625, 6.892693, 
    6.882741, 6.901014, 6.904687, 6.876927, 6.893965, 6.839377, 6.848181, 
    6.842937, 6.823811, 6.885036, 6.853576, 6.911733, 6.894641, 6.94459, 
    6.919725, 6.968614, 6.989576, 7.00933, 7.032462, 6.838167, 6.831513, 
    6.843428, 6.859934, 6.875267, 6.895683, 6.897773, 6.901603, 6.911527, 
    6.919878, 6.902816, 6.921972, 6.850227, 6.88777, 6.829, 6.846669, 
    6.85896, 6.853565, 6.881604, 6.888223, 6.915158, 6.901226, 6.984401, 
    6.947533, 7.050098, 7.021353, 6.82919, 6.838143, 6.869359, 6.854496, 
    6.897047, 6.907544, 6.916084, 6.927011, 6.92819, 6.934669, 6.924054, 
    6.934249, 6.895727, 6.912926, 6.865784, 6.877242, 6.871969, 6.866189, 
    6.884037, 6.903085, 6.903489, 6.909604, 6.926856, 6.897219, 6.989172, 
    6.932307, 6.847914, 6.865196, 6.867663, 6.860965, 6.906491, 6.889976, 
    6.934511, 6.922458, 6.942213, 6.932393, 6.930948, 6.918348, 6.910511, 
    6.890733, 6.874664, 6.861936, 6.864894, 6.87888, 6.90425, 6.928298, 
    6.923027, 6.94071, 6.893956, 6.91354, 6.905968, 6.925722, 6.882478, 
    6.919301, 6.873085, 6.877129, 6.889648, 6.914872, 6.920455, 6.926425, 
    6.92274, 6.904894, 6.901972, 6.889343, 6.88586, 6.876248, 6.868298, 
    6.875562, 6.883196, 6.904901, 6.924495, 6.945893, 6.951135, 6.976201, 
    6.955796, 6.98949, 6.960844, 7.010471, 6.921434, 6.959997, 6.890217, 
    6.897715, 6.911291, 6.942479, 6.925629, 6.945336, 6.901857, 6.879364, 
    6.873548, 6.86271, 6.873796, 6.872894, 6.883511, 6.880098, 6.905622, 
    6.891905, 6.930913, 6.94518, 6.985557, 7.010375, 7.035684, 7.046875, 
    7.050283, 7.051708,
  10.29746, 10.32976, 10.32347, 10.34956, 10.33508, 10.35217, 10.304, 
    10.33104, 10.31377, 10.30036, 10.40031, 10.35072, 10.45197, 10.42023, 
    10.50007, 10.44702, 10.51078, 10.49853, 10.53543, 10.52485, 10.57213, 
    10.54031, 10.59668, 10.56452, 10.56955, 10.53926, 10.36069, 10.39413, 
    10.35871, 10.36347, 10.36133, 10.33538, 10.32232, 10.29499, 10.29995, 
    10.32002, 10.36562, 10.35012, 10.38919, 10.38831, 10.43191, 10.41224, 
    10.4857, 10.46479, 10.52529, 10.51005, 10.52457, 10.52017, 10.52463, 
    10.50229, 10.51186, 10.49222, 10.41592, 10.43831, 10.37163, 10.33168, 
    10.30519, 10.28642, 10.28907, 10.29413, 10.32014, 10.34463, 10.36332, 
    10.37584, 10.38818, 10.4256, 10.44544, 10.48993, 10.48189, 10.49552, 
    10.50854, 10.53043, 10.52682, 10.53647, 10.49516, 10.52261, 10.47731, 
    10.48969, 10.39155, 10.3543, 10.3385, 10.32468, 10.29111, 10.31428, 
    10.30514, 10.3269, 10.34073, 10.33389, 10.37618, 10.35973, 10.44661, 
    10.40913, 10.50702, 10.48354, 10.51265, 10.49779, 10.52326, 10.50034, 
    10.54007, 10.54873, 10.54281, 10.56556, 10.49907, 10.52457, 10.3337, 
    10.33481, 10.34001, 10.31716, 10.31577, 10.29486, 10.31346, 10.32139, 
    10.34154, 10.35347, 10.36481, 10.38979, 10.41773, 10.45688, 10.48506, 
    10.50398, 10.49238, 10.50262, 10.49117, 10.48581, 10.54548, 10.51195, 
    10.56229, 10.5595, 10.5367, 10.55981, 10.3356, 10.32917, 10.3069, 
    10.32433, 10.29258, 10.31034, 10.32057, 10.36007, 10.36876, 10.37683, 
    10.39277, 10.41325, 10.44923, 10.48061, 10.5093, 10.50719, 10.50793, 
    10.51435, 10.49846, 10.51696, 10.52007, 10.51194, 10.55912, 10.54563, 
    10.55944, 10.55065, 10.33126, 10.34207, 10.33623, 10.34722, 10.33948, 
    10.37393, 10.38428, 10.43276, 10.41284, 10.44455, 10.41606, 10.42111, 
    10.44559, 10.4176, 10.47888, 10.43731, 10.5146, 10.47301, 10.51721, 
    10.50917, 10.52248, 10.53441, 10.54942, 10.57717, 10.57074, 10.59397, 
    10.3582, 10.37225, 10.37101, 10.38572, 10.39661, 10.42023, 10.45819, 
    10.44391, 10.47014, 10.47541, 10.43556, 10.46002, 10.38165, 10.39429, 
    10.38677, 10.35931, 10.4472, 10.40204, 10.48553, 10.46099, 10.53271, 
    10.49701, 10.5672, 10.5973, 10.62567, 10.65889, 10.37992, 10.37037, 
    10.38747, 10.41117, 10.43318, 10.46249, 10.46549, 10.47099, 10.48524, 
    10.49722, 10.47273, 10.50023, 10.39723, 10.45113, 10.36676, 10.39212, 
    10.40977, 10.40202, 10.44228, 10.45178, 10.49045, 10.47044, 10.58987, 
    10.53693, 10.68422, 10.64294, 10.36703, 10.37988, 10.4247, 10.40336, 
    10.46445, 10.47952, 10.49178, 10.50747, 10.50916, 10.51846, 10.50322, 
    10.51786, 10.46255, 10.48724, 10.41956, 10.43601, 10.42844, 10.42015, 
    10.44577, 10.47311, 10.47369, 10.48247, 10.50724, 10.46469, 10.59672, 
    10.51507, 10.39391, 10.41872, 10.42226, 10.41265, 10.47801, 10.45429, 
    10.51824, 10.50093, 10.52929, 10.51519, 10.51312, 10.49503, 10.48378, 
    10.45538, 10.43231, 10.41404, 10.41829, 10.43836, 10.47479, 10.50931, 
    10.50175, 10.52714, 10.46001, 10.48813, 10.47725, 10.50562, 10.44353, 
    10.4964, 10.43004, 10.43585, 10.45382, 10.49004, 10.49805, 10.50662, 
    10.50133, 10.47571, 10.47152, 10.45339, 10.44839, 10.43459, 10.42317, 
    10.4336, 10.44456, 10.47572, 10.50385, 10.53458, 10.5421, 10.5781, 
    10.5488, 10.59718, 10.55604, 10.62731, 10.49946, 10.55483, 10.45464, 
    10.4654, 10.4849, 10.52968, 10.50548, 10.53378, 10.47135, 10.43906, 
    10.43071, 10.41515, 10.43107, 10.42977, 10.44501, 10.44011, 10.47676, 
    10.45706, 10.51307, 10.53355, 10.59153, 10.62717, 10.66352, 10.67959, 
    10.68449, 10.68654,
  16.38581, 16.43751, 16.42745, 16.46922, 16.44604, 16.47341, 16.39628, 
    16.43957, 16.41192, 16.39046, 16.55054, 16.47109, 16.63336, 16.58246, 
    16.71055, 16.62543, 16.72775, 16.70808, 16.76732, 16.75033, 16.82629, 
    16.77516, 16.86576, 16.81406, 16.82215, 16.77348, 16.48705, 16.54063, 
    16.48388, 16.49151, 16.48808, 16.44652, 16.42561, 16.38186, 16.3898, 
    16.42192, 16.49494, 16.47012, 16.53271, 16.5313, 16.6012, 16.56965, 
    16.68749, 16.65393, 16.75104, 16.72658, 16.74989, 16.74282, 16.74998, 
    16.71412, 16.72948, 16.69794, 16.57556, 16.61146, 16.50458, 16.44059, 
    16.39818, 16.36814, 16.37238, 16.38048, 16.42211, 16.46133, 16.49127, 
    16.51132, 16.5311, 16.59108, 16.62288, 16.69428, 16.68137, 16.70324, 
    16.72414, 16.75929, 16.7535, 16.769, 16.70266, 16.74673, 16.67403, 
    16.69389, 16.53649, 16.47681, 16.45152, 16.42938, 16.37565, 16.41274, 
    16.39811, 16.43293, 16.45509, 16.44413, 16.51187, 16.48551, 16.62477, 
    16.56467, 16.7217, 16.68402, 16.73075, 16.70689, 16.74778, 16.71098, 
    16.77477, 16.78869, 16.77918, 16.81574, 16.70894, 16.74989, 16.44382, 
    16.44561, 16.45394, 16.41735, 16.41512, 16.38165, 16.41142, 16.42412, 
    16.45637, 16.47548, 16.49365, 16.53367, 16.57846, 16.64124, 16.68646, 
    16.71683, 16.6982, 16.71465, 16.69626, 16.68765, 16.78348, 16.72962, 
    16.81047, 16.80599, 16.76937, 16.8065, 16.44686, 16.43658, 16.40091, 
    16.42882, 16.378, 16.40644, 16.4228, 16.48606, 16.49998, 16.5129, 
    16.53844, 16.57127, 16.62897, 16.67931, 16.72536, 16.72198, 16.72317, 
    16.73347, 16.70797, 16.73766, 16.74265, 16.72961, 16.80539, 16.78371, 
    16.8059, 16.79178, 16.43992, 16.45723, 16.44787, 16.46547, 16.45307, 
    16.50826, 16.52484, 16.60256, 16.57062, 16.62147, 16.57578, 16.58387, 
    16.62314, 16.57825, 16.67653, 16.60986, 16.73387, 16.66712, 16.73806, 
    16.72516, 16.74653, 16.76568, 16.7898, 16.83439, 16.82405, 16.86139, 
    16.48306, 16.50557, 16.50358, 16.52715, 16.5446, 16.58247, 16.64335, 
    16.62043, 16.66252, 16.67098, 16.60705, 16.64628, 16.52064, 16.54089, 
    16.52883, 16.48484, 16.62572, 16.5533, 16.68721, 16.64784, 16.76295, 
    16.70563, 16.81837, 16.86675, 16.91237, 16.96583, 16.51785, 16.50255, 
    16.52995, 16.56793, 16.60322, 16.65024, 16.65505, 16.66387, 16.68674, 
    16.70598, 16.66667, 16.71081, 16.5456, 16.63201, 16.49677, 16.53741, 
    16.56569, 16.55328, 16.61782, 16.63306, 16.6951, 16.663, 16.85481, 
    16.76974, 17.0066, 16.94015, 16.49721, 16.5178, 16.58962, 16.55542, 
    16.65338, 16.67756, 16.69724, 16.72242, 16.72514, 16.74008, 16.71561, 
    16.73911, 16.65034, 16.68996, 16.5814, 16.60777, 16.59563, 16.58233, 
    16.62342, 16.66729, 16.66822, 16.68231, 16.72206, 16.65377, 16.86582, 
    16.73463, 16.54028, 16.58004, 16.58572, 16.5703, 16.67513, 16.63709, 
    16.73971, 16.71193, 16.75747, 16.73483, 16.7315, 16.70246, 16.6844, 
    16.63884, 16.60184, 16.57254, 16.57935, 16.61154, 16.66997, 16.72539, 
    16.71324, 16.75401, 16.64626, 16.69138, 16.67393, 16.71945, 16.61983, 
    16.70465, 16.5982, 16.60751, 16.63634, 16.69444, 16.70731, 16.72107, 
    16.71258, 16.67146, 16.66472, 16.63564, 16.62761, 16.60548, 16.58718, 
    16.6039, 16.62148, 16.67147, 16.71662, 16.76596, 16.77805, 16.83588, 
    16.7888, 16.86656, 16.80044, 16.91501, 16.70957, 16.79849, 16.63765, 
    16.65492, 16.68619, 16.75809, 16.71924, 16.76467, 16.66446, 16.61266, 
    16.59927, 16.57432, 16.59984, 16.59776, 16.62221, 16.61435, 16.67313, 
    16.64153, 16.73142, 16.76431, 16.85748, 16.91479, 16.97327, 16.99915, 
    17.00703, 17.01032,
  26.07266, 26.16243, 26.14495, 26.21754, 26.17724, 26.22482, 26.09083, 
    26.166, 26.11799, 26.08072, 26.35905, 26.22079, 26.50347, 26.41468, 
    26.63831, 26.48964, 26.6684, 26.634, 26.73765, 26.70791, 26.84098, 
    26.75138, 26.91022, 26.81955, 26.83371, 26.74844, 26.24854, 26.3418, 
    26.24303, 26.2563, 26.25034, 26.17808, 26.14175, 26.06581, 26.07958, 
    26.13536, 26.26227, 26.21911, 26.32802, 26.32555, 26.44736, 26.39237, 
    26.598, 26.53938, 26.70915, 26.66635, 26.70714, 26.69476, 26.7073, 
    26.64455, 26.67142, 26.61627, 26.40266, 26.46525, 26.27905, 26.16778, 
    26.09413, 26.042, 26.04936, 26.06341, 26.13568, 26.20383, 26.25589, 
    26.29078, 26.3252, 26.42971, 26.48519, 26.60987, 26.58732, 26.62554, 
    26.66209, 26.72359, 26.71346, 26.7406, 26.62452, 26.70161, 26.57448, 
    26.60919, 26.3346, 26.23075, 26.18677, 26.14831, 26.05503, 26.11941, 
    26.09401, 26.15447, 26.19298, 26.17393, 26.29173, 26.24586, 26.48848, 
    26.38368, 26.65782, 26.59194, 26.67364, 26.63192, 26.70345, 26.63906, 
    26.7507, 26.77508, 26.75842, 26.82248, 26.6355, 26.70714, 26.17339, 
    26.1765, 26.19097, 26.12742, 26.12353, 26.06543, 26.11712, 26.13917, 
    26.19521, 26.22842, 26.26004, 26.32969, 26.40772, 26.51723, 26.59621, 
    26.64929, 26.61673, 26.64548, 26.61334, 26.59829, 26.76595, 26.67167, 
    26.81325, 26.8054, 26.74124, 26.80628, 26.17868, 26.16081, 26.09888, 
    26.14733, 26.05911, 26.10846, 26.13688, 26.24683, 26.27105, 26.29353, 
    26.33799, 26.39518, 26.49582, 26.58371, 26.66422, 26.65831, 26.66039, 
    26.67841, 26.6338, 26.68574, 26.69447, 26.67165, 26.80434, 26.76636, 
    26.80523, 26.78049, 26.16662, 26.1967, 26.18044, 26.21103, 26.18948, 
    26.28545, 26.3143, 26.44973, 26.39405, 26.48272, 26.40304, 26.41714, 
    26.48563, 26.40734, 26.57886, 26.46246, 26.67911, 26.56241, 26.68644, 
    26.66387, 26.70125, 26.73479, 26.77703, 26.85518, 26.83706, 26.90255, 
    26.24161, 26.28076, 26.27731, 26.31833, 26.34872, 26.4147, 26.52091, 
    26.48091, 26.55438, 26.56915, 26.45756, 26.52602, 26.30699, 26.34225, 
    26.32125, 26.2447, 26.49013, 26.36387, 26.59752, 26.52874, 26.73, 
    26.62971, 26.82709, 26.91197, 26.99209, 27.08608, 26.30215, 26.27552, 
    26.32321, 26.38937, 26.45089, 26.53293, 26.54134, 26.55674, 26.59669, 
    26.63033, 26.56162, 26.63877, 26.35045, 26.50112, 26.26546, 26.33619, 
    26.38546, 26.36383, 26.47634, 26.50294, 26.61131, 26.55523, 26.891, 
    26.74188, 27.15787, 27.04092, 26.26622, 26.30205, 26.42717, 26.36756, 
    26.53841, 26.58066, 26.61504, 26.65908, 26.66383, 26.68996, 26.64716, 
    26.68827, 26.53311, 26.60233, 26.41283, 26.45882, 26.43765, 26.41446, 
    26.48612, 26.56271, 26.56433, 26.58895, 26.65845, 26.53911, 26.91033, 
    26.68044, 26.34118, 26.41047, 26.42037, 26.3935, 26.57642, 26.50998, 
    26.68933, 26.64073, 26.7204, 26.68078, 26.67496, 26.62417, 26.5926, 
    26.51303, 26.44847, 26.39739, 26.40926, 26.4654, 26.5674, 26.66427, 
    26.64302, 26.71434, 26.52599, 26.6048, 26.57431, 26.65388, 26.47985, 
    26.628, 26.44213, 26.45837, 26.50867, 26.61016, 26.63265, 26.65671, 
    26.64186, 26.56999, 26.55823, 26.50744, 26.49344, 26.45483, 26.42292, 
    26.45208, 26.48274, 26.57001, 26.64894, 26.73527, 26.75643, 26.8578, 
    26.77527, 26.91162, 26.79567, 26.99672, 26.6366, 26.79224, 26.51096, 
    26.5411, 26.59574, 26.72148, 26.65351, 26.73302, 26.55777, 26.46734, 
    26.44399, 26.4005, 26.44499, 26.44136, 26.484, 26.47029, 26.57292, 
    26.51774, 26.67481, 26.73238, 26.89568, 26.99633, 27.09919, 27.14474, 
    27.15862, 27.16442,
  44.5972, 44.76147, 44.72947, 44.8625, 44.78862, 44.87584, 44.63042, 
    44.76802, 44.6801, 44.61194, 45.12241, 44.86844, 45.38848, 45.2248, 
    45.6377, 45.36296, 45.69341, 45.62972, 45.82178, 45.76663, 46.01371, 
    45.84727, 46.14259, 45.97387, 46.0002, 45.8418, 44.91936, 45.09068, 
    44.90924, 44.93361, 44.92267, 44.79015, 44.72361, 44.58467, 44.60984, 
    44.7119, 44.94456, 44.86537, 45.06534, 45.06081, 45.28502, 45.18371, 
    45.56312, 45.45478, 45.76893, 45.68961, 45.7652, 45.74226, 45.7655, 
    45.64926, 45.69901, 45.59692, 45.20266, 45.31799, 44.97536, 44.77127, 
    44.63645, 44.54116, 44.55461, 44.58028, 44.7125, 44.83735, 44.93285, 
    44.9969, 45.06015, 45.25249, 45.35476, 45.58508, 45.54337, 45.61406, 
    45.68173, 45.79572, 45.77692, 45.82726, 45.61218, 45.75495, 45.51964, 
    45.58381, 45.07743, 44.88671, 44.80607, 44.73562, 44.56496, 44.68271, 
    44.63624, 44.74691, 44.81745, 44.78254, 44.99866, 44.91445, 45.36083, 
    45.16773, 45.67383, 45.55193, 45.70312, 45.62587, 45.75837, 45.63909, 
    45.84601, 45.89126, 45.86033, 45.97931, 45.6325, 45.76521, 44.78156, 
    44.78725, 44.81378, 44.69736, 44.69025, 44.58398, 44.67852, 44.71888, 
    44.82154, 44.88245, 44.94046, 45.06841, 45.21198, 45.41389, 45.55981, 
    45.65803, 45.59776, 45.65097, 45.5915, 45.56366, 45.8743, 45.69947, 
    45.96217, 45.94757, 45.82846, 45.94921, 44.79125, 44.75851, 44.64514, 
    44.73383, 44.57243, 44.66267, 44.71469, 44.91622, 44.96067, 45.00196, 
    45.08368, 45.18889, 45.37437, 45.5367, 45.68567, 45.67473, 45.67858, 
    45.71196, 45.62935, 45.72554, 45.74173, 45.69945, 45.94562, 45.87508, 
    45.94726, 45.90131, 44.76915, 44.82428, 44.79448, 44.85054, 44.81104, 
    44.98713, 45.04013, 45.28939, 45.18682, 45.35021, 45.20337, 45.22934, 
    45.35558, 45.21128, 45.52774, 45.31284, 45.71326, 45.49733, 45.72684, 
    45.68502, 45.75429, 45.81647, 45.89488, 46.04013, 46.00643, 46.1283, 
    44.90665, 44.97851, 44.97216, 45.04753, 45.1034, 45.22484, 45.42067, 
    45.34687, 45.48249, 45.50979, 45.30381, 45.43012, 45.02669, 45.09151, 
    45.05289, 44.91232, 45.36388, 45.13128, 45.56223, 45.43514, 45.8076, 
    45.62179, 45.9879, 46.14585, 46.29523, 46.47085, 45.01779, 44.96888, 
    45.0565, 45.17819, 45.29152, 45.44288, 45.4584, 45.48686, 45.5607, 
    45.62293, 45.49588, 45.63855, 45.10659, 45.38415, 44.95042, 45.08037, 
    45.171, 45.1312, 45.33845, 45.38751, 45.58774, 45.48406, 46.10679, 
    45.82964, 46.60524, 46.38642, 44.95181, 45.01762, 45.24781, 45.13806, 
    45.453, 45.53105, 45.59464, 45.67615, 45.68496, 45.73337, 45.65408, 
    45.73023, 45.4432, 45.57112, 45.2214, 45.30614, 45.26712, 45.22439, 
    45.35648, 45.49788, 45.50089, 45.54638, 45.67499, 45.45428, 46.14279, 
    45.71571, 45.08954, 45.21705, 45.23528, 45.1858, 45.52322, 45.40051, 
    45.73219, 45.64217, 45.7898, 45.71635, 45.70556, 45.61153, 45.55313, 
    45.40613, 45.28706, 45.19297, 45.21482, 45.31827, 45.50655, 45.68576, 
    45.64642, 45.77855, 45.43005, 45.5757, 45.51933, 45.66653, 45.34492, 
    45.61862, 45.27537, 45.30531, 45.39808, 45.58561, 45.62723, 45.67178, 
    45.64428, 45.51134, 45.4896, 45.39582, 45.36999, 45.29878, 45.23997, 
    45.2937, 45.35025, 45.51139, 45.65737, 45.81736, 45.85664, 46.045, 
    45.89161, 46.1452, 45.9295, 46.30387, 45.63453, 45.92314, 45.40231, 
    45.45797, 45.55894, 45.7918, 45.66584, 45.81319, 45.48875, 45.32185, 
    45.2788, 45.19868, 45.28064, 45.27396, 45.35258, 45.32729, 45.51675, 
    45.41483, 45.7053, 45.81202, 46.11551, 46.30315, 46.49537, 46.58065, 
    46.60666, 46.61754,
  75.10475, 75.4586, 75.38952, 75.67706, 75.51723, 75.70596, 75.17618, 
    75.47274, 75.28311, 75.13644, 76.24215, 75.68993, 76.82531, 76.466, 
    77.37594, 76.76917, 77.49962, 77.35824, 77.78547, 77.66251, 78.21509, 
    77.84237, 78.5051, 78.12567, 78.18476, 77.83015, 75.80031, 76.17292, 
    75.77837, 75.83121, 75.80749, 75.52055, 75.37688, 75.07783, 75.13192, 
    75.35164, 75.855, 75.68327, 76.11768, 76.10781, 76.59796, 76.37608, 
    77.21069, 76.97136, 77.66764, 77.49117, 77.65934, 77.60825, 77.66, 
    77.40157, 77.51205, 77.28553, 76.41753, 76.67033, 75.92191, 75.47976, 
    75.18914, 74.98443, 75.01329, 75.0684, 75.35293, 75.6226, 75.82957, 
    75.96873, 76.10639, 76.52664, 76.75113, 77.25932, 77.167, 77.32351, 
    77.47367, 77.72734, 77.68545, 77.79769, 77.31935, 77.63651, 77.11454, 
    77.2565, 76.14404, 75.72952, 75.55495, 75.40279, 75.03551, 75.28873, 
    75.18868, 75.42715, 75.57957, 75.50409, 75.97253, 75.78966, 76.76448, 
    76.34114, 77.45612, 77.18593, 77.5212, 77.34969, 77.64411, 77.37902, 
    77.83955, 77.94069, 77.87154, 78.13789, 77.36439, 77.65935, 75.50198, 
    75.51428, 75.57162, 75.3203, 75.30499, 75.07635, 75.2797, 75.36668, 
    75.58841, 75.72028, 75.84609, 76.12437, 76.43791, 76.88125, 77.20338, 
    77.42105, 77.2874, 77.40536, 77.27352, 77.2119, 77.90276, 77.51309, 
    78.09945, 78.06673, 77.80037, 78.07042, 75.52292, 75.4522, 75.20783, 
    75.39893, 75.05154, 75.24557, 75.35764, 75.7935, 75.88998, 75.97973, 
    76.15766, 76.38741, 76.79425, 77.15226, 77.48242, 77.45811, 77.46667, 
    77.54086, 77.35742, 77.57106, 77.60706, 77.51303, 78.06236, 77.90449, 
    78.06604, 77.96315, 75.47517, 75.59432, 75.52988, 75.65117, 75.56569, 
    75.94746, 76.06277, 76.60755, 76.38287, 76.74112, 76.41908, 76.47593, 
    76.75292, 76.43639, 77.13245, 76.65903, 77.54374, 77.06526, 77.57395, 
    77.48099, 77.63504, 77.77363, 77.94878, 78.27444, 78.19874, 78.47289, 
    75.77273, 75.92873, 75.91495, 76.0789, 76.20066, 76.46607, 76.89619, 
    76.7338, 77.03249, 77.09279, 76.63921, 76.917, 76.03352, 76.17474, 
    76.09057, 75.78503, 76.77118, 76.26151, 77.20873, 76.92806, 77.75384, 
    77.34065, 78.15714, 78.51244, 78.85021, 79.24949, 76.01415, 75.90781, 
    76.09844, 76.36401, 76.61223, 76.94511, 76.97935, 77.04215, 77.20534, 
    77.34318, 77.06206, 77.37782, 76.20762, 76.81577, 75.86771, 76.15044, 
    76.34829, 76.26133, 76.71528, 76.82317, 77.26521, 77.03596, 78.42442, 
    77.80302, 79.55668, 79.05722, 75.87074, 76.01378, 76.5164, 76.27631, 
    76.96745, 77.13977, 77.28049, 77.46128, 77.48083, 77.58848, 77.41228, 
    77.58149, 76.94583, 77.2284, 76.45854, 76.64433, 76.55872, 76.46509, 
    76.75491, 77.06647, 77.07312, 77.17366, 77.4587, 76.97027, 78.50556, 
    77.54919, 76.17045, 76.44902, 76.48895, 76.38065, 77.12245, 76.85178, 
    77.58584, 77.38586, 77.71414, 77.55061, 77.52663, 77.31789, 77.18861, 
    76.86416, 76.60245, 76.39633, 76.44414, 76.67094, 77.08561, 77.48263, 
    77.39526, 77.68908, 76.91685, 77.23853, 77.11385, 77.43991, 76.7295, 
    77.33363, 76.57681, 76.64249, 76.84644, 77.26048, 77.35272, 77.45156, 
    77.39053, 77.0962, 77.0482, 76.84145, 76.78461, 76.62817, 76.49922, 
    76.61703, 76.7412, 77.09631, 77.41959, 77.77561, 77.8633, 78.28538, 
    77.94145, 78.51097, 78.02625, 78.86981, 77.3689, 78.01201, 76.85573, 
    76.97839, 77.20144, 77.7186, 77.43837, 77.7663, 77.04633, 76.67882, 
    76.58434, 76.40883, 76.58836, 76.57372, 76.74633, 76.69076, 77.10816, 
    76.88331, 77.52603, 77.76369, 78.44407, 78.86816, 79.30544, 79.50036, 
    79.55991, 79.58485,
  138.2295, 139.2781, 139.0721, 139.9332, 139.4533, 140.0204, 138.4399, 
    139.3203, 138.7561, 138.3228, 141.6568, 139.972, 143.4813, 142.3514, 
    145.2499, 143.3036, 145.6535, 145.1923, 146.5958, 146.1889, 148.0374, 
    146.785, 149.0286, 147.7348, 147.9347, 146.7443, 140.3055, 141.4433, 
    140.2391, 140.3992, 140.3273, 139.4632, 139.0345, 138.1504, 138.3095, 
    138.9595, 140.4714, 139.952, 141.2735, 141.2432, 142.7643, 142.0716, 
    144.7143, 143.946, 146.2058, 145.6259, 146.1784, 146.0101, 146.1806, 
    145.3333, 145.6942, 144.9563, 142.2004, 142.9917, 140.6748, 139.3413, 
    138.4782, 137.8764, 137.961, 138.1226, 138.9633, 139.7693, 140.3942, 
    140.8175, 141.2388, 142.5409, 143.2465, 144.8714, 144.5734, 145.0795, 
    145.5686, 146.4031, 146.2646, 146.6364, 145.066, 146.1031, 144.4046, 
    144.8623, 141.3545, 140.0914, 139.5663, 139.1116, 138.0261, 138.7728, 
    138.4768, 139.1842, 139.6401, 139.414, 140.8291, 140.2733, 143.2887, 
    141.9631, 145.5113, 144.6344, 145.7242, 145.1645, 146.1282, 145.2599, 
    146.7756, 147.1131, 146.8822, 147.7761, 145.2123, 146.1784, 139.4077, 
    139.4445, 139.6163, 138.8664, 138.821, 138.146, 138.746, 139.0042, 
    139.6666, 140.0636, 140.4444, 141.294, 142.2639, 143.6589, 144.6907, 
    145.3968, 144.9624, 145.3457, 144.9174, 144.7182, 146.9863, 145.6976, 
    147.6463, 147.5361, 146.6453, 147.5485, 139.4703, 139.259, 138.5334, 
    139.1001, 138.0732, 138.645, 138.9773, 140.2849, 140.5777, 140.8511, 
    141.3963, 142.1067, 143.3829, 144.5259, 145.5972, 145.5178, 145.5457, 
    145.7886, 145.1896, 145.8878, 146.0062, 145.6974, 147.5213, 146.9921, 
    147.5338, 147.1883, 139.3275, 139.6844, 139.4912, 139.8553, 139.5985, 
    140.7527, 141.105, 142.7944, 142.0927, 143.2149, 142.2053, 142.3824, 
    143.2522, 142.2592, 144.4621, 142.9561, 145.7981, 144.2464, 145.8973, 
    145.5925, 146.0983, 146.5565, 147.1402, 148.2391, 147.982, 148.9178, 
    140.2221, 140.6956, 140.6536, 141.1545, 141.5288, 142.3517, 143.7064, 
    143.1918, 144.1414, 144.3347, 142.8938, 143.7727, 141.0155, 141.4489, 
    141.1903, 140.2593, 143.3099, 141.7166, 144.7079, 143.8079, 146.4909, 
    145.1351, 147.8412, 149.0539, 150.2278, 151.6432, 140.9563, 140.6319, 
    141.2144, 142.0341, 142.8091, 143.8622, 143.9715, 144.1723, 144.697, 
    145.1433, 144.2361, 145.256, 141.5502, 143.4511, 140.51, 141.3741, 
    141.9853, 141.716, 143.1333, 143.4745, 144.8905, 144.1525, 148.7514, 
    146.6541, 152.7535, 150.9578, 140.5192, 140.9551, 142.5088, 141.7623, 
    143.9335, 144.4857, 144.94, 145.5281, 145.5921, 145.945, 145.3682, 
    145.922, 143.8645, 144.7715, 142.3282, 142.9099, 142.6413, 142.3486, 
    143.2585, 144.2503, 144.2716, 144.5948, 145.5197, 143.9425, 149.0302, 
    145.816, 141.4357, 142.2985, 142.4231, 142.0857, 144.43, 143.5653, 
    145.9364, 145.2821, 146.3595, 145.8207, 145.742, 145.0612, 144.643, 
    143.6046, 142.7783, 142.1345, 142.2833, 142.9937, 144.3117, 145.5979, 
    145.3128, 146.2766, 143.7722, 144.8042, 144.4023, 145.4583, 143.1782, 
    145.1123, 142.6979, 142.9041, 143.5483, 144.8752, 145.1743, 145.4964, 
    145.2973, 144.3456, 144.1917, 143.5325, 143.3524, 142.8591, 142.4551, 
    142.8241, 143.2152, 144.346, 145.392, 146.5631, 146.8547, 148.2763, 
    147.1156, 149.0488, 147.3999, 150.2966, 145.227, 147.3521, 143.5779, 
    143.9684, 144.6844, 146.3742, 145.4533, 146.5322, 144.1857, 143.0184, 
    142.7215, 142.1734, 142.7341, 142.6882, 143.2314, 143.0561, 144.3841, 
    143.6655, 145.74, 146.5235, 148.8188, 150.2908, 151.844, 152.5485, 
    152.7653, 152.8563,
  366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466,
  603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILPSI =
  -0.01747912, -0.01720452, -0.01725754, -0.01703871, -0.01715974, 
    -0.01701698, -0.01742308, -0.0171937, -0.01733976, -0.01745422, 
    -0.01662254, -0.01702903, -0.01621154, -0.01646261, -0.0158398, 
    -0.01625032, -0.0157584, -0.01585151, -0.01557314, -0.01565234, 
    -0.01530204, -0.01553674, -0.01512387, -0.01535775, -0.0153209, 
    -0.01554454, -0.01694639, -0.01667256, -0.01696276, -0.01692338, 
    -0.01694104, -0.01715722, -0.01726727, -0.01750032, -0.01745776, 
    -0.01728673, -0.0169057, -0.01703403, -0.01671267, -0.01671985, 
    -0.01636961, -0.01652653, -0.01594974, -0.01611142, -0.01564903, 
    -0.01576394, -0.0156544, -0.01568753, -0.01565397, -0.01582287, 
    -0.01575026, -0.01589978, -0.01649701, -0.01631899, -0.01685617, 
    -0.01718833, -0.01741294, -0.01757423, -0.01755133, -0.01750776, 
    -0.01728573, -0.01707978, -0.01692461, -0.01682166, -0.01672089, 
    -0.01641975, -0.01626281, -0.01591725, -0.01597904, -0.01587453, 
    -0.01577542, -0.0156105, -0.01563752, -0.01556531, -0.0158773, 
    -0.01566919, -0.01601435, -0.01591913, -0.0166935, -0.01699931, 
    -0.01713104, -0.01724733, -0.01753374, -0.0173354, -0.0174133, 
    -0.01722862, -0.01711236, -0.01716976, -0.01681885, -0.01695434, 
    -0.01625356, -0.01655148, -0.01578695, -0.01596634, -0.01574428, 
    -0.01585717, -0.01566426, -0.01583776, -0.01553854, -0.01547419, 
    -0.01551813, -0.01535012, -0.01584744, -0.01565439, -0.01717136, 
    -0.01716199, -0.01711839, -0.01731094, -0.0173228, -0.01750148, 
    -0.01734241, -0.01727513, -0.01710566, -0.01700624, -0.01691232, 
    -0.0167078, -0.01648253, -0.01617306, -0.01595464, -0.01581003, 
    -0.01589854, -0.01582037, -0.01590778, -0.01594893, -0.01549826, 
    -0.01574958, -0.01537416, -0.01539468, -0.0155636, -0.01539237, 
    -0.01715541, -0.01720942, -0.01739834, -0.0172503, -0.01752106, 
    -0.01736893, -0.01728209, -0.01695147, -0.01687978, -0.01681356, 
    -0.01668363, -0.01651846, -0.01623297, -0.01598895, -0.01576968, 
    -0.01578563, -0.01578001, -0.01573144, -0.01585205, -0.01571173, 
    -0.0156883, -0.01574962, -0.01539743, -0.01549717, -0.01539512, 
    -0.01545997, -0.01719185, -0.01710118, -0.0171501, -0.01705822, 
    -0.01712289, -0.01683731, -0.0167527, -0.01636288, -0.01652169, 
    -0.01626976, -0.01649591, -0.01645558, -0.01626157, -0.01648361, 
    -0.01600228, -0.01632687, -0.01572955, -0.01604764, -0.01570985, 
    -0.01577062, -0.01567014, -0.01558074, -0.01546907, -0.01526527, 
    -0.0153122, -0.01514347, -0.01696698, -0.01685113, -0.01686131, 
    -0.01674093, -0.01665249, -0.01646256, -0.01616282, -0.01627484, 
    -0.01606985, -0.01602903, -0.01634073, -0.01614856, -0.01677409, 
    -0.01667125, -0.01673241, -0.0169578, -0.01624892, -0.01660861, 
    -0.01595106, -0.01614099, -0.01559345, -0.01586316, -0.0153381, 
    -0.0151194, -0.01491676, -0.01468361, -0.01678828, -0.01686659, 
    -0.01672668, -0.01653514, -0.0163596, -0.01612933, -0.01610598, 
    -0.0160633, -0.01595333, -0.01586149, -0.01604981, -0.01583856, 
    -0.01664746, -0.01621811, -0.01689628, -0.01668886, -0.01654637, 
    -0.01660873, -0.0162877, -0.01621301, -0.01591332, -0.0160675, 
    -0.01517305, -0.0155619, -0.01450882, -0.01479503, -0.01689403, 
    -0.01678856, -0.01642698, -0.01659796, -0.0161141, -0.01599735, 
    -0.01590314, -0.01578356, -0.01577072, -0.01570039, -0.01581581, 
    -0.01570494, -0.01612885, -0.01593789, -0.0164679, -0.01633715, 
    -0.01639717, -0.01646326, -0.0162602, -0.01604682, -0.01604233, 
    -0.01597457, -0.01578525, -0.01611217, -0.01512359, -0.01572599, 
    -0.01667436, -0.01647465, -0.01644637, -0.01652327, -0.01600901, 
    -0.01619331, -0.01570211, -0.01583325, -0.015619, -0.01572506, 
    -0.01574073, -0.01587826, -0.01596454, -0.0161848, -0.01636646, 
    -0.0165121, -0.01647811, -0.01631856, -0.01603387, -0.01576954, 
    -0.01582703, -0.01563517, -0.01614866, -0.01593113, -0.01601481, 
    -0.01579761, -0.01627782, -0.01586782, -0.01638445, -0.01633843, 
    -0.01619699, -0.01591647, -0.01585517, -0.01578994, -0.01583016, 
    -0.01602672, -0.01605919, -0.01620042, -0.01623963, -0.01634844, 
    -0.01643911, -0.01635624, -0.0162697, -0.01602665, -0.01581099, 
    -0.01557946, -0.01552338, -0.01525851, -0.01547371, -0.0151203, 
    -0.01542014, -0.01490515, -0.01584445, -0.01542911, -0.01619059, 
    -0.01610663, -0.01595594, -0.01561613, -0.01579862, -0.01558544, 
    -0.01606047, -0.01631307, -0.01637917, -0.0165032, -0.01637634, 
    -0.01638662, -0.01626614, -0.01630476, -0.01601865, -0.01617165, 
    -0.01574112, -0.01558712, -0.01516105, -0.01490613, -0.01465149, 
    -0.01454057, -0.014507, -0.01449298,
  -0.02241809, -0.0220693, -0.02213665, -0.02185867, -0.02201241, 
    -0.02183107, -0.02234691, -0.02205556, -0.02224108, -0.02238647, 
    -0.02132993, -0.02184637, -0.02080766, -0.02112672, -0.0203352, 
    -0.02085695, -0.02023173, -0.02035008, -0.01999623, -0.02009691, 
    -0.01965156, -0.01994994, -0.01942501, -0.01972239, -0.01967553, 
    -0.01995987, -0.02174139, -0.02139349, -0.02176219, -0.02171215, 
    -0.0217346, -0.02200921, -0.02214901, -0.02244502, -0.02239097, 
    -0.02217372, -0.02168969, -0.02185273, -0.02144445, -0.02145357, 
    -0.02100854, -0.02120794, -0.02047494, -0.02068043, -0.0200927, 
    -0.02023877, -0.02009953, -0.02014164, -0.02009898, -0.02031368, 
    -0.02022138, -0.02041144, -0.02117043, -0.02094422, -0.02162677, 
    -0.02204874, -0.02233404, -0.02253889, -0.02250981, -0.02245447, 
    -0.02217246, -0.02191084, -0.02171371, -0.02158292, -0.02145489, 
    -0.02107226, -0.02087283, -0.02043364, -0.02051218, -0.02037934, 
    -0.02025336, -0.02004372, -0.02007806, -0.01998627, -0.02038286, 
    -0.02011833, -0.02055706, -0.02043603, -0.0214201, -0.02180862, 
    -0.02197596, -0.02212368, -0.02248747, -0.02223555, -0.02233449, 
    -0.02209991, -0.02195223, -0.02202514, -0.02157935, -0.02175148, 
    -0.02086107, -0.02123965, -0.02026801, -0.02049603, -0.02021378, 
    -0.02035728, -0.02011206, -0.02033261, -0.01995224, -0.01987044, 
    -0.01992629, -0.01971269, -0.02034491, -0.02009952, -0.02202718, 
    -0.02201527, -0.02195989, -0.02220448, -0.02221955, -0.0224465, 
    -0.02224445, -0.02215899, -0.02194371, -0.02181742, -0.02169811, 
    -0.02143826, -0.02115203, -0.02075876, -0.02048117, -0.02029735, 
    -0.02040986, -0.02031049, -0.0204216, -0.02047391, -0.01990104, 
    -0.02022052, -0.01974326, -0.01976934, -0.01998409, -0.0197664, 
    -0.02200691, -0.02207552, -0.02231549, -0.02212746, -0.02247137, 
    -0.02227814, -0.02216784, -0.02174784, -0.02165676, -0.02157263, 
    -0.02140755, -0.02119768, -0.0208349, -0.02052477, -0.02024606, 
    -0.02026635, -0.0202592, -0.02019745, -0.02035077, -0.0201724, 
    -0.02014262, -0.02022057, -0.01977284, -0.01989964, -0.0197699, 
    -0.01985235, -0.0220532, -0.02193802, -0.02200017, -0.02188345, 
    -0.0219656, -0.02160281, -0.02149531, -0.02099999, -0.02120178, 
    -0.02088165, -0.02116903, -0.02111779, -0.02087124, -0.0211534, 
    -0.02054172, -0.02095423, -0.02019506, -0.02059937, -0.02017001, 
    -0.02024726, -0.02011954, -0.02000588, -0.01986391, -0.01960481, 
    -0.01966448, -0.01944993, -0.02176754, -0.02162036, -0.0216333, 
    -0.02148035, -0.02136798, -0.02112666, -0.02074574, -0.02088811, 
    -0.02062759, -0.02057571, -0.02097184, -0.02072763, -0.02152248, 
    -0.02139182, -0.02146953, -0.02175587, -0.02085518, -0.02131223, 
    -0.02047661, -0.02071801, -0.02002204, -0.02036489, -0.01969741, 
    -0.01941933, -0.01916164, -0.01886511, -0.02154052, -0.02164, 
    -0.02146224, -0.02121888, -0.02099583, -0.02070319, -0.02067351, 
    -0.02061927, -0.02047949, -0.02036277, -0.02060212, -0.02033362, 
    -0.0213616, -0.02081602, -0.02167772, -0.0214142, -0.02123315, 
    -0.02131239, -0.02090445, -0.02080954, -0.02042865, -0.0206246, 
    -0.01948754, -0.01998194, -0.01864277, -0.01900682, -0.02167487, 
    -0.02154087, -0.02108144, -0.0212987, -0.02068383, -0.02053545, 
    -0.0204157, -0.0202637, -0.02024738, -0.02015799, -0.0203047, 
    -0.02016377, -0.02070257, -0.02045988, -0.02113344, -0.02096729, 
    -0.02104356, -0.02112754, -0.0208695, -0.02059832, -0.02059261, 
    -0.02050649, -0.02026585, -0.02068138, -0.01942465, -0.02019053, 
    -0.02139577, -0.02114201, -0.02110608, -0.0212038, -0.02055027, 
    -0.02078449, -0.02016017, -0.02032687, -0.02005452, -0.02018935, 
    -0.02020927, -0.02038409, -0.02049375, -0.02077368, -0.02100454, 
    -0.0211896, -0.02114642, -0.02094367, -0.02058187, -0.02024589, 
    -0.02031897, -0.02007508, -0.02072775, -0.02045128, -0.02055765, 
    -0.02028156, -0.0208919, -0.02037081, -0.0210274, -0.02096892, 
    -0.02078917, -0.02043265, -0.02035473, -0.02027182, -0.02032295, 
    -0.02057278, -0.02061405, -0.02079353, -0.02084337, -0.02098164, 
    -0.02109686, -0.02099155, -0.02088157, -0.02057269, -0.02029858, 
    -0.02000427, -0.01993297, -0.01959621, -0.01986982, -0.01942047, 
    -0.01980171, -0.01914688, -0.02034111, -0.01981311, -0.02078105, 
    -0.02067434, -0.02048281, -0.02005088, -0.02028286, -0.02001186, 
    -0.02061567, -0.0209367, -0.02102069, -0.02117829, -0.0210171, 
    -0.02103016, -0.02087706, -0.02092613, -0.02056252, -0.02075697, 
    -0.02020976, -0.020014, -0.01947229, -0.01914812, -0.01882425, 
    -0.01868317, -0.01864046, -0.01862263,
  -0.02349889, -0.02313164, -0.02320256, -0.02290984, -0.02307174, 
    -0.02288077, -0.02342395, -0.02311717, -0.02331252, -0.02346559, 
    -0.02235299, -0.02289688, -0.02180281, -0.02213893, -0.021305, 
    -0.02185474, -0.02119597, -0.02132069, -0.02094778, -0.02105389, 
    -0.02058451, -0.02089901, -0.02034569, -0.02065917, -0.02060977, 
    -0.02090946, -0.02278633, -0.02241993, -0.02280824, -0.02275554, 
    -0.02277918, -0.02306837, -0.02321557, -0.02352724, -0.02347033, 
    -0.02324159, -0.02273189, -0.02290358, -0.0224736, -0.02248321, 
    -0.02201443, -0.02222448, -0.02145225, -0.02166877, -0.02104945, 
    -0.02120339, -0.02105665, -0.02110103, -0.02105607, -0.02128232, 
    -0.02118507, -0.02138534, -0.02218497, -0.02194667, -0.02266562, 
    -0.02310999, -0.02341039, -0.02362607, -0.02359545, -0.02353719, 
    -0.02324026, -0.02296478, -0.02275719, -0.02261944, -0.02248459, 
    -0.02208156, -0.02187147, -0.02140873, -0.02149149, -0.02135152, 
    -0.02121877, -0.02099783, -0.02103403, -0.02093729, -0.02135523, 
    -0.02107647, -0.02153877, -0.02141125, -0.02244795, -0.02285714, 
    -0.02303335, -0.0231889, -0.02357193, -0.02330669, -0.02341086, 
    -0.02316387, -0.02300837, -0.02308514, -0.02261568, -0.02279696, 
    -0.02185908, -0.02225788, -0.0212342, -0.02147448, -0.02117705, 
    -0.02132827, -0.02106986, -0.02130227, -0.02090142, -0.0208152, 
    -0.02087408, -0.02064894, -0.02131524, -0.02105664, -0.02308729, 
    -0.02307475, -0.02301643, -0.02327398, -0.02328984, -0.02352879, 
    -0.02331606, -0.02322608, -0.0229994, -0.0228664, -0.02274075, 
    -0.02246708, -0.02216559, -0.0217513, -0.02145881, -0.02126512, 
    -0.02138367, -0.02127897, -0.02139605, -0.02145117, -0.02084746, 
    -0.02118416, -0.02068116, -0.02070866, -0.02093499, -0.02070555, 
    -0.02306595, -0.02313819, -0.02339086, -0.02319288, -0.02355497, 
    -0.02335153, -0.0232354, -0.02279313, -0.02269721, -0.02260861, 
    -0.02243474, -0.02221368, -0.02183151, -0.02150476, -0.02121108, 
    -0.02123245, -0.02122492, -0.02115985, -0.02132142, -0.02113345, 
    -0.02110207, -0.02118421, -0.02071234, -0.02084599, -0.02070924, 
    -0.02079614, -0.02311469, -0.0229934, -0.02305885, -0.02293593, 
    -0.02302245, -0.02264039, -0.02252717, -0.02200543, -0.022218, 
    -0.02188076, -0.0221835, -0.02212952, -0.0218698, -0.02216703, 
    -0.02152261, -0.02195723, -0.02115732, -0.02158336, -0.02113093, 
    -0.02121234, -0.02107774, -0.02095796, -0.02080833, -0.02053522, 
    -0.02059812, -0.02037196, -0.02281387, -0.02265887, -0.0226725, 
    -0.02251141, -0.02239306, -0.02213886, -0.02173758, -0.02188757, 
    -0.02161309, -0.02155843, -0.02197577, -0.02171849, -0.02255579, 
    -0.02241817, -0.02250002, -0.02280159, -0.02185287, -0.02233434, 
    -0.02145401, -0.02170836, -0.02097499, -0.02133629, -0.02063283, 
    -0.02033971, -0.02006803, -0.01975537, -0.02257478, -0.02267956, 
    -0.02249234, -0.02223601, -0.02200104, -0.02169275, -0.02166148, 
    -0.02160432, -0.02145705, -0.02133405, -0.02158626, -0.02130334, 
    -0.02238633, -0.02181162, -0.02271928, -0.02244174, -0.02225104, 
    -0.0223345, -0.02190478, -0.02180479, -0.02140347, -0.02160995, 
    -0.02041161, -0.02093272, -0.0195209, -0.01990479, -0.02271628, 
    -0.02257515, -0.02209123, -0.02232008, -0.02167234, -0.02151601, 
    -0.02138983, -0.02122966, -0.02121247, -0.02111826, -0.02127287, 
    -0.02112435, -0.02169209, -0.02143638, -0.02214601, -0.02197098, 
    -0.02205133, -0.0221398, -0.02186796, -0.02158226, -0.02157624, 
    -0.0214855, -0.02123193, -0.02166976, -0.02034531, -0.02115255, 
    -0.02242233, -0.02215504, -0.02211719, -0.02222013, -0.02153163, 
    -0.0217784, -0.02112056, -0.02129622, -0.02100922, -0.02115131, 
    -0.0211723, -0.02135652, -0.02147207, -0.02176702, -0.02201022, 
    -0.02220517, -0.02215968, -0.0219461, -0.02156492, -0.02121089, 
    -0.0212879, -0.02103089, -0.02171862, -0.02142732, -0.0215394, 
    -0.02124849, -0.02189156, -0.02134253, -0.0220343, -0.0219727, 
    -0.02178334, -0.02140769, -0.02132558, -0.02123822, -0.02129209, 
    -0.02155535, -0.02159883, -0.02178792, -0.02184043, -0.0219861, 
    -0.02210747, -0.02199654, -0.02188068, -0.02155525, -0.02126641, 
    -0.02095625, -0.02088111, -0.02052616, -0.02081455, -0.0203409, 
    -0.02074277, -0.02005246, -0.02131123, -0.02075479, -0.02177477, 
    -0.02166235, -0.02146055, -0.02100538, -0.02124984, -0.02096426, 
    -0.02160053, -0.02193875, -0.02202723, -0.02219326, -0.02202345, 
    -0.02203721, -0.02187592, -0.02192762, -0.02154453, -0.02174941, 
    -0.02117282, -0.02096651, -0.02039553, -0.02005377, -0.01971228, 
    -0.0195635, -0.01951846, -0.01949967,
  -0.02299437, -0.02262586, -0.02269703, -0.02240331, -0.02256576, 
    -0.02237413, -0.02291918, -0.02261135, -0.02280737, -0.02296097, 
    -0.02184449, -0.0223903, -0.02129234, -0.02162967, -0.0207927, 
    -0.02134445, -0.02068327, -0.02080845, -0.02043416, -0.02054066, 
    -0.02006951, -0.02038519, -0.01982979, -0.02014445, -0.02009487, 
    -0.02039569, -0.02227936, -0.02191167, -0.02230134, -0.02224846, 
    -0.02227218, -0.02256238, -0.02271008, -0.02302282, -0.02296572, 
    -0.0227362, -0.02222473, -0.02239702, -0.02196552, -0.02197517, 
    -0.02150472, -0.02171552, -0.02094049, -0.0211578, -0.0205362, 
    -0.02069071, -0.02054343, -0.02058798, -0.02054285, -0.02076994, 
    -0.02067232, -0.02087334, -0.02167587, -0.02143672, -0.02215823, 
    -0.02260414, -0.02290558, -0.02312198, -0.02309126, -0.0230328, 
    -0.02273486, -0.02245843, -0.02225011, -0.02211188, -0.02197656, 
    -0.02157209, -0.02136124, -0.02089682, -0.02097988, -0.02083939, 
    -0.02070615, -0.02048439, -0.02052072, -0.02042363, -0.02084311, 
    -0.02056332, -0.02102733, -0.02089934, -0.02193979, -0.02235041, 
    -0.02252724, -0.02268333, -0.02306767, -0.02280152, -0.02290605, 
    -0.02265821, -0.02250217, -0.02257921, -0.02210811, -0.02229003, 
    -0.02134881, -0.02174905, -0.02072164, -0.0209628, -0.02066428, 
    -0.02081606, -0.02055669, -0.02078996, -0.02038762, -0.02030108, 
    -0.02036018, -0.02013418, -0.02080297, -0.02054342, -0.02258137, 
    -0.02256878, -0.02251026, -0.0227687, -0.02278461, -0.02302438, 
    -0.02281092, -0.02272064, -0.02249317, -0.02235971, -0.02223362, 
    -0.02195899, -0.02165642, -0.02124063, -0.02094708, -0.02075267, 
    -0.02087167, -0.02076657, -0.02088409, -0.02093941, -0.02033345, 
    -0.02067141, -0.02016653, -0.02019413, -0.02042132, -0.02019102, 
    -0.02255995, -0.02263244, -0.02288598, -0.02268732, -0.02305065, 
    -0.02284652, -0.02272998, -0.02228618, -0.02218992, -0.02210101, 
    -0.02192652, -0.02170468, -0.02132114, -0.02099319, -0.02069843, 
    -0.02071988, -0.02071233, -0.02064701, -0.02080918, -0.02062051, 
    -0.02058901, -0.02067146, -0.02019783, -0.02033198, -0.02019471, 
    -0.02028194, -0.02260886, -0.02248715, -0.02255283, -0.02242948, 
    -0.0225163, -0.0221329, -0.02201929, -0.02149569, -0.02170902, 
    -0.02137056, -0.02167439, -0.02162023, -0.02135956, -0.02165787, 
    -0.02101111, -0.02144731, -0.02064447, -0.02107208, -0.02061798, 
    -0.02069969, -0.0205646, -0.02044437, -0.02029418, -0.02002004, 
    -0.02008318, -0.01985616, -0.022307, -0.02215145, -0.02216513, 
    -0.02200347, -0.0218847, -0.0216296, -0.02122687, -0.02137739, 
    -0.02110192, -0.02104706, -0.02146592, -0.02120771, -0.02204801, 
    -0.0219099, -0.02199204, -0.02229467, -0.02134258, -0.02182577, 
    -0.02094226, -0.02119754, -0.02046146, -0.02082411, -0.02011802, 
    -0.01982378, -0.01955106, -0.01923719, -0.02206707, -0.02217221, 
    -0.02198434, -0.02172709, -0.02149128, -0.02118187, -0.02115049, 
    -0.02109312, -0.02094531, -0.02082186, -0.02107499, -0.02079103, 
    -0.02187795, -0.02130117, -0.02221208, -0.02193356, -0.02174218, 
    -0.02182594, -0.02139468, -0.02129432, -0.02089154, -0.02109876, 
    -0.01989596, -0.02041904, -0.01900181, -0.01938719, -0.02220906, 
    -0.02206744, -0.0215818, -0.02181147, -0.02116139, -0.02100448, 
    -0.02087785, -0.02071709, -0.02069982, -0.02060527, -0.02076045, 
    -0.02061138, -0.02118121, -0.02092457, -0.02163677, -0.02146111, 
    -0.02154174, -0.02163053, -0.02135772, -0.02107098, -0.02106493, 
    -0.02097386, -0.02071936, -0.0211588, -0.01982941, -0.02063969, 
    -0.02191408, -0.02164583, -0.02160785, -0.02171115, -0.02102016, 
    -0.02126784, -0.02060757, -0.02078389, -0.02049582, -0.02063844, 
    -0.02065951, -0.02084441, -0.02096038, -0.02125641, -0.02150049, 
    -0.02169614, -0.02165049, -0.02143614, -0.02105358, -0.02069824, 
    -0.02077554, -0.02051757, -0.02120784, -0.02091547, -0.02102796, 
    -0.02073598, -0.0213814, -0.02083037, -0.02152466, -0.02146284, 
    -0.02127279, -0.02089577, -0.02081336, -0.02072567, -0.02077974, 
    -0.02104397, -0.02108761, -0.02127739, -0.02133009, -0.02147629, 
    -0.0215981, -0.02148676, -0.02137048, -0.02104387, -0.02075397, 
    -0.02044266, -0.02036723, -0.02001094, -0.02030043, -0.01982498, 
    -0.02022837, -0.01953544, -0.02079896, -0.02024044, -0.02126419, 
    -0.02115136, -0.02094882, -0.02049197, -0.02073734, -0.02045069, 
    -0.02108932, -0.02142877, -0.02151757, -0.02168419, -0.02151377, 
    -0.02152758, -0.02136571, -0.02141759, -0.02103312, -0.02123874, 
    -0.02066003, -0.02045295, -0.01987981, -0.01953675, -0.01919393, 
    -0.01904457, -0.01899936, -0.01898049,
  -0.02071496, -0.02036216, -0.02043028, -0.0201491, -0.02030462, 
    -0.02012118, -0.02064297, -0.02034826, -0.02053592, -0.02068298, 
    -0.01961423, -0.02013665, -0.01908586, -0.01940865, -0.01860785, 
    -0.01913572, -0.01850316, -0.01862291, -0.01826488, -0.01836675, 
    -0.01791614, -0.01821805, -0.01768691, -0.01798781, -0.01794039, 
    -0.01822809, -0.02003046, -0.01967853, -0.0200515, -0.02000089, 
    -0.02002359, -0.02030138, -0.02044279, -0.0207422, -0.02068753, 
    -0.02046779, -0.01997817, -0.02014309, -0.01973007, -0.01973931, 
    -0.01928908, -0.01949081, -0.01874923, -0.01895713, -0.01836249, 
    -0.01851028, -0.0183694, -0.01841201, -0.01836885, -0.01858607, 
    -0.01849269, -0.01868499, -0.01945287, -0.01922401, -0.01991451, 
    -0.02034136, -0.02062995, -0.02083715, -0.02080773, -0.02075176, 
    -0.02046651, -0.02020187, -0.02000246, -0.01987015, -0.01974063, 
    -0.01935355, -0.01915179, -0.01870745, -0.01878691, -0.01865251, 
    -0.01852505, -0.01831293, -0.01834768, -0.01825481, -0.01865607, 
    -0.01838842, -0.01883231, -0.01870986, -0.01970545, -0.02009847, 
    -0.02026775, -0.02041717, -0.02078514, -0.02053032, -0.0206304, 
    -0.02039313, -0.02024374, -0.02031749, -0.01986655, -0.02004067, 
    -0.01913989, -0.01952289, -0.01853987, -0.01877057, -0.01848499, 
    -0.01863019, -0.01838208, -0.01860523, -0.01822037, -0.0181376, 
    -0.01819412, -0.01797799, -0.01861767, -0.01836939, -0.02031956, 
    -0.02030751, -0.02025148, -0.0204989, -0.02051414, -0.02074369, 
    -0.02053932, -0.02045289, -0.02023512, -0.02010737, -0.01998668, 
    -0.01972382, -0.01943425, -0.01903639, -0.01875553, -0.01856955, 
    -0.01868339, -0.01858285, -0.01869527, -0.01874819, -0.01816856, 
    -0.01849182, -0.01800892, -0.01803531, -0.0182526, -0.01803234, 
    -0.02029905, -0.02036845, -0.02061119, -0.02042099, -0.02076885, 
    -0.0205734, -0.02046183, -0.02003699, -0.01994485, -0.01985975, 
    -0.01969275, -0.01948044, -0.01911342, -0.01879965, -0.01851766, 
    -0.01853818, -0.01853096, -0.01846848, -0.01862361, -0.01844313, 
    -0.018413, -0.01849187, -0.01803885, -0.01816715, -0.01803588, 
    -0.0181193, -0.02034587, -0.02022937, -0.02029224, -0.02017416, 
    -0.02025727, -0.01989028, -0.01978153, -0.01928044, -0.01948459, 
    -0.01916071, -0.01945145, -0.01939961, -0.01915019, -0.01943564, 
    -0.01881679, -0.01923415, -0.01846605, -0.01887512, -0.01844071, 
    -0.01851887, -0.01838965, -0.01827465, -0.018131, -0.01786883, 
    -0.01792921, -0.01771212, -0.02005691, -0.01990803, -0.01992112, 
    -0.01976639, -0.01965272, -0.01940858, -0.01902322, -0.01916725, 
    -0.01890367, -0.01885119, -0.01925196, -0.01900488, -0.01980902, 
    -0.01967684, -0.01975545, -0.02004511, -0.01913393, -0.01959632, 
    -0.01875092, -0.01899515, -0.018291, -0.01863789, -0.01796253, 
    -0.01768116, -0.01742041, -0.01712036, -0.01982726, -0.0199279, 
    -0.01974808, -0.01950188, -0.01927622, -0.01898016, -0.01895014, 
    -0.01889525, -0.01875384, -0.01863574, -0.01887791, -0.01860625, 
    -0.01964626, -0.01909432, -0.01996605, -0.01969948, -0.01951632, 
    -0.01959648, -0.01918378, -0.01908776, -0.0187024, -0.01890065, 
    -0.01775018, -0.01825042, -0.01689538, -0.01726375, -0.01996317, 
    -0.01982762, -0.01936284, -0.01958263, -0.01896057, -0.01881045, 
    -0.0186893, -0.01853551, -0.018519, -0.01842855, -0.01857699, -0.0184344, 
    -0.01897954, -0.018734, -0.01941544, -0.01924736, -0.01932451, 
    -0.01940948, -0.01914842, -0.01887407, -0.01886828, -0.01878115, 
    -0.01853769, -0.01895809, -0.01768654, -0.01846147, -0.01968083, 
    -0.01942412, -0.01938777, -0.01948663, -0.01882545, -0.01906242, 
    -0.01843075, -0.01859942, -0.01832386, -0.01846028, -0.01848044, 
    -0.01865731, -0.01876826, -0.01905148, -0.01928504, -0.01947226, 
    -0.01942857, -0.01922346, -0.01885742, -0.01851749, -0.01859143, 
    -0.01834466, -0.01900501, -0.01872529, -0.01883291, -0.01855358, 
    -0.01917108, -0.01864388, -0.01930816, -0.01924901, -0.01906715, 
    -0.01870644, -0.01862761, -0.01854373, -0.01859545, -0.01884822, 
    -0.01888997, -0.01907156, -0.01912198, -0.01926187, -0.01937844, 
    -0.0192719, -0.01916063, -0.01884813, -0.01857079, -0.01827301, 
    -0.01820087, -0.01786013, -0.01813698, -0.01768231, -0.01806807, 
    -0.01740547, -0.01861383, -0.01807961, -0.01905893, -0.01895097, 
    -0.0187572, -0.01832017, -0.01855489, -0.0182807, -0.01889161, 
    -0.0192164, -0.01930138, -0.01946082, -0.01929775, -0.01931096, 
    -0.01915606, -0.01920571, -0.01883784, -0.01903457, -0.01848093, 
    -0.01828286, -0.01773474, -0.01740673, -0.01707901, -0.01693625, 
    -0.01689303, -0.016875,
  -0.01736272, -0.01703657, -0.01709955, -0.01683965, -0.01698339, 
    -0.01681384, -0.01729616, -0.01702373, -0.0171972, -0.01733314, 
    -0.01634534, -0.01682814, -0.01585715, -0.01615538, -0.0154156, 
    -0.01590321, -0.01531892, -0.01542951, -0.01509887, -0.01519294, 
    -0.01477687, -0.01505562, -0.01456524, -0.01484303, -0.01479926, 
    -0.01506489, -0.01672999, -0.01640475, -0.01674944, -0.01670266, 
    -0.01672364, -0.0169804, -0.01711111, -0.01738789, -0.01733735, 
    -0.01713422, -0.01668166, -0.01683409, -0.01645238, -0.01646091, 
    -0.0160449, -0.01623129, -0.01554619, -0.01573823, -0.015189, 
    -0.01532549, -0.01519539, -0.01523474, -0.01519487, -0.01539549, 
    -0.01530925, -0.01548685, -0.01619623, -0.01598478, -0.01662283, 
    -0.01701736, -0.01728412, -0.01747568, -0.01744848, -0.01739673, 
    -0.01713303, -0.01688842, -0.01670411, -0.01658184, -0.01646214, 
    -0.01610447, -0.01591806, -0.01550759, -0.01558099, -0.01545686, 
    -0.01533913, -0.01514324, -0.01517533, -0.01508957, -0.01546014, 
    -0.01521295, -0.01562293, -0.01550983, -0.01642963, -0.01679285, 
    -0.01694931, -0.01708742, -0.01742759, -0.01719203, -0.01728454, 
    -0.0170652, -0.01692712, -0.01699529, -0.0165785, -0.01673943, 
    -0.01590707, -0.01626093, -0.01535282, -0.0155659, -0.01530214, 
    -0.01543623, -0.0152071, -0.01541318, -0.01505777, -0.01498134, 
    -0.01503353, -0.01483396, -0.01542467, -0.01519538, -0.0169972, 
    -0.01698606, -0.01693428, -0.01716298, -0.01717706, -0.01738928, 
    -0.01720034, -0.01712044, -0.01691915, -0.01680108, -0.01668953, 
    -0.0164466, -0.01617903, -0.01581145, -0.01555201, -0.01538023, 
    -0.01548537, -0.01539251, -0.01549634, -0.01554523, -0.01500993, 
    -0.01530844, -0.01486252, -0.0148869, -0.01508753, -0.01488415, 
    -0.01697825, -0.0170424, -0.01726678, -0.01709095, -0.01741253, 
    -0.01723185, -0.01712872, -0.01673603, -0.01665087, -0.01657222, 
    -0.01641789, -0.0162217, -0.01588261, -0.01559276, -0.01533231, 
    -0.01535126, -0.01534459, -0.01528689, -0.01543016, -0.01526348, 
    -0.01523565, -0.01530849, -0.01489016, -0.01500862, -0.01488741, 
    -0.01496444, -0.01702152, -0.01691383, -0.01697195, -0.01686281, 
    -0.01693962, -0.01660043, -0.01649993, -0.01603692, -0.01622554, 
    -0.0159263, -0.01619492, -0.01614702, -0.01591658, -0.01618031, 
    -0.0156086, -0.01599415, -0.01528465, -0.01566247, -0.01526124, 
    -0.01533343, -0.01521408, -0.01510789, -0.01497525, -0.01473319, 
    -0.01478893, -0.01458852, -0.01675444, -0.01661684, -0.01662893, 
    -0.01648595, -0.0163809, -0.01615531, -0.01579928, -0.01593234, 
    -0.01568885, -0.01564036, -0.0160106, -0.01578234, -0.01652534, 
    -0.01640319, -0.01647583, -0.01674354, -0.01590156, -0.01632879, 
    -0.01554775, -0.01577335, -0.01512299, -0.01544335, -0.01481969, 
    -0.01455994, -0.01431926, -0.01404235, -0.01654219, -0.0166352, 
    -0.01646902, -0.01624152, -0.01603302, -0.01575951, -0.01573177, 
    -0.01568107, -0.01555045, -0.01544136, -0.01566505, -0.01541413, 
    -0.01637493, -0.01586496, -0.01667047, -0.01642411, -0.01625486, 
    -0.01632893, -0.01594761, -0.0158589, -0.01550293, -0.01568606, 
    -0.01462365, -0.01508551, -0.01383476, -0.01417468, -0.0166678, 
    -0.01654252, -0.01611305, -0.01631613, -0.01574141, -0.01560274, 
    -0.01549083, -0.01534879, -0.01533354, -0.01525001, -0.0153871, 
    -0.01525541, -0.01575893, -0.01553212, -0.01616165, -0.01600635, 
    -0.01607764, -0.01615614, -0.01591495, -0.0156615, -0.01565616, 
    -0.01557568, -0.01535081, -0.01573912, -0.01456491, -0.01528042, 
    -0.01640688, -0.01616967, -0.01613608, -0.01622742, -0.01561659, 
    -0.01583549, -0.01525205, -0.01540782, -0.01515334, -0.01527932, 
    -0.01529793, -0.01546129, -0.01556377, -0.01582539, -0.01604116, 
    -0.01621415, -0.01617378, -0.01598427, -0.01564612, -0.01533215, 
    -0.01540044, -0.01517254, -0.01578246, -0.01552408, -0.01562348, 
    -0.01536548, -0.01593588, -0.01544889, -0.01606253, -0.01600787, 
    -0.01583987, -0.01550667, -0.01543385, -0.01535638, -0.01540415, 
    -0.01563763, -0.01567619, -0.01584394, -0.01589052, -0.01601976, 
    -0.01612746, -0.01602903, -0.01592623, -0.01563754, -0.01538138, 
    -0.01510638, -0.01503976, -0.01472516, -0.01498077, -0.014561, 
    -0.01491714, -0.01430547, -0.01542113, -0.01492779, -0.01583227, 
    -0.01573254, -0.01555355, -0.01514993, -0.01536669, -0.01511348, 
    -0.01567771, -0.01597775, -0.01605626, -0.01620358, -0.0160529, 
    -0.01606511, -0.01592201, -0.01596787, -0.01562804, -0.01580977, 
    -0.01529839, -0.01511547, -0.0146094, -0.01430663, -0.0140042, 
    -0.01387247, -0.0138326, -0.01381596,
  -0.01391834, -0.01359567, -0.01365795, -0.01340094, -0.01354307, 
    -0.01337543, -0.01385247, -0.01358296, -0.01375456, -0.01388907, 
    -0.01291255, -0.01338957, -0.01243078, -0.01272502, -0.01199555, 
    -0.01247621, -0.01190033, -0.01200926, -0.01168368, -0.01177628, 
    -0.01136692, -0.01164113, -0.01115891, -0.01143199, -0.01138894, 
    -0.01165025, -0.01329255, -0.01297122, -0.01331177, -0.01326554, 
    -0.01328627, -0.01354011, -0.01366939, -0.01394326, -0.01389324, 
    -0.01369225, -0.01324479, -0.01339545, -0.01301827, -0.01302669, 
    -0.01261599, -0.01279995, -0.01212422, -0.01231351, -0.01177241, 
    -0.0119068, -0.01177869, -0.01181743, -0.01177819, -0.01197574, 
    -0.0118908, -0.01206574, -0.01276534, -0.01255668, -0.01318666, 
    -0.01357666, -0.01384056, -0.01403015, -0.01400323, -0.01395201, 
    -0.01369108, -0.01344916, -0.01326698, -0.01314615, -0.01302791, 
    -0.01267477, -0.01249085, -0.01208619, -0.01215851, -0.0120362, 
    -0.01192023, -0.01172736, -0.01175895, -0.01167453, -0.01203943, 
    -0.01179599, -0.01219985, -0.01208839, -0.01299579, -0.01335468, 
    -0.01350937, -0.01364596, -0.01398255, -0.01374944, -0.01384098, 
    -0.01362398, -0.01348742, -0.01355484, -0.01314285, -0.01330188, 
    -0.01248001, -0.01282921, -0.01193372, -0.01214364, -0.0118838, 
    -0.01201588, -0.01179022, -0.01199317, -0.01164324, -0.01156803, 
    -0.01161938, -0.01142307, -0.01200449, -0.01177868, -0.01355672, 
    -0.01354571, -0.0134945, -0.0137207, -0.01373463, -0.01394463, 
    -0.01375767, -0.01367862, -0.01347955, -0.01336281, -0.01325256, 
    -0.01301255, -0.01274836, -0.01238571, -0.01212995, -0.01196072, 
    -0.01206429, -0.01197281, -0.0120751, -0.01212327, -0.01159616, 
    -0.01189001, -0.01145115, -0.01147513, -0.01167253, -0.01147242, 
    -0.01353798, -0.01360142, -0.0138234, -0.01364945, -0.01396764, 
    -0.01378884, -0.0136868, -0.01329852, -0.01321436, -0.01313665, 
    -0.0129842, -0.01279049, -0.01245589, -0.01217011, -0.01191352, 
    -0.01193218, -0.01192561, -0.01186878, -0.01200989, -0.01184573, 
    -0.01181833, -0.01189005, -0.01147834, -0.01159488, -0.01147564, 
    -0.01155141, -0.01358078, -0.01347429, -0.01353175, -0.01342384, 
    -0.01349979, -0.01316452, -0.01306523, -0.01260811, -0.01279427, 
    -0.01249898, -0.01276405, -0.01271677, -0.01248939, -0.01274963, 
    -0.01218572, -0.01256592, -0.01186658, -0.01223883, -0.01184353, 
    -0.01191462, -0.0117971, -0.01169256, -0.01156204, -0.01132398, 
    -0.01137879, -0.01118178, -0.01331672, -0.01318073, -0.01319268, 
    -0.01305142, -0.01294767, -0.01272495, -0.01237371, -0.01250494, 
    -0.01226483, -0.01221703, -0.01258215, -0.01235701, -0.01309033, 
    -0.01296968, -0.01304143, -0.01330594, -0.01247458, -0.01289621, 
    -0.01212576, -0.01234814, -0.01170742, -0.01202289, -0.01140904, 
    -0.0111537, -0.0109173, -0.01064556, -0.01310698, -0.01319888, 
    -0.0130347, -0.01281005, -0.01260427, -0.01233449, -0.01230714, 
    -0.01225716, -0.01212841, -0.01202093, -0.01224137, -0.0119941, 
    -0.01294178, -0.01243848, -0.01323372, -0.01299034, -0.01282322, 
    -0.01289635, -0.01252001, -0.01243251, -0.01208159, -0.01226208, 
    -0.01121631, -0.01167054, -0.01044201, -0.01077539, -0.01323109, 
    -0.01310731, -0.01268324, -0.01288371, -0.01231664, -0.01217995, 
    -0.01206967, -0.01192975, -0.01191473, -0.01183247, -0.01196748, 
    -0.01183779, -0.01233392, -0.01211035, -0.01273121, -0.01257795, 
    -0.01264829, -0.01272577, -0.01248778, -0.01223787, -0.0122326, 
    -0.01215328, -0.01193173, -0.01231439, -0.01115858, -0.01186241, 
    -0.01297333, -0.01273912, -0.01270597, -0.01279613, -0.0121936, 
    -0.01240942, -0.01183448, -0.01198789, -0.0117373, -0.01186133, 
    -0.01187966, -0.01204056, -0.01214154, -0.01239946, -0.0126123, 
    -0.01278303, -0.01274318, -0.01255617, -0.01222271, -0.01191336, 
    -0.01198062, -0.0117562, -0.01235712, -0.01210243, -0.01220039, 
    -0.01194619, -0.01250843, -0.01202834, -0.01263339, -0.01257946, 
    -0.01241373, -0.01208528, -0.01201354, -0.01193722, -0.01198428, 
    -0.01221434, -0.01225235, -0.01241775, -0.01246369, -0.01259119, 
    -0.01269746, -0.01260033, -0.01249891, -0.01221425, -0.01196185, 
    -0.01169107, -0.01162552, -0.01131608, -0.01156747, -0.01115474, 
    -0.01150487, -0.01090377, -0.012001, -0.01151535, -0.01240624, 
    -0.0123079, -0.01213147, -0.01173394, -0.01194737, -0.01169806, 
    -0.01225385, -0.01254974, -0.0126272, -0.0127726, -0.01262389, 
    -0.01263594, -0.01249475, -0.01253999, -0.01220489, -0.01238405, 
    -0.01188011, -0.01170002, -0.0112023, -0.0109049, -0.01060814, 
    -0.01047897, -0.01043989, -0.01042358,
  -0.008339484, -0.008031336, -0.008090762, -0.00784574, -0.007981176, 
    -0.007821442, -0.008276521, -0.008019218, -0.008182981, -0.008311507, 
    -0.007381527, -0.007834906, -0.006925563, -0.007203795, -0.006515509, 
    -0.006968473, -0.006426044, -0.006528391, -0.006222868, -0.006309649, 
    -0.005926748, -0.006183017, -0.005732945, -0.005987478, -0.005947292, 
    -0.006191558, -0.007742554, -0.007437192, -0.007760842, -0.00771685, 
    -0.00773658, -0.007978356, -0.008101672, -0.008363314, -0.008315488, 
    -0.008123491, -0.007697112, -0.007840505, -0.007481845, -0.007489848, 
    -0.007100612, -0.007274777, -0.006636536, -0.006814899, -0.006306015, 
    -0.006432121, -0.006311907, -0.006348243, -0.006311433, -0.00649689, 
    -0.006417101, -0.006581514, -0.007241987, -0.007044516, -0.007641828, 
    -0.008013207, -0.00826514, -0.00844643, -0.008420671, -0.008371679, 
    -0.008122374, -0.007891675, -0.00771822, -0.007603322, -0.007490999, 
    -0.007156228, -0.006982304, -0.006600746, -0.006668826, -0.006553721, 
    -0.006444736, -0.006263785, -0.006293395, -0.006214296, -0.006556764, 
    -0.006328126, -0.006707756, -0.006602814, -0.007460509, -0.007801688, 
    -0.007949048, -0.008079317, -0.008400894, -0.008178094, -0.008265537, 
    -0.008058345, -0.007928134, -0.007992398, -0.007600192, -0.00775143, 
    -0.006972064, -0.00730251, -0.006457401, -0.006654826, -0.006410528, 
    -0.006534618, -0.006322717, -0.006513269, -0.006184992, -0.006114619, 
    -0.006162664, -0.005979151, -0.006523912, -0.006311897, -0.007994197, 
    -0.007983696, -0.00793488, -0.008150652, -0.008163958, -0.008364622, 
    -0.008185953, -0.008110487, -0.007920629, -0.007809432, -0.007704504, 
    -0.007476423, -0.007225905, -0.006883011, -0.006641936, -0.006482768, 
    -0.006580144, -0.006494136, -0.006590317, -0.006635646, -0.006140934, 
    -0.006416353, -0.006005378, -0.00602777, -0.006212417, -0.006025245, 
    -0.007976328, -0.008036828, -0.008248742, -0.00808265, -0.008386634, 
    -0.008215723, -0.008118297, -0.00774823, -0.007668172, -0.007594293, 
    -0.007449508, -0.007265809, -0.006949276, -0.006679748, -0.006438428, 
    -0.00645596, -0.006449784, -0.006396427, -0.006528988, -0.006374795, 
    -0.006349089, -0.006416398, -0.006030771, -0.006139733, -0.006028247, 
    -0.006099071, -0.008017138, -0.007915615, -0.007970387, -0.007867551, 
    -0.007939918, -0.007620787, -0.007526447, -0.007093158, -0.007269396, 
    -0.006989988, -0.007240764, -0.007195991, -0.006980926, -0.007227103, 
    -0.006694449, -0.007053253, -0.006394357, -0.006744486, -0.006372727, 
    -0.006439462, -0.006329169, -0.006231185, -0.006109013, -0.005886693, 
    -0.005937818, -0.005754231, -0.007765549, -0.007636199, -0.007647561, 
    -0.007513325, -0.007414845, -0.007203737, -0.006871687, -0.006995615, 
    -0.00676899, -0.006723946, -0.0070686, -0.006855928, -0.007550283, 
    -0.007435729, -0.007503838, -0.007755292, -0.00696693, -0.007366024, 
    -0.006637985, -0.006847565, -0.006245106, -0.006541211, -0.00596605, 
    -0.005728099, -0.005508537, -0.005257096, -0.007566107, -0.007653448, 
    -0.00749745, -0.007284347, -0.007089522, -0.006834683, -0.006808889, 
    -0.006761762, -0.006640486, -0.006539368, -0.006746877, -0.006514144, 
    -0.007409253, -0.006932837, -0.007686588, -0.007455338, -0.007296829, 
    -0.007366164, -0.007009856, -0.006927195, -0.006596421, -0.006766397, 
    -0.005786372, -0.00621056, -0.005069459, -0.005377093, -0.007684084, 
    -0.007566417, -0.007164246, -0.007354178, -0.006817851, -0.006689011, 
    -0.006585207, -0.006453675, -0.006439568, -0.006362352, -0.006489127, 
    -0.006367343, -0.006834146, -0.006623484, -0.007209662, -0.007064636, 
    -0.007131171, -0.007204509, -0.006979407, -0.00674358, -0.006738617, 
    -0.006663894, -0.006455539, -0.006815721, -0.005732642, -0.00639045, 
    -0.007439188, -0.007217155, -0.007185764, -0.00727116, -0.00670187, 
    -0.006905397, -0.006364232, -0.006508301, -0.006273099, -0.006389431, 
    -0.006406635, -0.006557826, -0.006652844, -0.006895992, -0.007097123, 
    -0.007258746, -0.007220999, -0.007044042, -0.006729296, -0.006438278, 
    -0.006501468, -0.006290823, -0.006856038, -0.006616031, -0.006708271, 
    -0.006469117, -0.006998917, -0.006546337, -0.007117067, -0.007066059, 
    -0.006909469, -0.006599889, -0.006532413, -0.006460696, -0.006504909, 
    -0.006721407, -0.006757231, -0.006913261, -0.006956646, -0.007077151, 
    -0.007177707, -0.007085796, -0.006989922, -0.006721327, -0.00648383, 
    -0.006229791, -0.006168405, -0.005879332, -0.006114091, -0.00572907, 
    -0.006055566, -0.005495992, -0.006520626, -0.006065361, -0.006902397, 
    -0.006809607, -0.006643364, -0.006269956, -0.006470232, -0.006236337, 
    -0.006758639, -0.007037961, -0.007111212, -0.00724886, -0.007108082, 
    -0.00711948, -0.006985987, -0.007028745, -0.006712502, -0.006881452, 
    -0.00640706, -0.006238175, -0.005773329, -0.005497045, -0.005222552, 
    -0.005103488, -0.00506751, -0.005052503,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15 ;

 SOILWATER_10CM =
  439.2047, 440.8188, 440.505, 441.8078, 441.0847, 441.9382, 439.532, 
    440.8831, 440.0208, 439.3499, 444.3429, 441.8659, 446.9229, 445.337, 
    449.3265, 446.6761, 449.8619, 449.2495, 451.0932, 450.5646, 452.9283, 
    451.3373, 454.1558, 452.5479, 452.7993, 451.285, 442.3633, 444.0341, 
    442.2646, 442.5025, 442.3957, 441.0998, 440.4478, 439.0811, 439.3292, 
    440.3329, 442.6096, 441.8357, 443.7868, 443.7427, 445.921, 444.938, 
    448.6083, 447.5633, 450.5866, 449.8252, 450.5509, 450.3307, 450.5538, 
    449.4374, 449.9155, 448.9338, 445.1221, 446.2405, 442.91, 440.9151, 
    439.5913, 438.6521, 438.7848, 439.0379, 440.3387, 441.5616, 442.495, 
    443.12, 443.7364, 445.606, 446.5966, 448.82, 448.4179, 449.0989, 
    449.7495, 450.8435, 450.6633, 451.1458, 449.0807, 450.4526, 448.1891, 
    448.8076, 443.9053, 442.0443, 441.2559, 440.5654, 438.8869, 440.0464, 
    439.5893, 440.676, 441.3669, 441.0251, 443.1371, 442.3153, 446.6554, 
    444.7829, 449.6736, 448.5004, 449.955, 449.2123, 450.4854, 449.3396, 
    451.3253, 451.7585, 451.4624, 452.5998, 449.2761, 450.551, 441.0155, 
    441.0713, 441.331, 440.1903, 440.1205, 439.0744, 440.0052, 440.4012, 
    441.4069, 442.0027, 442.5693, 443.8168, 445.2126, 447.1684, 448.5764, 
    449.5217, 448.9418, 449.4538, 448.8816, 448.6135, 451.5962, 449.9201, 
    452.4361, 452.2966, 451.1573, 452.3123, 441.1104, 440.7897, 439.6768, 
    440.5477, 438.9605, 439.8495, 440.3602, 442.3328, 442.7666, 443.1694, 
    443.9654, 444.9883, 446.7862, 448.3538, 449.7873, 449.6822, 449.7192, 
    450.0399, 449.2459, 450.1703, 450.3257, 449.9197, 452.2779, 451.6035, 
    452.2936, 451.8544, 440.8939, 441.4337, 441.142, 441.6907, 441.3042, 
    443.0249, 443.5415, 445.9635, 444.9683, 446.5524, 445.1289, 445.381, 
    446.6047, 445.2057, 448.2675, 446.1908, 450.0524, 447.9744, 450.1828, 
    449.7811, 450.4462, 451.0424, 451.793, 453.1801, 452.8586, 454.0198, 
    442.2391, 442.9407, 442.8787, 443.6134, 444.1573, 445.3373, 447.2339, 
    446.52, 447.8307, 448.0942, 446.103, 447.3252, 443.4105, 444.0419, 
    443.6657, 442.2946, 446.6848, 444.4287, 448.5998, 447.3736, 450.9574, 
    449.1733, 452.6818, 454.187, 455.605, 457.2668, 443.3237, 442.8466, 
    443.7008, 444.8846, 445.984, 447.4484, 447.5982, 447.873, 448.5849, 
    449.1841, 447.9601, 449.3344, 444.1888, 446.8808, 442.6666, 443.9334, 
    444.8147, 444.4277, 446.4384, 446.9132, 448.8456, 447.8459, 453.8154, 
    451.1688, 458.5334, 456.4687, 442.6801, 443.3219, 445.5603, 444.4944, 
    447.5461, 448.2993, 448.9118, 449.696, 449.7805, 450.2455, 449.4837, 
    450.2153, 447.4515, 448.6853, 445.3039, 446.1256, 445.7474, 445.3329, 
    446.6129, 447.9795, 448.0083, 448.4471, 449.6855, 447.5585, 454.1584, 
    450.0766, 444.0225, 445.262, 445.4387, 444.9583, 448.2237, 447.039, 
    450.2341, 449.3692, 450.7867, 450.0821, 449.9785, 449.0743, 448.5121, 
    447.0933, 445.9408, 445.0279, 445.24, 446.2432, 448.063, 449.7883, 
    449.4101, 450.6789, 447.3244, 448.7295, 448.1862, 449.6034, 446.5012, 
    449.1433, 445.8274, 446.1175, 447.0155, 448.8251, 449.2255, 449.6539, 
    449.3894, 448.1092, 447.8995, 446.9935, 446.7438, 446.0543, 445.4841, 
    446.0051, 446.5528, 448.1096, 449.5155, 451.051, 451.4271, 453.2268, 
    451.762, 454.1813, 452.1248, 455.6876, 449.2961, 452.0636, 447.0562, 
    447.594, 448.5682, 450.8062, 449.5967, 451.0112, 447.8913, 446.278, 
    445.8607, 445.0834, 445.8784, 445.8137, 446.5752, 446.3304, 448.1613, 
    447.1773, 449.976, 450.9999, 453.8982, 455.6804, 457.4979, 458.3018, 
    458.5466, 458.649 ;

 SOMC_FIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOMHR =
  7.62417e-08, 7.645039e-08, 7.640983e-08, 7.657811e-08, 7.648478e-08, 
    7.659495e-08, 7.628402e-08, 7.645866e-08, 7.634719e-08, 7.626051e-08, 
    7.690453e-08, 7.658562e-08, 7.72358e-08, 7.70325e-08, 7.754317e-08, 
    7.720416e-08, 7.761152e-08, 7.753343e-08, 7.776852e-08, 7.770118e-08, 
    7.800173e-08, 7.77996e-08, 7.815754e-08, 7.795349e-08, 7.79854e-08, 
    7.779293e-08, 7.664984e-08, 7.686482e-08, 7.663709e-08, 7.666775e-08, 
    7.6654e-08, 7.648669e-08, 7.640234e-08, 7.622577e-08, 7.625783e-08, 
    7.638754e-08, 7.668154e-08, 7.658178e-08, 7.683326e-08, 7.682758e-08, 
    7.710744e-08, 7.698127e-08, 7.745152e-08, 7.731791e-08, 7.770399e-08, 
    7.760691e-08, 7.769943e-08, 7.767138e-08, 7.769979e-08, 7.755741e-08, 
    7.761841e-08, 7.749312e-08, 7.700489e-08, 7.71484e-08, 7.67203e-08, 
    7.646273e-08, 7.629168e-08, 7.617025e-08, 7.618742e-08, 7.622014e-08, 
    7.63883e-08, 7.654639e-08, 7.666684e-08, 7.674739e-08, 7.682677e-08, 
    7.706688e-08, 7.719401e-08, 7.747852e-08, 7.742722e-08, 7.751416e-08, 
    7.759725e-08, 7.773669e-08, 7.771375e-08, 7.777518e-08, 7.751189e-08, 
    7.768687e-08, 7.739798e-08, 7.7477e-08, 7.684823e-08, 7.66087e-08, 
    7.650677e-08, 7.641763e-08, 7.620062e-08, 7.635047e-08, 7.62914e-08, 
    7.643196e-08, 7.652125e-08, 7.647709e-08, 7.674959e-08, 7.664367e-08, 
    7.720153e-08, 7.696129e-08, 7.758756e-08, 7.743775e-08, 7.762347e-08, 
    7.752871e-08, 7.769106e-08, 7.754495e-08, 7.779804e-08, 7.785313e-08, 
    7.781549e-08, 7.796012e-08, 7.753685e-08, 7.769941e-08, 7.647585e-08, 
    7.648305e-08, 7.651661e-08, 7.636908e-08, 7.636006e-08, 7.622488e-08, 
    7.634518e-08, 7.639639e-08, 7.652643e-08, 7.660332e-08, 7.667641e-08, 
    7.683709e-08, 7.701648e-08, 7.726729e-08, 7.744746e-08, 7.75682e-08, 
    7.749417e-08, 7.755953e-08, 7.748646e-08, 7.745222e-08, 7.783248e-08, 
    7.761898e-08, 7.793933e-08, 7.792161e-08, 7.777663e-08, 7.79236e-08, 
    7.648811e-08, 7.644667e-08, 7.630274e-08, 7.641538e-08, 7.621016e-08, 
    7.632502e-08, 7.639106e-08, 7.664585e-08, 7.670185e-08, 7.675374e-08, 
    7.685622e-08, 7.698772e-08, 7.721835e-08, 7.741897e-08, 7.760209e-08, 
    7.758867e-08, 7.75934e-08, 7.763429e-08, 7.753298e-08, 7.765092e-08, 
    7.76707e-08, 7.761896e-08, 7.791923e-08, 7.783346e-08, 7.792123e-08, 
    7.786539e-08, 7.646015e-08, 7.652987e-08, 7.649219e-08, 7.656304e-08, 
    7.651312e-08, 7.673505e-08, 7.680158e-08, 7.711283e-08, 7.698513e-08, 
    7.718838e-08, 7.700579e-08, 7.703814e-08, 7.719496e-08, 7.701567e-08, 
    7.740789e-08, 7.714196e-08, 7.763587e-08, 7.737035e-08, 7.765251e-08, 
    7.76013e-08, 7.76861e-08, 7.776203e-08, 7.785756e-08, 7.803377e-08, 
    7.799298e-08, 7.814034e-08, 7.663383e-08, 7.672424e-08, 7.67163e-08, 
    7.681093e-08, 7.68809e-08, 7.703256e-08, 7.727571e-08, 7.718429e-08, 
    7.735214e-08, 7.738582e-08, 7.713083e-08, 7.728738e-08, 7.678477e-08, 
    7.686597e-08, 7.681763e-08, 7.664095e-08, 7.720533e-08, 7.691573e-08, 
    7.745043e-08, 7.729361e-08, 7.77512e-08, 7.752365e-08, 7.797052e-08, 
    7.816141e-08, 7.834114e-08, 7.8551e-08, 7.677361e-08, 7.671218e-08, 
    7.682219e-08, 7.697433e-08, 7.711554e-08, 7.730318e-08, 7.732238e-08, 
    7.735753e-08, 7.744857e-08, 7.75251e-08, 7.736862e-08, 7.754428e-08, 
    7.688477e-08, 7.723047e-08, 7.668893e-08, 7.685201e-08, 7.696537e-08, 
    7.691567e-08, 7.717384e-08, 7.723467e-08, 7.748181e-08, 7.735408e-08, 
    7.811428e-08, 7.777804e-08, 7.871082e-08, 7.845025e-08, 7.669071e-08, 
    7.677341e-08, 7.706114e-08, 7.692425e-08, 7.731571e-08, 7.741203e-08, 
    7.749034e-08, 7.759039e-08, 7.760121e-08, 7.766049e-08, 7.756335e-08, 
    7.765666e-08, 7.730358e-08, 7.746139e-08, 7.702828e-08, 7.713371e-08, 
    7.708522e-08, 7.703201e-08, 7.719621e-08, 7.737107e-08, 7.737484e-08, 
    7.74309e-08, 7.758878e-08, 7.73173e-08, 7.815761e-08, 7.763871e-08, 
    7.686358e-08, 7.702278e-08, 7.704556e-08, 7.698389e-08, 7.740237e-08, 
    7.725077e-08, 7.765905e-08, 7.754873e-08, 7.772948e-08, 7.763967e-08, 
    7.762645e-08, 7.751108e-08, 7.743924e-08, 7.725771e-08, 7.710998e-08, 
    7.699284e-08, 7.702008e-08, 7.714876e-08, 7.738178e-08, 7.760217e-08, 
    7.75539e-08, 7.771575e-08, 7.728734e-08, 7.746699e-08, 7.739755e-08, 
    7.75786e-08, 7.718186e-08, 7.751962e-08, 7.709549e-08, 7.713269e-08, 
    7.724775e-08, 7.747915e-08, 7.753039e-08, 7.758502e-08, 7.755131e-08, 
    7.73877e-08, 7.73609e-08, 7.724496e-08, 7.721293e-08, 7.712459e-08, 
    7.705142e-08, 7.711827e-08, 7.718845e-08, 7.738778e-08, 7.756736e-08, 
    7.77631e-08, 7.781102e-08, 7.803957e-08, 7.785348e-08, 7.81605e-08, 
    7.789941e-08, 7.835134e-08, 7.753925e-08, 7.789179e-08, 7.7253e-08, 
    7.732185e-08, 7.744634e-08, 7.773184e-08, 7.757776e-08, 7.775797e-08, 
    7.735986e-08, 7.715318e-08, 7.709974e-08, 7.699995e-08, 7.710202e-08, 
    7.709372e-08, 7.719137e-08, 7.716e-08, 7.73944e-08, 7.72685e-08, 
    7.762611e-08, 7.775656e-08, 7.812488e-08, 7.835057e-08, 7.858029e-08, 
    7.868167e-08, 7.871252e-08, 7.872543e-08 ;

 SOM_C_LEACHED =
  7.939695e-21, -2.654235e-20, -1.490632e-20, -5.089133e-20, -4.024473e-20, 
    1.172645e-19, 5.7726e-21, -5.84036e-21, 1.320764e-19, -4.989288e-20, 
    -1.387068e-20, -1.053238e-21, -5.226247e-20, 4.599828e-20, 4.729424e-20, 
    5.049176e-21, 1.950474e-21, 5.953245e-20, -2.228078e-20, -1.696911e-20, 
    -4.709543e-20, -1.951801e-20, -3.00313e-20, -1.74163e-20, -1.341106e-20, 
    -6.751767e-21, 6.294123e-21, -2.386452e-20, 4.134675e-20, 1.8652e-20, 
    1.974116e-20, -6.509668e-21, -1.205469e-20, -5.431513e-20, 3.109031e-20, 
    -3.929474e-20, -3.337577e-20, -1.062331e-19, -8.855361e-22, 
    -3.133699e-20, 2.023745e-20, 6.572702e-21, 1.956144e-21, -1.011344e-20, 
    4.968032e-20, -2.795793e-20, 4.939962e-20, -1.276805e-20, -4.078856e-20, 
    -5.142739e-21, -3.778742e-20, -8.048927e-20, -1.785106e-20, 1.50827e-20, 
    -1.831331e-20, -2.537412e-20, 1.119418e-21, -3.404177e-20, 4.146702e-22, 
    1.652078e-20, -1.165759e-20, 2.627175e-20, -6.167769e-22, -1.257942e-20, 
    1.998146e-20, 1.934019e-20, 1.002654e-19, -4.487015e-20, 4.450347e-20, 
    5.462449e-20, -2.8215e-20, -5.221893e-20, -3.950489e-20, -2.330974e-20, 
    -1.019402e-20, -2.003679e-20, 7.306861e-20, -1.755924e-20, -1.664644e-20, 
    -7.186419e-20, -1.126794e-20, -8.671549e-21, -2.584965e-20, 
    -1.513617e-21, 4.742063e-20, -2.113936e-20, -2.475167e-20, -3.12999e-20, 
    2.727747e-20, 2.158088e-20, -7.218732e-20, -1.553229e-21, 2.217378e-20, 
    3.470204e-21, 3.832439e-20, 5.977244e-20, -3.161453e-20, 7.535694e-20, 
    2.070424e-20, -9.568163e-21, 9.350686e-21, 8.320031e-20, 3.929183e-20, 
    8.537322e-23, 1.256103e-20, -5.447596e-20, -2.394943e-21, 6.973808e-20, 
    3.687124e-20, -5.113503e-20, -1.844153e-20, -3.433467e-22, 5.451583e-22, 
    3.274132e-20, 1.776737e-20, -3.349303e-20, -1.5243e-21, -2.701631e-20, 
    -2.027858e-20, -6.317533e-20, -2.727937e-20, 5.864468e-20, 1.334368e-20, 
    -1.367576e-20, -9.68362e-21, -1.134765e-20, 6.147209e-20, 3.724722e-20, 
    -2.979411e-20, -5.09447e-20, 1.623161e-20, 5.156021e-21, 5.672346e-20, 
    -3.140157e-20, 2.724152e-20, -3.57644e-20, 1.777411e-20, 2.94294e-20, 
    2.050826e-20, 1.27849e-20, -1.305542e-20, 7.336536e-20, -1.222341e-20, 
    4.453564e-20, 2.696583e-21, 2.363765e-20, -2.615166e-22, 5.554006e-20, 
    4.428068e-20, 5.088885e-21, -3.187777e-20, 3.011855e-20, -4.137695e-20, 
    -3.155841e-20, 4.030381e-21, -5.373741e-20, 3.491989e-20, 6.257735e-20, 
    -6.716697e-20, 1.052289e-20, -2.886607e-20, -1.311904e-20, 2.708065e-20, 
    -5.400357e-20, -3.671145e-20, -7.032332e-20, 5.09361e-20, 1.091246e-20, 
    -7.811077e-20, -1.938287e-20, 3.916781e-21, -4.999275e-20, -1.239309e-21, 
    2.102347e-20, 5.833533e-21, 2.274171e-20, 7.243316e-21, 3.193779e-21, 
    5.90839e-21, 1.991197e-20, -5.856275e-20, 2.727801e-22, -1.998648e-20, 
    -2.187989e-20, -3.443385e-20, 6.413966e-20, 1.446641e-20, 6.158044e-21, 
    1.344803e-20, 4.098172e-20, 9.055734e-21, -2.467451e-20, 6.849534e-21, 
    -2.052354e-20, -9.619456e-21, -4.962593e-20, 1.249975e-20, -9.069749e-21, 
    1.970008e-20, -4.259498e-20, 5.48214e-21, 9.257028e-21, -5.800523e-20, 
    -3.618251e-20, -1.60812e-21, -8.165273e-20, 5.190372e-20, -3.089055e-20, 
    -3.125651e-20, 1.328062e-20, 2.184683e-21, 2.832634e-20, -8.971611e-21, 
    -5.772057e-20, 4.674072e-21, -1.497352e-20, 9.792427e-21, -4.190195e-20, 
    4.620727e-20, -2.000292e-20, -8.648556e-21, 3.672302e-20, 7.441684e-20, 
    8.416885e-20, 2.813496e-20, 1.799908e-20, 3.918652e-20, 3.592479e-20, 
    -4.562384e-20, -1.472318e-20, -6.935011e-20, -6.901571e-21, 
    -2.763537e-20, -6.286242e-22, -3.471469e-20, 2.938166e-20, -2.252842e-20, 
    2.942307e-21, -3.784024e-20, 1.917576e-20, -2.181268e-21, -4.528149e-20, 
    -2.370833e-20, 2.883235e-21, -4.62452e-20, -2.263879e-20, -5.165297e-20, 
    -8.049011e-20, -6.695302e-22, -3.2065e-20, -3.836759e-20, -1.875059e-20, 
    4.101676e-20, 1.340455e-20, -1.360674e-20, -2.171467e-20, 9.404941e-20, 
    1.56226e-20, 2.430786e-20, 1.99281e-20, 2.818827e-20, -4.149741e-20, 
    5.00542e-20, 6.310025e-21, 2.939956e-21, -1.766585e-20, 5.41498e-20, 
    -3.892064e-20, -4.099066e-20, -4.085752e-21, -5.273604e-21, 4.421088e-20, 
    -2.060672e-20, 7.842344e-21, -2.015592e-20, 5.012503e-23, 3.590905e-20, 
    8.073685e-20, 1.417206e-20, 1.443865e-21, -7.414053e-20, 7.493831e-20, 
    -2.712259e-20, -1.35336e-20, 9.088423e-20, -2.727638e-20, 7.199219e-21, 
    6.77109e-20, -4.510791e-20, -6.539e-21, 1.306359e-20, -1.81773e-20, 
    2.60678e-20, 7.030175e-20, -9.495211e-21, 3.500623e-20, 5.00521e-20, 
    -6.904201e-20, -5.969431e-20, -2.412609e-20, 1.614833e-20, -5.997084e-21, 
    -9.28415e-22, 1.086351e-20, -9.526411e-21, 4.44363e-20, -4.277652e-20, 
    -1.026701e-20, 2.245122e-21, -1.058314e-21, -1.792009e-20, 3.949564e-20, 
    -4.510076e-20, -2.468206e-20, 2.977173e-20, 4.460849e-20, -8.889932e-20, 
    -1.978026e-20, 8.427996e-20, -4.84611e-20, -6.021599e-22, 1.353617e-20, 
    -1.948004e-20, 2.068666e-20, -1.142898e-20, -1.134058e-20, 5.050566e-20, 
    1.998355e-20, 3.113246e-20, -2.501845e-21, -9.570195e-21, -2.28972e-20, 
    3.098313e-20, 7.145115e-21, 7.341972e-21, 2.642847e-20, -3.088166e-20, 
    4.84502e-20 ;

 SR =
  7.624269e-08, 7.645139e-08, 7.641083e-08, 7.657911e-08, 7.648578e-08, 
    7.659595e-08, 7.628502e-08, 7.645966e-08, 7.634819e-08, 7.62615e-08, 
    7.690554e-08, 7.658662e-08, 7.723681e-08, 7.70335e-08, 7.754418e-08, 
    7.720516e-08, 7.761253e-08, 7.753444e-08, 7.776953e-08, 7.77022e-08, 
    7.800275e-08, 7.780061e-08, 7.815856e-08, 7.79545e-08, 7.798641e-08, 
    7.779394e-08, 7.665084e-08, 7.686582e-08, 7.663809e-08, 7.666875e-08, 
    7.6655e-08, 7.648769e-08, 7.640334e-08, 7.622676e-08, 7.625883e-08, 
    7.638853e-08, 7.668255e-08, 7.658277e-08, 7.683426e-08, 7.682858e-08, 
    7.710845e-08, 7.698227e-08, 7.745253e-08, 7.731892e-08, 7.7705e-08, 
    7.760792e-08, 7.770044e-08, 7.767239e-08, 7.77008e-08, 7.755842e-08, 
    7.761943e-08, 7.749413e-08, 7.700589e-08, 7.71494e-08, 7.67213e-08, 
    7.646373e-08, 7.629267e-08, 7.617125e-08, 7.618841e-08, 7.622113e-08, 
    7.638929e-08, 7.654739e-08, 7.666784e-08, 7.674839e-08, 7.682777e-08, 
    7.706788e-08, 7.719501e-08, 7.747953e-08, 7.742823e-08, 7.751517e-08, 
    7.759827e-08, 7.773771e-08, 7.771477e-08, 7.777619e-08, 7.75129e-08, 
    7.768788e-08, 7.739899e-08, 7.747801e-08, 7.684923e-08, 7.66097e-08, 
    7.650777e-08, 7.641862e-08, 7.620162e-08, 7.635147e-08, 7.629239e-08, 
    7.643295e-08, 7.652225e-08, 7.647809e-08, 7.67506e-08, 7.664466e-08, 
    7.720254e-08, 7.696229e-08, 7.758857e-08, 7.743876e-08, 7.762448e-08, 
    7.752973e-08, 7.769207e-08, 7.754596e-08, 7.779906e-08, 7.785415e-08, 
    7.78165e-08, 7.796114e-08, 7.753786e-08, 7.770043e-08, 7.647685e-08, 
    7.648405e-08, 7.651761e-08, 7.637008e-08, 7.636106e-08, 7.622587e-08, 
    7.634618e-08, 7.639739e-08, 7.652743e-08, 7.660432e-08, 7.667741e-08, 
    7.683809e-08, 7.701749e-08, 7.72683e-08, 7.744847e-08, 7.75692e-08, 
    7.749518e-08, 7.756054e-08, 7.748747e-08, 7.745323e-08, 7.78335e-08, 
    7.761999e-08, 7.794034e-08, 7.792262e-08, 7.777765e-08, 7.792462e-08, 
    7.648911e-08, 7.644767e-08, 7.630373e-08, 7.641638e-08, 7.621115e-08, 
    7.632602e-08, 7.639206e-08, 7.664685e-08, 7.670285e-08, 7.675474e-08, 
    7.685723e-08, 7.698873e-08, 7.721936e-08, 7.741998e-08, 7.76031e-08, 
    7.758969e-08, 7.759441e-08, 7.76353e-08, 7.7534e-08, 7.765193e-08, 
    7.767171e-08, 7.761997e-08, 7.792025e-08, 7.783448e-08, 7.792224e-08, 
    7.78664e-08, 7.646114e-08, 7.653087e-08, 7.649319e-08, 7.656404e-08, 
    7.651412e-08, 7.673605e-08, 7.680259e-08, 7.711383e-08, 7.698614e-08, 
    7.718939e-08, 7.70068e-08, 7.703915e-08, 7.719597e-08, 7.701667e-08, 
    7.74089e-08, 7.714296e-08, 7.763688e-08, 7.737135e-08, 7.765352e-08, 
    7.760231e-08, 7.768711e-08, 7.776304e-08, 7.785858e-08, 7.803479e-08, 
    7.7994e-08, 7.814135e-08, 7.663483e-08, 7.672524e-08, 7.671731e-08, 
    7.681193e-08, 7.68819e-08, 7.703356e-08, 7.727672e-08, 7.71853e-08, 
    7.735314e-08, 7.738683e-08, 7.713184e-08, 7.728839e-08, 7.678577e-08, 
    7.686698e-08, 7.681864e-08, 7.664195e-08, 7.720634e-08, 7.691673e-08, 
    7.745144e-08, 7.729462e-08, 7.775221e-08, 7.752466e-08, 7.797154e-08, 
    7.816244e-08, 7.834216e-08, 7.855203e-08, 7.677461e-08, 7.671318e-08, 
    7.682319e-08, 7.697533e-08, 7.711654e-08, 7.730418e-08, 7.732339e-08, 
    7.735854e-08, 7.744958e-08, 7.752611e-08, 7.736963e-08, 7.754529e-08, 
    7.688577e-08, 7.723148e-08, 7.668994e-08, 7.685301e-08, 7.696638e-08, 
    7.691667e-08, 7.717485e-08, 7.723568e-08, 7.748282e-08, 7.735509e-08, 
    7.811531e-08, 7.777906e-08, 7.871185e-08, 7.845127e-08, 7.669171e-08, 
    7.677441e-08, 7.706215e-08, 7.692525e-08, 7.731672e-08, 7.741303e-08, 
    7.749135e-08, 7.75914e-08, 7.760222e-08, 7.76615e-08, 7.756436e-08, 
    7.765767e-08, 7.730458e-08, 7.74624e-08, 7.702928e-08, 7.713471e-08, 
    7.708622e-08, 7.703301e-08, 7.719722e-08, 7.737208e-08, 7.737585e-08, 
    7.743191e-08, 7.758979e-08, 7.731831e-08, 7.815863e-08, 7.763973e-08, 
    7.686458e-08, 7.702379e-08, 7.704657e-08, 7.698489e-08, 7.740338e-08, 
    7.725177e-08, 7.766006e-08, 7.754974e-08, 7.77305e-08, 7.764068e-08, 
    7.762746e-08, 7.75121e-08, 7.744025e-08, 7.725872e-08, 7.711099e-08, 
    7.699384e-08, 7.702109e-08, 7.714976e-08, 7.738279e-08, 7.760318e-08, 
    7.755491e-08, 7.771676e-08, 7.728835e-08, 7.7468e-08, 7.739856e-08, 
    7.757962e-08, 7.718286e-08, 7.752063e-08, 7.709649e-08, 7.713369e-08, 
    7.724876e-08, 7.748016e-08, 7.75314e-08, 7.758604e-08, 7.755232e-08, 
    7.738871e-08, 7.736191e-08, 7.724597e-08, 7.721394e-08, 7.71256e-08, 
    7.705243e-08, 7.711927e-08, 7.718945e-08, 7.738879e-08, 7.756837e-08, 
    7.776411e-08, 7.781203e-08, 7.804059e-08, 7.785449e-08, 7.816151e-08, 
    7.790043e-08, 7.835236e-08, 7.754026e-08, 7.789281e-08, 7.725401e-08, 
    7.732286e-08, 7.744735e-08, 7.773286e-08, 7.757877e-08, 7.775899e-08, 
    7.736087e-08, 7.715419e-08, 7.710074e-08, 7.700096e-08, 7.710302e-08, 
    7.709473e-08, 7.719238e-08, 7.7161e-08, 7.739541e-08, 7.72695e-08, 
    7.762712e-08, 7.775758e-08, 7.812591e-08, 7.835159e-08, 7.858132e-08, 
    7.86827e-08, 7.871355e-08, 7.872645e-08 ;

 STORVEGC =
  0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545 ;

 STORVEGN =
  0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061 ;

 SUPPLEMENT_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SoilAlpha =
  0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 0.9999956, 
    0.9999956, 0.9999956 ;

 SoilAlpha_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TAUX =
  -0.3413633, -0.3413851, -0.3413841, -0.3413882, -0.341386, -0.3413886, 
    -0.341381, -0.3413852, -0.3413826, -0.3413639, -0.3413959, -0.3413884, 
    -0.34143, -0.341425, -0.3414377, -0.3414291, -0.3414395, -0.3414376, 
    -0.3414435, -0.3414418, -0.3414492, -0.3414443, -0.3414532, -0.3414481, 
    -0.3414488, -0.3414441, -0.34139, -0.341395, -0.3413897, -0.3413904, 
    -0.3413901, -0.341386, -0.3413838, -0.341363, -0.3413638, -0.3413835, 
    -0.3413907, -0.3413884, -0.3413945, -0.3413944, -0.3414269, -0.3413981, 
    -0.3414356, -0.3414322, -0.3414419, -0.3414395, -0.3414418, -0.3414411, 
    -0.3414418, -0.3414382, -0.3414397, -0.3414366, -0.3413987, -0.3414279, 
    -0.3413917, -0.3413852, -0.3413812, -0.3413617, -0.3413621, -0.3413629, 
    -0.3413835, -0.3413875, -0.3413905, -0.3413924, -0.3413944, -0.3414256, 
    -0.3414289, -0.3414361, -0.341435, -0.3414371, -0.3414392, -0.3414427, 
    -0.3414421, -0.3414437, -0.3414371, -0.3414414, -0.3414342, -0.3414362, 
    -0.3413945, -0.341389, -0.3413863, -0.3413843, -0.3413624, -0.3413826, 
    -0.3413812, -0.3413847, -0.3413869, -0.3413858, -0.3413925, -0.3413899, 
    -0.3414291, -0.3413976, -0.341439, -0.3414352, -0.3414399, -0.3414375, 
    -0.3414415, -0.3414379, -0.3414443, -0.3414456, -0.3414447, -0.3414483, 
    -0.3414377, -0.3414418, -0.3413858, -0.3413859, -0.3413868, -0.3413831, 
    -0.3413829, -0.341363, -0.3413825, -0.3413838, -0.341387, -0.3413889, 
    -0.3413907, -0.3413946, -0.3413989, -0.3414308, -0.3414355, -0.3414385, 
    -0.3414367, -0.3414383, -0.3414364, -0.3414356, -0.3414451, -0.3414397, 
    -0.3414478, -0.3414474, -0.3414437, -0.3414474, -0.3413861, -0.3413851, 
    -0.3413815, -0.3413843, -0.3413627, -0.341382, -0.3413836, -0.3413899, 
    -0.3413913, -0.3413926, -0.3413951, -0.3413983, -0.3414296, -0.3414347, 
    -0.3414394, -0.341439, -0.3414392, -0.3414401, -0.3414376, -0.3414406, 
    -0.341441, -0.3414398, -0.3414473, -0.3414452, -0.3414474, -0.341446, 
    -0.3413854, -0.3413871, -0.3413862, -0.3413879, -0.3413866, -0.341392, 
    -0.3413936, -0.3414269, -0.3413982, -0.3414288, -0.3413987, -0.3414251, 
    -0.3414288, -0.3414246, -0.3414343, -0.3414276, -0.3414402, -0.3414333, 
    -0.3414406, -0.3414393, -0.3414415, -0.3414433, -0.3414458, -0.3414501, 
    -0.3414491, -0.3414528, -0.3413897, -0.3413918, -0.3413917, -0.341394, 
    -0.3413957, -0.341425, -0.3414311, -0.3414288, -0.3414331, -0.3414339, 
    -0.3414275, -0.3414313, -0.3413933, -0.3413952, -0.3413941, -0.3413898, 
    -0.3414293, -0.3413965, -0.3414355, -0.3414316, -0.3414431, -0.3414373, 
    -0.3414485, -0.3414532, -0.3414579, -0.341463, -0.3413931, -0.3413916, 
    -0.3413943, -0.3413979, -0.3414271, -0.3414318, -0.3414323, -0.3414332, 
    -0.3414355, -0.3414374, -0.3414334, -0.3414379, -0.3413955, -0.3414299, 
    -0.341391, -0.3413949, -0.3413977, -0.3413965, -0.3414286, -0.3414301, 
    -0.3414363, -0.3414331, -0.341452, -0.3414436, -0.3414671, -0.3414605, 
    -0.3413911, -0.3413931, -0.3414257, -0.3413967, -0.3414322, -0.3414345, 
    -0.3414366, -0.341439, -0.3414393, -0.3414408, -0.3414384, -0.3414407, 
    -0.3414318, -0.3414358, -0.3414249, -0.3414275, -0.3414264, -0.341425, 
    -0.3414291, -0.3414334, -0.3414336, -0.341435, -0.3414386, -0.3414322, 
    -0.3414528, -0.3414399, -0.3413953, -0.3414246, -0.3414253, -0.3413982, 
    -0.3414343, -0.3414305, -0.3414408, -0.341438, -0.3414426, -0.3414403, 
    -0.34144, -0.3414371, -0.3414353, -0.3414306, -0.3414269, -0.3413985, 
    -0.3414247, -0.3414279, -0.3414337, -0.3414393, -0.3414381, -0.3414422, 
    -0.3414314, -0.3414359, -0.3414341, -0.3414387, -0.3414288, -0.3414369, 
    -0.3414266, -0.3414275, -0.3414304, -0.3414361, -0.3414375, -0.3414389, 
    -0.3414381, -0.3414339, -0.3414333, -0.3414304, -0.3414295, -0.3414274, 
    -0.3414255, -0.3414272, -0.3414289, -0.3414339, -0.3414384, -0.3414434, 
    -0.3414446, -0.3414501, -0.3414454, -0.3414529, -0.3414463, -0.3414578, 
    -0.3414375, -0.3414464, -0.3414306, -0.3414323, -0.3414353, -0.3414425, 
    -0.3414387, -0.3414432, -0.3414332, -0.341428, -0.3414267, -0.3413986, 
    -0.3414268, -0.3414266, -0.341429, -0.3414283, -0.3414341, -0.341431, 
    -0.3414399, -0.3414432, -0.3414524, -0.341458, -0.3414639, -0.3414665, 
    -0.3414673, -0.3414676 ;

 TAUY =
  -0.3413633, -0.3413851, -0.3413841, -0.3413882, -0.341386, -0.3413886, 
    -0.341381, -0.3413852, -0.3413826, -0.3413639, -0.3413959, -0.3413884, 
    -0.34143, -0.341425, -0.3414377, -0.3414291, -0.3414395, -0.3414376, 
    -0.3414435, -0.3414418, -0.3414492, -0.3414443, -0.3414532, -0.3414481, 
    -0.3414488, -0.3414441, -0.34139, -0.341395, -0.3413897, -0.3413904, 
    -0.3413901, -0.341386, -0.3413838, -0.341363, -0.3413638, -0.3413835, 
    -0.3413907, -0.3413884, -0.3413945, -0.3413944, -0.3414269, -0.3413981, 
    -0.3414356, -0.3414322, -0.3414419, -0.3414395, -0.3414418, -0.3414411, 
    -0.3414418, -0.3414382, -0.3414397, -0.3414366, -0.3413987, -0.3414279, 
    -0.3413917, -0.3413852, -0.3413812, -0.3413617, -0.3413621, -0.3413629, 
    -0.3413835, -0.3413875, -0.3413905, -0.3413924, -0.3413944, -0.3414256, 
    -0.3414289, -0.3414361, -0.341435, -0.3414371, -0.3414392, -0.3414427, 
    -0.3414421, -0.3414437, -0.3414371, -0.3414414, -0.3414342, -0.3414362, 
    -0.3413945, -0.341389, -0.3413863, -0.3413843, -0.3413624, -0.3413826, 
    -0.3413812, -0.3413847, -0.3413869, -0.3413858, -0.3413925, -0.3413899, 
    -0.3414291, -0.3413976, -0.341439, -0.3414352, -0.3414399, -0.3414375, 
    -0.3414415, -0.3414379, -0.3414443, -0.3414456, -0.3414447, -0.3414483, 
    -0.3414377, -0.3414418, -0.3413858, -0.3413859, -0.3413868, -0.3413831, 
    -0.3413829, -0.341363, -0.3413825, -0.3413838, -0.341387, -0.3413889, 
    -0.3413907, -0.3413946, -0.3413989, -0.3414308, -0.3414355, -0.3414385, 
    -0.3414367, -0.3414383, -0.3414364, -0.3414356, -0.3414451, -0.3414397, 
    -0.3414478, -0.3414474, -0.3414437, -0.3414474, -0.3413861, -0.3413851, 
    -0.3413815, -0.3413843, -0.3413627, -0.341382, -0.3413836, -0.3413899, 
    -0.3413913, -0.3413926, -0.3413951, -0.3413983, -0.3414296, -0.3414347, 
    -0.3414394, -0.341439, -0.3414392, -0.3414401, -0.3414376, -0.3414406, 
    -0.341441, -0.3414398, -0.3414473, -0.3414452, -0.3414474, -0.341446, 
    -0.3413854, -0.3413871, -0.3413862, -0.3413879, -0.3413866, -0.341392, 
    -0.3413936, -0.3414269, -0.3413982, -0.3414288, -0.3413987, -0.3414251, 
    -0.3414288, -0.3414246, -0.3414343, -0.3414276, -0.3414402, -0.3414333, 
    -0.3414406, -0.3414393, -0.3414415, -0.3414433, -0.3414458, -0.3414501, 
    -0.3414491, -0.3414528, -0.3413897, -0.3413918, -0.3413917, -0.341394, 
    -0.3413957, -0.341425, -0.3414311, -0.3414288, -0.3414331, -0.3414339, 
    -0.3414275, -0.3414313, -0.3413933, -0.3413952, -0.3413941, -0.3413898, 
    -0.3414293, -0.3413965, -0.3414355, -0.3414316, -0.3414431, -0.3414373, 
    -0.3414485, -0.3414532, -0.3414579, -0.341463, -0.3413931, -0.3413916, 
    -0.3413943, -0.3413979, -0.3414271, -0.3414318, -0.3414323, -0.3414332, 
    -0.3414355, -0.3414374, -0.3414334, -0.3414379, -0.3413955, -0.3414299, 
    -0.341391, -0.3413949, -0.3413977, -0.3413965, -0.3414286, -0.3414301, 
    -0.3414363, -0.3414331, -0.341452, -0.3414436, -0.3414671, -0.3414605, 
    -0.3413911, -0.3413931, -0.3414257, -0.3413967, -0.3414322, -0.3414345, 
    -0.3414366, -0.341439, -0.3414393, -0.3414408, -0.3414384, -0.3414407, 
    -0.3414318, -0.3414358, -0.3414249, -0.3414275, -0.3414264, -0.341425, 
    -0.3414291, -0.3414334, -0.3414336, -0.341435, -0.3414386, -0.3414322, 
    -0.3414528, -0.3414399, -0.3413953, -0.3414246, -0.3414253, -0.3413982, 
    -0.3414343, -0.3414305, -0.3414408, -0.341438, -0.3414426, -0.3414403, 
    -0.34144, -0.3414371, -0.3414353, -0.3414306, -0.3414269, -0.3413985, 
    -0.3414247, -0.3414279, -0.3414337, -0.3414393, -0.3414381, -0.3414422, 
    -0.3414314, -0.3414359, -0.3414341, -0.3414387, -0.3414288, -0.3414369, 
    -0.3414266, -0.3414275, -0.3414304, -0.3414361, -0.3414375, -0.3414389, 
    -0.3414381, -0.3414339, -0.3414333, -0.3414304, -0.3414295, -0.3414274, 
    -0.3414255, -0.3414272, -0.3414289, -0.3414339, -0.3414384, -0.3414434, 
    -0.3414446, -0.3414501, -0.3414454, -0.3414529, -0.3414463, -0.3414578, 
    -0.3414375, -0.3414464, -0.3414306, -0.3414323, -0.3414353, -0.3414425, 
    -0.3414387, -0.3414432, -0.3414332, -0.341428, -0.3414267, -0.3413986, 
    -0.3414268, -0.3414266, -0.341429, -0.3414283, -0.3414341, -0.341431, 
    -0.3414399, -0.3414432, -0.3414524, -0.341458, -0.3414639, -0.3414665, 
    -0.3414673, -0.3414676 ;

 TBOT =
  253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605 ;

 TBUILD =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TG =
  261.7208, 261.7411, 261.7372, 261.7536, 261.7445, 261.7553, 261.7249, 
    261.7419, 261.731, 261.7226, 261.7856, 261.7544, 261.8176, 261.7977, 
    261.8476, 261.8145, 261.8543, 261.8467, 261.8697, 261.8631, 261.8924, 
    261.8727, 261.9076, 261.8877, 261.8908, 261.872, 261.7607, 261.7817, 
    261.7594, 261.7624, 261.7611, 261.7447, 261.7364, 261.7192, 261.7224, 
    261.735, 261.7638, 261.754, 261.7786, 261.7781, 261.805, 261.7931, 
    261.8387, 261.8256, 261.8633, 261.8539, 261.8629, 261.8602, 261.8629, 
    261.849, 261.855, 261.8427, 261.7954, 261.809, 261.7676, 261.7423, 
    261.7256, 261.7138, 261.7155, 261.7187, 261.7351, 261.7505, 261.7623, 
    261.7702, 261.778, 261.801, 261.8135, 261.8413, 261.8363, 261.8448, 
    261.8529, 261.8665, 261.8643, 261.8703, 261.8446, 261.8617, 261.8334, 
    261.8412, 261.7801, 261.7567, 261.7466, 261.7379, 261.7168, 261.7314, 
    261.7256, 261.7393, 261.7481, 261.7438, 261.7704, 261.7601, 261.8142, 
    261.7911, 261.852, 261.8373, 261.8555, 261.8462, 261.8621, 261.8478, 
    261.8725, 261.8779, 261.8742, 261.8884, 261.847, 261.8629, 261.7437, 
    261.7444, 261.7477, 261.7332, 261.7323, 261.7191, 261.7308, 261.7359, 
    261.7486, 261.7561, 261.7633, 261.779, 261.7965, 261.8206, 261.8383, 
    261.8501, 261.8428, 261.8492, 261.8421, 261.8387, 261.8759, 261.855, 
    261.8863, 261.8846, 261.8704, 261.8848, 261.7448, 261.7408, 261.7267, 
    261.7377, 261.7177, 261.7289, 261.7353, 261.7603, 261.7658, 261.7708, 
    261.7809, 261.7937, 261.8159, 261.8355, 261.8534, 261.8521, 261.8525, 
    261.8565, 261.8466, 261.8582, 261.8601, 261.855, 261.8844, 261.876, 
    261.8846, 261.8791, 261.7421, 261.7489, 261.7452, 261.7522, 261.7473, 
    261.769, 261.7755, 261.8055, 261.7935, 261.8129, 261.7955, 261.7982, 
    261.8136, 261.7961, 261.8344, 261.8084, 261.8567, 261.8307, 261.8583, 
    261.8533, 261.8616, 261.869, 261.8784, 261.8955, 261.8916, 261.9059, 
    261.7591, 261.7679, 261.7672, 261.7764, 261.7833, 261.7977, 261.8215, 
    261.8125, 261.8289, 261.8322, 261.8073, 261.8226, 261.7739, 261.7818, 
    261.7771, 261.7598, 261.8146, 261.7867, 261.8386, 261.8232, 261.868, 
    261.8457, 261.8894, 261.908, 261.9256, 261.946, 261.7728, 261.7668, 
    261.7776, 261.7924, 261.8058, 261.8242, 261.826, 261.8295, 261.8384, 
    261.8459, 261.8306, 261.8477, 261.7836, 261.817, 261.7645, 261.7805, 
    261.7915, 261.7867, 261.8115, 261.8175, 261.8416, 261.8291, 261.9034, 
    261.8706, 261.9616, 261.9362, 261.7647, 261.7728, 261.8005, 261.7875, 
    261.8254, 261.8348, 261.8425, 261.8522, 261.8533, 261.8591, 261.8496, 
    261.8587, 261.8242, 261.8396, 261.7973, 261.8076, 261.8029, 261.7976, 
    261.8137, 261.8308, 261.8312, 261.8366, 261.852, 261.8256, 261.9076, 
    261.8569, 261.7816, 261.7967, 261.799, 261.7934, 261.8339, 261.819, 
    261.8589, 261.8482, 261.8658, 261.8571, 261.8558, 261.8445, 261.8375, 
    261.8197, 261.8053, 261.7943, 261.7965, 261.8091, 261.8318, 261.8534, 
    261.8487, 261.8645, 261.8226, 261.8402, 261.8334, 261.8511, 261.8123, 
    261.8453, 261.8039, 261.8075, 261.8188, 261.8413, 261.8464, 261.8517, 
    261.8484, 261.8324, 261.8298, 261.8185, 261.8153, 261.8067, 261.7996, 
    261.8061, 261.8129, 261.8324, 261.85, 261.8691, 261.8738, 261.8961, 
    261.8779, 261.9079, 261.8824, 261.9265, 261.8472, 261.8817, 261.8193, 
    261.826, 261.8381, 261.8661, 261.851, 261.8686, 261.8297, 261.8095, 
    261.8043, 261.7949, 261.8045, 261.8037, 261.8132, 261.8102, 261.8331, 
    261.8208, 261.8557, 261.8685, 261.9044, 261.9265, 261.9489, 261.9588, 
    261.9618, 261.963 ;

 TG_R =
  261.7208, 261.7411, 261.7372, 261.7536, 261.7445, 261.7553, 261.7249, 
    261.7419, 261.731, 261.7226, 261.7856, 261.7544, 261.8176, 261.7977, 
    261.8476, 261.8145, 261.8543, 261.8467, 261.8697, 261.8631, 261.8924, 
    261.8727, 261.9076, 261.8877, 261.8908, 261.872, 261.7607, 261.7817, 
    261.7594, 261.7624, 261.7611, 261.7447, 261.7364, 261.7192, 261.7224, 
    261.735, 261.7638, 261.754, 261.7786, 261.7781, 261.805, 261.7931, 
    261.8387, 261.8256, 261.8633, 261.8539, 261.8629, 261.8602, 261.8629, 
    261.849, 261.855, 261.8427, 261.7954, 261.809, 261.7676, 261.7423, 
    261.7256, 261.7138, 261.7155, 261.7187, 261.7351, 261.7505, 261.7623, 
    261.7702, 261.778, 261.801, 261.8135, 261.8413, 261.8363, 261.8448, 
    261.8529, 261.8665, 261.8643, 261.8703, 261.8446, 261.8617, 261.8334, 
    261.8412, 261.7801, 261.7567, 261.7466, 261.7379, 261.7168, 261.7314, 
    261.7256, 261.7393, 261.7481, 261.7438, 261.7704, 261.7601, 261.8142, 
    261.7911, 261.852, 261.8373, 261.8555, 261.8462, 261.8621, 261.8478, 
    261.8725, 261.8779, 261.8742, 261.8884, 261.847, 261.8629, 261.7437, 
    261.7444, 261.7477, 261.7332, 261.7323, 261.7191, 261.7308, 261.7359, 
    261.7486, 261.7561, 261.7633, 261.779, 261.7965, 261.8206, 261.8383, 
    261.8501, 261.8428, 261.8492, 261.8421, 261.8387, 261.8759, 261.855, 
    261.8863, 261.8846, 261.8704, 261.8848, 261.7448, 261.7408, 261.7267, 
    261.7377, 261.7177, 261.7289, 261.7353, 261.7603, 261.7658, 261.7708, 
    261.7809, 261.7937, 261.8159, 261.8355, 261.8534, 261.8521, 261.8525, 
    261.8565, 261.8466, 261.8582, 261.8601, 261.855, 261.8844, 261.876, 
    261.8846, 261.8791, 261.7421, 261.7489, 261.7452, 261.7522, 261.7473, 
    261.769, 261.7755, 261.8055, 261.7935, 261.8129, 261.7955, 261.7982, 
    261.8136, 261.7961, 261.8344, 261.8084, 261.8567, 261.8307, 261.8583, 
    261.8533, 261.8616, 261.869, 261.8784, 261.8955, 261.8916, 261.9059, 
    261.7591, 261.7679, 261.7672, 261.7764, 261.7833, 261.7977, 261.8215, 
    261.8125, 261.8289, 261.8322, 261.8073, 261.8226, 261.7739, 261.7818, 
    261.7771, 261.7598, 261.8146, 261.7867, 261.8386, 261.8232, 261.868, 
    261.8457, 261.8894, 261.908, 261.9256, 261.946, 261.7728, 261.7668, 
    261.7776, 261.7924, 261.8058, 261.8242, 261.826, 261.8295, 261.8384, 
    261.8459, 261.8306, 261.8477, 261.7836, 261.817, 261.7645, 261.7805, 
    261.7915, 261.7867, 261.8115, 261.8175, 261.8416, 261.8291, 261.9034, 
    261.8706, 261.9616, 261.9362, 261.7647, 261.7728, 261.8005, 261.7875, 
    261.8254, 261.8348, 261.8425, 261.8522, 261.8533, 261.8591, 261.8496, 
    261.8587, 261.8242, 261.8396, 261.7973, 261.8076, 261.8029, 261.7976, 
    261.8137, 261.8308, 261.8312, 261.8366, 261.852, 261.8256, 261.9076, 
    261.8569, 261.7816, 261.7967, 261.799, 261.7934, 261.8339, 261.819, 
    261.8589, 261.8482, 261.8658, 261.8571, 261.8558, 261.8445, 261.8375, 
    261.8197, 261.8053, 261.7943, 261.7965, 261.8091, 261.8318, 261.8534, 
    261.8487, 261.8645, 261.8226, 261.8402, 261.8334, 261.8511, 261.8123, 
    261.8453, 261.8039, 261.8075, 261.8188, 261.8413, 261.8464, 261.8517, 
    261.8484, 261.8324, 261.8298, 261.8185, 261.8153, 261.8067, 261.7996, 
    261.8061, 261.8129, 261.8324, 261.85, 261.8691, 261.8738, 261.8961, 
    261.8779, 261.9079, 261.8824, 261.9265, 261.8472, 261.8817, 261.8193, 
    261.826, 261.8381, 261.8661, 261.851, 261.8686, 261.8297, 261.8095, 
    261.8043, 261.7949, 261.8045, 261.8037, 261.8132, 261.8102, 261.8331, 
    261.8208, 261.8557, 261.8685, 261.9044, 261.9265, 261.9489, 261.9588, 
    261.9618, 261.963 ;

 TG_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TH2OSFC =
  254.6773, 254.6788, 254.6785, 254.6797, 254.6791, 254.6799, 254.6776, 
    254.6788, 254.6781, 254.6774, 254.6821, 254.6798, 254.6846, 254.6831, 
    254.6869, 254.6843, 254.6874, 254.6868, 254.6886, 254.6881, 254.6903, 
    254.6888, 254.6915, 254.6899, 254.6902, 254.6888, 254.6803, 254.6818, 
    254.6802, 254.6804, 254.6803, 254.6791, 254.6784, 254.6772, 254.6774, 
    254.6783, 254.6805, 254.6798, 254.6816, 254.6816, 254.6837, 254.6827, 
    254.6862, 254.6852, 254.6881, 254.6874, 254.688, 254.6879, 254.688, 
    254.687, 254.6875, 254.6865, 254.6829, 254.684, 254.6808, 254.6789, 
    254.6776, 254.6768, 254.6769, 254.6771, 254.6783, 254.6795, 254.6804, 
    254.681, 254.6816, 254.6833, 254.6843, 254.6864, 254.686, 254.6867, 
    254.6873, 254.6883, 254.6882, 254.6886, 254.6867, 254.688, 254.6858, 
    254.6864, 254.6817, 254.68, 254.6792, 254.6786, 254.677, 254.6781, 
    254.6776, 254.6787, 254.6793, 254.679, 254.681, 254.6802, 254.6843, 
    254.6826, 254.6872, 254.6861, 254.6875, 254.6868, 254.688, 254.6869, 
    254.6888, 254.6892, 254.6889, 254.69, 254.6868, 254.688, 254.679, 
    254.679, 254.6793, 254.6782, 254.6781, 254.6772, 254.678, 254.6784, 
    254.6794, 254.6799, 254.6805, 254.6817, 254.683, 254.6848, 254.6862, 
    254.6871, 254.6865, 254.687, 254.6865, 254.6862, 254.689, 254.6875, 
    254.6898, 254.6897, 254.6886, 254.6897, 254.6791, 254.6788, 254.6777, 
    254.6786, 254.677, 254.6779, 254.6784, 254.6802, 254.6807, 254.681, 
    254.6818, 254.6828, 254.6845, 254.686, 254.6873, 254.6872, 254.6873, 
    254.6876, 254.6868, 254.6877, 254.6878, 254.6875, 254.6897, 254.6891, 
    254.6897, 254.6893, 254.6789, 254.6794, 254.6791, 254.6796, 254.6793, 
    254.6809, 254.6814, 254.6837, 254.6828, 254.6842, 254.6829, 254.6831, 
    254.6843, 254.683, 254.6859, 254.6839, 254.6876, 254.6856, 254.6877, 
    254.6873, 254.688, 254.6885, 254.6892, 254.6905, 254.6902, 254.6913, 
    254.6802, 254.6808, 254.6808, 254.6815, 254.682, 254.6831, 254.6849, 
    254.6842, 254.6855, 254.6857, 254.6838, 254.685, 254.6813, 254.6819, 
    254.6815, 254.6802, 254.6844, 254.6822, 254.6862, 254.685, 254.6884, 
    254.6867, 254.6901, 254.6915, 254.6928, 254.6944, 254.6812, 254.6807, 
    254.6816, 254.6827, 254.6837, 254.6851, 254.6853, 254.6855, 254.6862, 
    254.6868, 254.6856, 254.6869, 254.682, 254.6846, 254.6806, 254.6817, 
    254.6826, 254.6822, 254.6842, 254.6846, 254.6864, 254.6855, 254.6911, 
    254.6886, 254.6956, 254.6936, 254.6806, 254.6812, 254.6833, 254.6823, 
    254.6852, 254.6859, 254.6865, 254.6872, 254.6873, 254.6878, 254.687, 
    254.6877, 254.6851, 254.6863, 254.6831, 254.6839, 254.6835, 254.6831, 
    254.6843, 254.6856, 254.6856, 254.6861, 254.6871, 254.6852, 254.6914, 
    254.6875, 254.6819, 254.683, 254.6832, 254.6828, 254.6858, 254.6847, 
    254.6878, 254.6869, 254.6883, 254.6876, 254.6875, 254.6867, 254.6861, 
    254.6848, 254.6837, 254.6828, 254.683, 254.684, 254.6857, 254.6873, 
    254.687, 254.6882, 254.685, 254.6863, 254.6858, 254.6871, 254.6842, 
    254.6866, 254.6836, 254.6839, 254.6847, 254.6864, 254.6868, 254.6872, 
    254.687, 254.6857, 254.6855, 254.6847, 254.6844, 254.6838, 254.6833, 
    254.6837, 254.6842, 254.6857, 254.6871, 254.6885, 254.6889, 254.6905, 
    254.6892, 254.6914, 254.6895, 254.6929, 254.6868, 254.6894, 254.6847, 
    254.6853, 254.6862, 254.6883, 254.6871, 254.6885, 254.6855, 254.684, 
    254.6836, 254.6829, 254.6836, 254.6836, 254.6843, 254.6841, 254.6858, 
    254.6849, 254.6875, 254.6885, 254.6912, 254.6929, 254.6946, 254.6954, 
    254.6956, 254.6957 ;

 THBOT =
  253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605 ;

 TKE1 =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TLAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 TLAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TOTCOLC =
  18.2395, 18.23949, 18.23949, 18.23948, 18.23949, 18.23948, 18.2395, 
    18.23949, 18.2395, 18.2395, 18.23947, 18.23948, 18.23945, 18.23946, 
    18.23944, 18.23945, 18.23944, 18.23944, 18.23943, 18.23943, 18.23942, 
    18.23943, 18.23941, 18.23942, 18.23942, 18.23943, 18.23948, 18.23947, 
    18.23948, 18.23948, 18.23948, 18.23949, 18.23949, 18.2395, 18.2395, 
    18.23949, 18.23948, 18.23948, 18.23947, 18.23947, 18.23946, 18.23947, 
    18.23944, 18.23945, 18.23943, 18.23944, 18.23943, 18.23943, 18.23943, 
    18.23944, 18.23944, 18.23944, 18.23946, 18.23946, 18.23948, 18.23949, 
    18.2395, 18.2395, 18.2395, 18.2395, 18.23949, 18.23949, 18.23948, 
    18.23948, 18.23947, 18.23946, 18.23945, 18.23944, 18.23944, 18.23944, 
    18.23944, 18.23943, 18.23943, 18.23943, 18.23944, 18.23943, 18.23944, 
    18.23944, 18.23947, 18.23948, 18.23949, 18.23949, 18.2395, 18.23949, 
    18.2395, 18.23949, 18.23949, 18.23949, 18.23948, 18.23948, 18.23945, 
    18.23947, 18.23944, 18.23944, 18.23944, 18.23944, 18.23943, 18.23944, 
    18.23943, 18.23942, 18.23943, 18.23942, 18.23944, 18.23943, 18.23949, 
    18.23949, 18.23949, 18.23949, 18.23949, 18.2395, 18.2395, 18.23949, 
    18.23949, 18.23948, 18.23948, 18.23947, 18.23946, 18.23945, 18.23944, 
    18.23944, 18.23944, 18.23944, 18.23944, 18.23944, 18.23942, 18.23944, 
    18.23942, 18.23942, 18.23943, 18.23942, 18.23949, 18.23949, 18.2395, 
    18.23949, 18.2395, 18.2395, 18.23949, 18.23948, 18.23948, 18.23948, 
    18.23947, 18.23947, 18.23945, 18.23944, 18.23944, 18.23944, 18.23944, 
    18.23943, 18.23944, 18.23943, 18.23943, 18.23944, 18.23942, 18.23942, 
    18.23942, 18.23942, 18.23949, 18.23949, 18.23949, 18.23948, 18.23949, 
    18.23948, 18.23947, 18.23946, 18.23947, 18.23945, 18.23946, 18.23946, 
    18.23945, 18.23946, 18.23944, 18.23946, 18.23943, 18.23945, 18.23943, 
    18.23944, 18.23943, 18.23943, 18.23942, 18.23941, 18.23942, 18.23941, 
    18.23948, 18.23948, 18.23948, 18.23947, 18.23947, 18.23946, 18.23945, 
    18.23946, 18.23945, 18.23945, 18.23946, 18.23945, 18.23948, 18.23947, 
    18.23947, 18.23948, 18.23945, 18.23947, 18.23944, 18.23945, 18.23943, 
    18.23944, 18.23942, 18.23941, 18.2394, 18.23939, 18.23948, 18.23948, 
    18.23947, 18.23947, 18.23946, 18.23945, 18.23945, 18.23945, 18.23944, 
    18.23944, 18.23945, 18.23944, 18.23947, 18.23945, 18.23948, 18.23947, 
    18.23947, 18.23947, 18.23946, 18.23945, 18.23944, 18.23945, 18.23941, 
    18.23943, 18.23938, 18.2394, 18.23948, 18.23948, 18.23946, 18.23947, 
    18.23945, 18.23944, 18.23944, 18.23944, 18.23944, 18.23943, 18.23944, 
    18.23943, 18.23945, 18.23944, 18.23946, 18.23946, 18.23946, 18.23946, 
    18.23945, 18.23945, 18.23945, 18.23944, 18.23944, 18.23945, 18.23941, 
    18.23943, 18.23947, 18.23946, 18.23946, 18.23947, 18.23944, 18.23945, 
    18.23943, 18.23944, 18.23943, 18.23943, 18.23944, 18.23944, 18.23944, 
    18.23945, 18.23946, 18.23946, 18.23946, 18.23946, 18.23945, 18.23944, 
    18.23944, 18.23943, 18.23945, 18.23944, 18.23944, 18.23944, 18.23946, 
    18.23944, 18.23946, 18.23946, 18.23945, 18.23944, 18.23944, 18.23944, 
    18.23944, 18.23944, 18.23945, 18.23945, 18.23945, 18.23946, 18.23946, 
    18.23946, 18.23945, 18.23944, 18.23944, 18.23943, 18.23943, 18.23941, 
    18.23942, 18.23941, 18.23942, 18.2394, 18.23944, 18.23942, 18.23945, 
    18.23945, 18.23944, 18.23943, 18.23944, 18.23943, 18.23945, 18.23946, 
    18.23946, 18.23946, 18.23946, 18.23946, 18.23945, 18.23946, 18.23944, 
    18.23945, 18.23944, 18.23943, 18.23941, 18.2394, 18.23939, 18.23938, 
    18.23938, 18.23938 ;

 TOTCOLCH4 =
  1.320662e-05, 1.302441e-05, 1.30598e-05, 1.291305e-05, 1.299444e-05, 
    1.289838e-05, 1.316966e-05, 1.301717e-05, 1.311449e-05, 1.319022e-05, 
    1.262899e-05, 1.290651e-05, 1.234188e-05, 1.251807e-05, 1.207633e-05, 
    1.236926e-05, 1.201742e-05, 1.208479e-05, 1.188229e-05, 1.194024e-05, 
    1.168187e-05, 1.185556e-05, 1.154839e-05, 1.172332e-05, 1.169591e-05, 
    1.18613e-05, 1.285061e-05, 1.266348e-05, 1.28617e-05, 1.283499e-05, 
    1.284698e-05, 1.299275e-05, 1.306628e-05, 1.322058e-05, 1.319255e-05, 
    1.307924e-05, 1.282298e-05, 1.29099e-05, 1.269108e-05, 1.269601e-05, 
    1.24531e-05, 1.256253e-05, 1.215546e-05, 1.227093e-05, 1.193782e-05, 
    1.202143e-05, 1.194174e-05, 1.19659e-05, 1.194143e-05, 1.20641e-05, 
    1.201151e-05, 1.211957e-05, 1.254202e-05, 1.24176e-05, 1.278927e-05, 
    1.301357e-05, 1.316296e-05, 1.32691e-05, 1.325409e-05, 1.322547e-05, 
    1.307858e-05, 1.294073e-05, 1.283583e-05, 1.276573e-05, 1.269672e-05, 
    1.248816e-05, 1.237807e-05, 1.213213e-05, 1.217647e-05, 1.210138e-05, 
    1.202976e-05, 1.190965e-05, 1.192941e-05, 1.187654e-05, 1.210338e-05, 
    1.195253e-05, 1.220173e-05, 1.213348e-05, 1.267789e-05, 1.288644e-05, 
    1.297518e-05, 1.3053e-05, 1.324255e-05, 1.31116e-05, 1.316319e-05, 
    1.304051e-05, 1.296264e-05, 1.300115e-05, 1.276381e-05, 1.2856e-05, 
    1.237155e-05, 1.257984e-05, 1.203811e-05, 1.216737e-05, 1.200717e-05, 
    1.208887e-05, 1.194893e-05, 1.207486e-05, 1.185689e-05, 1.180951e-05, 
    1.184188e-05, 1.171765e-05, 1.208185e-05, 1.194173e-05, 1.300223e-05, 
    1.299594e-05, 1.296669e-05, 1.309535e-05, 1.310323e-05, 1.322134e-05, 
    1.311625e-05, 1.307153e-05, 1.295814e-05, 1.289113e-05, 1.282748e-05, 
    1.268773e-05, 1.253194e-05, 1.231466e-05, 1.215898e-05, 1.205482e-05, 
    1.211867e-05, 1.206229e-05, 1.212532e-05, 1.215489e-05, 1.182725e-05, 
    1.201102e-05, 1.17355e-05, 1.175072e-05, 1.187528e-05, 1.174901e-05, 
    1.299153e-05, 1.302769e-05, 1.31533e-05, 1.305498e-05, 1.323422e-05, 
    1.313383e-05, 1.307616e-05, 1.285405e-05, 1.280535e-05, 1.27602e-05, 
    1.267111e-05, 1.255692e-05, 1.235702e-05, 1.218356e-05, 1.20256e-05, 
    1.203716e-05, 1.203309e-05, 1.199784e-05, 1.208518e-05, 1.198351e-05, 
    1.196646e-05, 1.201105e-05, 1.175276e-05, 1.182645e-05, 1.175104e-05, 
    1.179901e-05, 1.301594e-05, 1.295513e-05, 1.298798e-05, 1.292621e-05, 
    1.296971e-05, 1.277641e-05, 1.271854e-05, 1.244839e-05, 1.255916e-05, 
    1.238296e-05, 1.254125e-05, 1.251318e-05, 1.237719e-05, 1.25327e-05, 
    1.21931e-05, 1.242313e-05, 1.199647e-05, 1.22255e-05, 1.198214e-05, 
    1.202628e-05, 1.195323e-05, 1.188786e-05, 1.180573e-05, 1.165444e-05, 
    1.168944e-05, 1.156315e-05, 1.286456e-05, 1.278583e-05, 1.279278e-05, 
    1.271048e-05, 1.264966e-05, 1.251804e-05, 1.23074e-05, 1.238655e-05, 
    1.224134e-05, 1.221222e-05, 1.243286e-05, 1.229729e-05, 1.27332e-05, 
    1.266259e-05, 1.270463e-05, 1.285834e-05, 1.236828e-05, 1.261937e-05, 
    1.215641e-05, 1.229193e-05, 1.189717e-05, 1.209319e-05, 1.170872e-05, 
    1.154502e-05, 1.139144e-05, 1.121238e-05, 1.274292e-05, 1.279637e-05, 
    1.27007e-05, 1.25685e-05, 1.244609e-05, 1.228365e-05, 1.226706e-05, 
    1.223667e-05, 1.215804e-05, 1.209198e-05, 1.222705e-05, 1.207544e-05, 
    1.264618e-05, 1.234653e-05, 1.281657e-05, 1.267471e-05, 1.257629e-05, 
    1.261947e-05, 1.23956e-05, 1.234293e-05, 1.21293e-05, 1.223967e-05, 
    1.158537e-05, 1.187403e-05, 1.107648e-05, 1.129827e-05, 1.281505e-05, 
    1.274311e-05, 1.249322e-05, 1.261202e-05, 1.227283e-05, 1.218957e-05, 
    1.212198e-05, 1.203565e-05, 1.202635e-05, 1.197526e-05, 1.2059e-05, 
    1.197857e-05, 1.22833e-05, 1.214696e-05, 1.252176e-05, 1.243035e-05, 
    1.247239e-05, 1.251853e-05, 1.237623e-05, 1.222492e-05, 1.222171e-05, 
    1.217326e-05, 1.203686e-05, 1.227146e-05, 1.154816e-05, 1.199386e-05, 
    1.266473e-05, 1.252645e-05, 1.250675e-05, 1.256027e-05, 1.219792e-05, 
    1.2329e-05, 1.197651e-05, 1.20716e-05, 1.191587e-05, 1.199321e-05, 
    1.200459e-05, 1.210407e-05, 1.216608e-05, 1.232297e-05, 1.24509e-05, 
    1.255251e-05, 1.252887e-05, 1.24173e-05, 1.221568e-05, 1.20255e-05, 
    1.206711e-05, 1.19277e-05, 1.229737e-05, 1.21421e-05, 1.220206e-05, 
    1.204583e-05, 1.238864e-05, 1.209653e-05, 1.24635e-05, 1.243125e-05, 
    1.23316e-05, 1.213156e-05, 1.208742e-05, 1.204028e-05, 1.206937e-05, 
    1.221057e-05, 1.223374e-05, 1.233403e-05, 1.236173e-05, 1.243827e-05, 
    1.250169e-05, 1.244374e-05, 1.238292e-05, 1.221052e-05, 1.205551e-05, 
    1.188692e-05, 1.184574e-05, 1.164938e-05, 1.180914e-05, 1.154568e-05, 
    1.176955e-05, 1.138257e-05, 1.207968e-05, 1.17762e-05, 1.232708e-05, 
    1.226752e-05, 1.21599e-05, 1.191377e-05, 1.204656e-05, 1.18913e-05, 
    1.223465e-05, 1.241344e-05, 1.24598e-05, 1.254632e-05, 1.245782e-05, 
    1.246502e-05, 1.238042e-05, 1.24076e-05, 1.220481e-05, 1.231367e-05, 
    1.200487e-05, 1.189253e-05, 1.157636e-05, 1.138333e-05, 1.118752e-05, 
    1.110128e-05, 1.107506e-05, 1.10641e-05 ;

 TOTCOLN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTECOSYSC =
  18.2395, 18.23949, 18.23949, 18.23948, 18.23949, 18.23948, 18.2395, 
    18.23949, 18.2395, 18.2395, 18.23947, 18.23948, 18.23945, 18.23946, 
    18.23944, 18.23945, 18.23944, 18.23944, 18.23943, 18.23943, 18.23942, 
    18.23943, 18.23941, 18.23942, 18.23942, 18.23943, 18.23948, 18.23947, 
    18.23948, 18.23948, 18.23948, 18.23949, 18.23949, 18.2395, 18.2395, 
    18.23949, 18.23948, 18.23948, 18.23947, 18.23947, 18.23946, 18.23947, 
    18.23944, 18.23945, 18.23943, 18.23944, 18.23943, 18.23943, 18.23943, 
    18.23944, 18.23944, 18.23944, 18.23946, 18.23946, 18.23948, 18.23949, 
    18.2395, 18.2395, 18.2395, 18.2395, 18.23949, 18.23949, 18.23948, 
    18.23948, 18.23947, 18.23946, 18.23945, 18.23944, 18.23944, 18.23944, 
    18.23944, 18.23943, 18.23943, 18.23943, 18.23944, 18.23943, 18.23944, 
    18.23944, 18.23947, 18.23948, 18.23949, 18.23949, 18.2395, 18.23949, 
    18.2395, 18.23949, 18.23949, 18.23949, 18.23948, 18.23948, 18.23945, 
    18.23947, 18.23944, 18.23944, 18.23944, 18.23944, 18.23943, 18.23944, 
    18.23943, 18.23942, 18.23943, 18.23942, 18.23944, 18.23943, 18.23949, 
    18.23949, 18.23949, 18.23949, 18.23949, 18.2395, 18.2395, 18.23949, 
    18.23949, 18.23948, 18.23948, 18.23947, 18.23946, 18.23945, 18.23944, 
    18.23944, 18.23944, 18.23944, 18.23944, 18.23944, 18.23942, 18.23944, 
    18.23942, 18.23942, 18.23943, 18.23942, 18.23949, 18.23949, 18.2395, 
    18.23949, 18.2395, 18.2395, 18.23949, 18.23948, 18.23948, 18.23948, 
    18.23947, 18.23947, 18.23945, 18.23944, 18.23944, 18.23944, 18.23944, 
    18.23943, 18.23944, 18.23943, 18.23943, 18.23944, 18.23942, 18.23942, 
    18.23942, 18.23942, 18.23949, 18.23949, 18.23949, 18.23948, 18.23949, 
    18.23948, 18.23947, 18.23946, 18.23947, 18.23945, 18.23946, 18.23946, 
    18.23945, 18.23946, 18.23944, 18.23946, 18.23943, 18.23945, 18.23943, 
    18.23944, 18.23943, 18.23943, 18.23942, 18.23941, 18.23942, 18.23941, 
    18.23948, 18.23948, 18.23948, 18.23947, 18.23947, 18.23946, 18.23945, 
    18.23946, 18.23945, 18.23945, 18.23946, 18.23945, 18.23948, 18.23947, 
    18.23947, 18.23948, 18.23945, 18.23947, 18.23944, 18.23945, 18.23943, 
    18.23944, 18.23942, 18.23941, 18.2394, 18.23939, 18.23948, 18.23948, 
    18.23947, 18.23947, 18.23946, 18.23945, 18.23945, 18.23945, 18.23944, 
    18.23944, 18.23945, 18.23944, 18.23947, 18.23945, 18.23948, 18.23947, 
    18.23947, 18.23947, 18.23946, 18.23945, 18.23944, 18.23945, 18.23941, 
    18.23943, 18.23938, 18.2394, 18.23948, 18.23948, 18.23946, 18.23947, 
    18.23945, 18.23944, 18.23944, 18.23944, 18.23944, 18.23943, 18.23944, 
    18.23943, 18.23945, 18.23944, 18.23946, 18.23946, 18.23946, 18.23946, 
    18.23945, 18.23945, 18.23945, 18.23944, 18.23944, 18.23945, 18.23941, 
    18.23943, 18.23947, 18.23946, 18.23946, 18.23947, 18.23944, 18.23945, 
    18.23943, 18.23944, 18.23943, 18.23943, 18.23944, 18.23944, 18.23944, 
    18.23945, 18.23946, 18.23946, 18.23946, 18.23946, 18.23945, 18.23944, 
    18.23944, 18.23943, 18.23945, 18.23944, 18.23944, 18.23944, 18.23946, 
    18.23944, 18.23946, 18.23946, 18.23945, 18.23944, 18.23944, 18.23944, 
    18.23944, 18.23944, 18.23945, 18.23945, 18.23945, 18.23946, 18.23946, 
    18.23946, 18.23945, 18.23944, 18.23944, 18.23943, 18.23943, 18.23941, 
    18.23942, 18.23941, 18.23942, 18.2394, 18.23944, 18.23942, 18.23945, 
    18.23945, 18.23944, 18.23943, 18.23944, 18.23943, 18.23945, 18.23946, 
    18.23946, 18.23946, 18.23946, 18.23946, 18.23945, 18.23946, 18.23944, 
    18.23945, 18.23944, 18.23943, 18.23941, 18.2394, 18.23939, 18.23938, 
    18.23938, 18.23938 ;

 TOTECOSYSN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTLITC =
  5.976081e-05, 5.976067e-05, 5.97607e-05, 5.976058e-05, 5.976064e-05, 
    5.976057e-05, 5.976078e-05, 5.976066e-05, 5.976074e-05, 5.97608e-05, 
    5.976036e-05, 5.976058e-05, 5.976013e-05, 5.976027e-05, 5.975992e-05, 
    5.976015e-05, 5.975987e-05, 5.975992e-05, 5.975976e-05, 5.975981e-05, 
    5.97596e-05, 5.975974e-05, 5.97595e-05, 5.975964e-05, 5.975962e-05, 
    5.975975e-05, 5.976053e-05, 5.976038e-05, 5.976054e-05, 5.976052e-05, 
    5.976053e-05, 5.976064e-05, 5.97607e-05, 5.976082e-05, 5.97608e-05, 
    5.976071e-05, 5.976051e-05, 5.976058e-05, 5.97604e-05, 5.976041e-05, 
    5.976022e-05, 5.97603e-05, 5.975998e-05, 5.976007e-05, 5.975981e-05, 
    5.975987e-05, 5.975981e-05, 5.975983e-05, 5.975981e-05, 5.975991e-05, 
    5.975987e-05, 5.975995e-05, 5.976029e-05, 5.976019e-05, 5.976048e-05, 
    5.976066e-05, 5.976078e-05, 5.976086e-05, 5.976085e-05, 5.976083e-05, 
    5.976071e-05, 5.97606e-05, 5.976052e-05, 5.976046e-05, 5.976041e-05, 
    5.976024e-05, 5.976016e-05, 5.975996e-05, 5.976e-05, 5.975994e-05, 
    5.975988e-05, 5.975979e-05, 5.97598e-05, 5.975976e-05, 5.975994e-05, 
    5.975982e-05, 5.976002e-05, 5.975996e-05, 5.976039e-05, 5.976056e-05, 
    5.976063e-05, 5.976069e-05, 5.976084e-05, 5.976074e-05, 5.976078e-05, 
    5.976068e-05, 5.976062e-05, 5.976065e-05, 5.976046e-05, 5.976054e-05, 
    5.976015e-05, 5.976032e-05, 5.975989e-05, 5.975999e-05, 5.975986e-05, 
    5.975993e-05, 5.975982e-05, 5.975992e-05, 5.975974e-05, 5.975971e-05, 
    5.975973e-05, 5.975963e-05, 5.975992e-05, 5.975981e-05, 5.976065e-05, 
    5.976064e-05, 5.976062e-05, 5.976072e-05, 5.976073e-05, 5.976082e-05, 
    5.976074e-05, 5.97607e-05, 5.976062e-05, 5.976056e-05, 5.976051e-05, 
    5.97604e-05, 5.976028e-05, 5.976011e-05, 5.975998e-05, 5.97599e-05, 
    5.975995e-05, 5.975991e-05, 5.975996e-05, 5.975998e-05, 5.975972e-05, 
    5.975987e-05, 5.975965e-05, 5.975966e-05, 5.975976e-05, 5.975966e-05, 
    5.976064e-05, 5.976067e-05, 5.976077e-05, 5.976069e-05, 5.976083e-05, 
    5.976075e-05, 5.976071e-05, 5.976053e-05, 5.97605e-05, 5.976046e-05, 
    5.976039e-05, 5.97603e-05, 5.976014e-05, 5.976e-05, 5.975988e-05, 
    5.975989e-05, 5.975988e-05, 5.975986e-05, 5.975992e-05, 5.975984e-05, 
    5.975983e-05, 5.975987e-05, 5.975966e-05, 5.975972e-05, 5.975966e-05, 
    5.97597e-05, 5.976066e-05, 5.976061e-05, 5.976064e-05, 5.976059e-05, 
    5.976062e-05, 5.976047e-05, 5.976043e-05, 5.976021e-05, 5.97603e-05, 
    5.976016e-05, 5.976028e-05, 5.976026e-05, 5.976016e-05, 5.976028e-05, 
    5.976001e-05, 5.976019e-05, 5.975986e-05, 5.976004e-05, 5.975984e-05, 
    5.975988e-05, 5.975982e-05, 5.975977e-05, 5.97597e-05, 5.975958e-05, 
    5.975961e-05, 5.975951e-05, 5.976054e-05, 5.976048e-05, 5.976048e-05, 
    5.976042e-05, 5.976037e-05, 5.976027e-05, 5.97601e-05, 5.976016e-05, 
    5.976005e-05, 5.976003e-05, 5.97602e-05, 5.976009e-05, 5.976044e-05, 
    5.976038e-05, 5.976042e-05, 5.976054e-05, 5.976015e-05, 5.976035e-05, 
    5.975998e-05, 5.976009e-05, 5.975978e-05, 5.975993e-05, 5.975963e-05, 
    5.97595e-05, 5.975938e-05, 5.975923e-05, 5.976044e-05, 5.976049e-05, 
    5.976041e-05, 5.976031e-05, 5.976021e-05, 5.976008e-05, 5.976007e-05, 
    5.976004e-05, 5.975998e-05, 5.975993e-05, 5.976004e-05, 5.975992e-05, 
    5.976037e-05, 5.976013e-05, 5.97605e-05, 5.976039e-05, 5.976031e-05, 
    5.976035e-05, 5.976017e-05, 5.976013e-05, 5.975996e-05, 5.976005e-05, 
    5.975953e-05, 5.975976e-05, 5.975912e-05, 5.97593e-05, 5.97605e-05, 
    5.976044e-05, 5.976025e-05, 5.976034e-05, 5.976007e-05, 5.976001e-05, 
    5.975995e-05, 5.975988e-05, 5.975988e-05, 5.975984e-05, 5.975991e-05, 
    5.975984e-05, 5.976008e-05, 5.975998e-05, 5.976027e-05, 5.97602e-05, 
    5.976023e-05, 5.976027e-05, 5.976016e-05, 5.976004e-05, 5.976003e-05, 
    5.975999e-05, 5.975989e-05, 5.976007e-05, 5.97595e-05, 5.975985e-05, 
    5.976038e-05, 5.976027e-05, 5.976026e-05, 5.97603e-05, 5.976002e-05, 
    5.976012e-05, 5.975984e-05, 5.975991e-05, 5.975979e-05, 5.975985e-05, 
    5.975986e-05, 5.975994e-05, 5.975999e-05, 5.976011e-05, 5.976022e-05, 
    5.97603e-05, 5.976028e-05, 5.976019e-05, 5.976003e-05, 5.975988e-05, 
    5.975991e-05, 5.97598e-05, 5.976009e-05, 5.975997e-05, 5.976002e-05, 
    5.97599e-05, 5.976016e-05, 5.975994e-05, 5.976023e-05, 5.97602e-05, 
    5.976012e-05, 5.975996e-05, 5.975993e-05, 5.975989e-05, 5.975991e-05, 
    5.976003e-05, 5.976004e-05, 5.976012e-05, 5.976014e-05, 5.97602e-05, 
    5.976026e-05, 5.976021e-05, 5.976016e-05, 5.976003e-05, 5.97599e-05, 
    5.975977e-05, 5.975974e-05, 5.975958e-05, 5.975971e-05, 5.97595e-05, 
    5.975968e-05, 5.975937e-05, 5.975992e-05, 5.975968e-05, 5.976012e-05, 
    5.976007e-05, 5.975999e-05, 5.975979e-05, 5.97599e-05, 5.975977e-05, 
    5.976004e-05, 5.976019e-05, 5.976022e-05, 5.976029e-05, 5.976022e-05, 
    5.976023e-05, 5.976016e-05, 5.976018e-05, 5.976002e-05, 5.976011e-05, 
    5.975986e-05, 5.975977e-05, 5.975952e-05, 5.975937e-05, 5.975921e-05, 
    5.975914e-05, 5.975912e-05, 5.975911e-05 ;

 TOTLITC_1m =
  5.976081e-05, 5.976067e-05, 5.97607e-05, 5.976058e-05, 5.976064e-05, 
    5.976057e-05, 5.976078e-05, 5.976066e-05, 5.976074e-05, 5.97608e-05, 
    5.976036e-05, 5.976058e-05, 5.976013e-05, 5.976027e-05, 5.975992e-05, 
    5.976015e-05, 5.975987e-05, 5.975992e-05, 5.975976e-05, 5.975981e-05, 
    5.97596e-05, 5.975974e-05, 5.97595e-05, 5.975964e-05, 5.975962e-05, 
    5.975975e-05, 5.976053e-05, 5.976038e-05, 5.976054e-05, 5.976052e-05, 
    5.976053e-05, 5.976064e-05, 5.97607e-05, 5.976082e-05, 5.97608e-05, 
    5.976071e-05, 5.976051e-05, 5.976058e-05, 5.97604e-05, 5.976041e-05, 
    5.976022e-05, 5.97603e-05, 5.975998e-05, 5.976007e-05, 5.975981e-05, 
    5.975987e-05, 5.975981e-05, 5.975983e-05, 5.975981e-05, 5.975991e-05, 
    5.975987e-05, 5.975995e-05, 5.976029e-05, 5.976019e-05, 5.976048e-05, 
    5.976066e-05, 5.976078e-05, 5.976086e-05, 5.976085e-05, 5.976083e-05, 
    5.976071e-05, 5.97606e-05, 5.976052e-05, 5.976046e-05, 5.976041e-05, 
    5.976024e-05, 5.976016e-05, 5.975996e-05, 5.976e-05, 5.975994e-05, 
    5.975988e-05, 5.975979e-05, 5.97598e-05, 5.975976e-05, 5.975994e-05, 
    5.975982e-05, 5.976002e-05, 5.975996e-05, 5.976039e-05, 5.976056e-05, 
    5.976063e-05, 5.976069e-05, 5.976084e-05, 5.976074e-05, 5.976078e-05, 
    5.976068e-05, 5.976062e-05, 5.976065e-05, 5.976046e-05, 5.976054e-05, 
    5.976015e-05, 5.976032e-05, 5.975989e-05, 5.975999e-05, 5.975986e-05, 
    5.975993e-05, 5.975982e-05, 5.975992e-05, 5.975974e-05, 5.975971e-05, 
    5.975973e-05, 5.975963e-05, 5.975992e-05, 5.975981e-05, 5.976065e-05, 
    5.976064e-05, 5.976062e-05, 5.976072e-05, 5.976073e-05, 5.976082e-05, 
    5.976074e-05, 5.97607e-05, 5.976062e-05, 5.976056e-05, 5.976051e-05, 
    5.97604e-05, 5.976028e-05, 5.976011e-05, 5.975998e-05, 5.97599e-05, 
    5.975995e-05, 5.975991e-05, 5.975996e-05, 5.975998e-05, 5.975972e-05, 
    5.975987e-05, 5.975965e-05, 5.975966e-05, 5.975976e-05, 5.975966e-05, 
    5.976064e-05, 5.976067e-05, 5.976077e-05, 5.976069e-05, 5.976083e-05, 
    5.976075e-05, 5.976071e-05, 5.976053e-05, 5.97605e-05, 5.976046e-05, 
    5.976039e-05, 5.97603e-05, 5.976014e-05, 5.976e-05, 5.975988e-05, 
    5.975989e-05, 5.975988e-05, 5.975986e-05, 5.975992e-05, 5.975984e-05, 
    5.975983e-05, 5.975987e-05, 5.975966e-05, 5.975972e-05, 5.975966e-05, 
    5.97597e-05, 5.976066e-05, 5.976061e-05, 5.976064e-05, 5.976059e-05, 
    5.976062e-05, 5.976047e-05, 5.976043e-05, 5.976021e-05, 5.97603e-05, 
    5.976016e-05, 5.976028e-05, 5.976026e-05, 5.976016e-05, 5.976028e-05, 
    5.976001e-05, 5.976019e-05, 5.975986e-05, 5.976004e-05, 5.975984e-05, 
    5.975988e-05, 5.975982e-05, 5.975977e-05, 5.97597e-05, 5.975958e-05, 
    5.975961e-05, 5.975951e-05, 5.976054e-05, 5.976048e-05, 5.976048e-05, 
    5.976042e-05, 5.976037e-05, 5.976027e-05, 5.97601e-05, 5.976016e-05, 
    5.976005e-05, 5.976003e-05, 5.97602e-05, 5.976009e-05, 5.976044e-05, 
    5.976038e-05, 5.976042e-05, 5.976054e-05, 5.976015e-05, 5.976035e-05, 
    5.975998e-05, 5.976009e-05, 5.975978e-05, 5.975993e-05, 5.975963e-05, 
    5.97595e-05, 5.975938e-05, 5.975923e-05, 5.976044e-05, 5.976049e-05, 
    5.976041e-05, 5.976031e-05, 5.976021e-05, 5.976008e-05, 5.976007e-05, 
    5.976004e-05, 5.975998e-05, 5.975993e-05, 5.976004e-05, 5.975992e-05, 
    5.976037e-05, 5.976013e-05, 5.97605e-05, 5.976039e-05, 5.976031e-05, 
    5.976035e-05, 5.976017e-05, 5.976013e-05, 5.975996e-05, 5.976005e-05, 
    5.975953e-05, 5.975976e-05, 5.975912e-05, 5.97593e-05, 5.97605e-05, 
    5.976044e-05, 5.976025e-05, 5.976034e-05, 5.976007e-05, 5.976001e-05, 
    5.975995e-05, 5.975988e-05, 5.975988e-05, 5.975984e-05, 5.975991e-05, 
    5.975984e-05, 5.976008e-05, 5.975998e-05, 5.976027e-05, 5.97602e-05, 
    5.976023e-05, 5.976027e-05, 5.976016e-05, 5.976004e-05, 5.976003e-05, 
    5.975999e-05, 5.975989e-05, 5.976007e-05, 5.97595e-05, 5.975985e-05, 
    5.976038e-05, 5.976027e-05, 5.976026e-05, 5.97603e-05, 5.976002e-05, 
    5.976012e-05, 5.975984e-05, 5.975991e-05, 5.975979e-05, 5.975985e-05, 
    5.975986e-05, 5.975994e-05, 5.975999e-05, 5.976011e-05, 5.976022e-05, 
    5.97603e-05, 5.976028e-05, 5.976019e-05, 5.976003e-05, 5.975988e-05, 
    5.975991e-05, 5.97598e-05, 5.976009e-05, 5.975997e-05, 5.976002e-05, 
    5.97599e-05, 5.976016e-05, 5.975994e-05, 5.976023e-05, 5.97602e-05, 
    5.976012e-05, 5.975996e-05, 5.975993e-05, 5.975989e-05, 5.975991e-05, 
    5.976003e-05, 5.976004e-05, 5.976012e-05, 5.976014e-05, 5.97602e-05, 
    5.976026e-05, 5.976021e-05, 5.976016e-05, 5.976003e-05, 5.97599e-05, 
    5.975977e-05, 5.975974e-05, 5.975958e-05, 5.975971e-05, 5.97595e-05, 
    5.975968e-05, 5.975937e-05, 5.975992e-05, 5.975968e-05, 5.976012e-05, 
    5.976007e-05, 5.975999e-05, 5.975979e-05, 5.97599e-05, 5.975977e-05, 
    5.976004e-05, 5.976019e-05, 5.976022e-05, 5.976029e-05, 5.976022e-05, 
    5.976023e-05, 5.976016e-05, 5.976018e-05, 5.976002e-05, 5.976011e-05, 
    5.975986e-05, 5.975977e-05, 5.975952e-05, 5.975937e-05, 5.975921e-05, 
    5.975914e-05, 5.975912e-05, 5.975911e-05 ;

 TOTLITN =
  1.375895e-06, 1.375891e-06, 1.375891e-06, 1.375888e-06, 1.37589e-06, 
    1.375888e-06, 1.375894e-06, 1.375891e-06, 1.375893e-06, 1.375894e-06, 
    1.375882e-06, 1.375888e-06, 1.375876e-06, 1.375879e-06, 1.37587e-06, 
    1.375876e-06, 1.375868e-06, 1.37587e-06, 1.375865e-06, 1.375867e-06, 
    1.375861e-06, 1.375865e-06, 1.375858e-06, 1.375862e-06, 1.375861e-06, 
    1.375865e-06, 1.375887e-06, 1.375883e-06, 1.375887e-06, 1.375886e-06, 
    1.375887e-06, 1.37589e-06, 1.375892e-06, 1.375895e-06, 1.375894e-06, 
    1.375892e-06, 1.375886e-06, 1.375888e-06, 1.375883e-06, 1.375883e-06, 
    1.375878e-06, 1.37588e-06, 1.375871e-06, 1.375874e-06, 1.375867e-06, 
    1.375868e-06, 1.375867e-06, 1.375867e-06, 1.375867e-06, 1.375869e-06, 
    1.375868e-06, 1.375871e-06, 1.37588e-06, 1.375877e-06, 1.375885e-06, 
    1.37589e-06, 1.375894e-06, 1.375896e-06, 1.375896e-06, 1.375895e-06, 
    1.375892e-06, 1.375889e-06, 1.375886e-06, 1.375885e-06, 1.375883e-06, 
    1.375879e-06, 1.375876e-06, 1.375871e-06, 1.375872e-06, 1.37587e-06, 
    1.375869e-06, 1.375866e-06, 1.375866e-06, 1.375865e-06, 1.37587e-06, 
    1.375867e-06, 1.375872e-06, 1.375871e-06, 1.375883e-06, 1.375888e-06, 
    1.37589e-06, 1.375891e-06, 1.375896e-06, 1.375893e-06, 1.375894e-06, 
    1.375891e-06, 1.375889e-06, 1.37589e-06, 1.375885e-06, 1.375887e-06, 
    1.375876e-06, 1.375881e-06, 1.375869e-06, 1.375872e-06, 1.375868e-06, 
    1.37587e-06, 1.375867e-06, 1.375869e-06, 1.375865e-06, 1.375864e-06, 
    1.375864e-06, 1.375862e-06, 1.37587e-06, 1.375867e-06, 1.37589e-06, 
    1.37589e-06, 1.375889e-06, 1.375892e-06, 1.375892e-06, 1.375895e-06, 
    1.375893e-06, 1.375892e-06, 1.375889e-06, 1.375888e-06, 1.375886e-06, 
    1.375883e-06, 1.37588e-06, 1.375875e-06, 1.375871e-06, 1.375869e-06, 
    1.375871e-06, 1.375869e-06, 1.375871e-06, 1.375871e-06, 1.375864e-06, 
    1.375868e-06, 1.375862e-06, 1.375862e-06, 1.375865e-06, 1.375862e-06, 
    1.37589e-06, 1.375891e-06, 1.375893e-06, 1.375891e-06, 1.375895e-06, 
    1.375893e-06, 1.375892e-06, 1.375887e-06, 1.375886e-06, 1.375885e-06, 
    1.375883e-06, 1.37588e-06, 1.375876e-06, 1.375872e-06, 1.375868e-06, 
    1.375869e-06, 1.375869e-06, 1.375868e-06, 1.37587e-06, 1.375868e-06, 
    1.375867e-06, 1.375868e-06, 1.375862e-06, 1.375864e-06, 1.375862e-06, 
    1.375863e-06, 1.375891e-06, 1.375889e-06, 1.37589e-06, 1.375888e-06, 
    1.375889e-06, 1.375885e-06, 1.375884e-06, 1.375878e-06, 1.37588e-06, 
    1.375876e-06, 1.37588e-06, 1.375879e-06, 1.375876e-06, 1.37588e-06, 
    1.375872e-06, 1.375877e-06, 1.375868e-06, 1.375873e-06, 1.375867e-06, 
    1.375868e-06, 1.375867e-06, 1.375865e-06, 1.375864e-06, 1.37586e-06, 
    1.375861e-06, 1.375858e-06, 1.375887e-06, 1.375885e-06, 1.375886e-06, 
    1.375884e-06, 1.375882e-06, 1.375879e-06, 1.375875e-06, 1.375877e-06, 
    1.375873e-06, 1.375873e-06, 1.375878e-06, 1.375874e-06, 1.375884e-06, 
    1.375883e-06, 1.375884e-06, 1.375887e-06, 1.375876e-06, 1.375882e-06, 
    1.375871e-06, 1.375874e-06, 1.375866e-06, 1.37587e-06, 1.375861e-06, 
    1.375858e-06, 1.375854e-06, 1.37585e-06, 1.375884e-06, 1.375886e-06, 
    1.375883e-06, 1.375881e-06, 1.375878e-06, 1.375874e-06, 1.375874e-06, 
    1.375873e-06, 1.375871e-06, 1.37587e-06, 1.375873e-06, 1.37587e-06, 
    1.375882e-06, 1.375876e-06, 1.375886e-06, 1.375883e-06, 1.375881e-06, 
    1.375882e-06, 1.375877e-06, 1.375876e-06, 1.375871e-06, 1.375873e-06, 
    1.375859e-06, 1.375865e-06, 1.375847e-06, 1.375852e-06, 1.375886e-06, 
    1.375884e-06, 1.375879e-06, 1.375882e-06, 1.375874e-06, 1.375872e-06, 
    1.375871e-06, 1.375869e-06, 1.375868e-06, 1.375867e-06, 1.375869e-06, 
    1.375867e-06, 1.375874e-06, 1.375871e-06, 1.375879e-06, 1.375877e-06, 
    1.375878e-06, 1.375879e-06, 1.375876e-06, 1.375873e-06, 1.375873e-06, 
    1.375872e-06, 1.375869e-06, 1.375874e-06, 1.375858e-06, 1.375868e-06, 
    1.375883e-06, 1.37588e-06, 1.375879e-06, 1.37588e-06, 1.375872e-06, 
    1.375875e-06, 1.375867e-06, 1.375869e-06, 1.375866e-06, 1.375868e-06, 
    1.375868e-06, 1.37587e-06, 1.375872e-06, 1.375875e-06, 1.375878e-06, 
    1.37588e-06, 1.37588e-06, 1.375877e-06, 1.375873e-06, 1.375868e-06, 
    1.375869e-06, 1.375866e-06, 1.375874e-06, 1.375871e-06, 1.375872e-06, 
    1.375869e-06, 1.375877e-06, 1.37587e-06, 1.375878e-06, 1.375877e-06, 
    1.375875e-06, 1.375871e-06, 1.37587e-06, 1.375869e-06, 1.375869e-06, 
    1.375873e-06, 1.375873e-06, 1.375875e-06, 1.375876e-06, 1.375878e-06, 
    1.375879e-06, 1.375878e-06, 1.375876e-06, 1.375873e-06, 1.375869e-06, 
    1.375865e-06, 1.375864e-06, 1.37586e-06, 1.375864e-06, 1.375858e-06, 
    1.375863e-06, 1.375854e-06, 1.37587e-06, 1.375863e-06, 1.375875e-06, 
    1.375874e-06, 1.375871e-06, 1.375866e-06, 1.375869e-06, 1.375865e-06, 
    1.375873e-06, 1.375877e-06, 1.375878e-06, 1.37588e-06, 1.375878e-06, 
    1.375878e-06, 1.375876e-06, 1.375877e-06, 1.375872e-06, 1.375875e-06, 
    1.375868e-06, 1.375866e-06, 1.375858e-06, 1.375854e-06, 1.37585e-06, 
    1.375848e-06, 1.375847e-06, 1.375847e-06 ;

 TOTLITN_1m =
  1.375895e-06, 1.375891e-06, 1.375891e-06, 1.375888e-06, 1.37589e-06, 
    1.375888e-06, 1.375894e-06, 1.375891e-06, 1.375893e-06, 1.375894e-06, 
    1.375882e-06, 1.375888e-06, 1.375876e-06, 1.375879e-06, 1.37587e-06, 
    1.375876e-06, 1.375868e-06, 1.37587e-06, 1.375865e-06, 1.375867e-06, 
    1.375861e-06, 1.375865e-06, 1.375858e-06, 1.375862e-06, 1.375861e-06, 
    1.375865e-06, 1.375887e-06, 1.375883e-06, 1.375887e-06, 1.375886e-06, 
    1.375887e-06, 1.37589e-06, 1.375892e-06, 1.375895e-06, 1.375894e-06, 
    1.375892e-06, 1.375886e-06, 1.375888e-06, 1.375883e-06, 1.375883e-06, 
    1.375878e-06, 1.37588e-06, 1.375871e-06, 1.375874e-06, 1.375867e-06, 
    1.375868e-06, 1.375867e-06, 1.375867e-06, 1.375867e-06, 1.375869e-06, 
    1.375868e-06, 1.375871e-06, 1.37588e-06, 1.375877e-06, 1.375885e-06, 
    1.37589e-06, 1.375894e-06, 1.375896e-06, 1.375896e-06, 1.375895e-06, 
    1.375892e-06, 1.375889e-06, 1.375886e-06, 1.375885e-06, 1.375883e-06, 
    1.375879e-06, 1.375876e-06, 1.375871e-06, 1.375872e-06, 1.37587e-06, 
    1.375869e-06, 1.375866e-06, 1.375866e-06, 1.375865e-06, 1.37587e-06, 
    1.375867e-06, 1.375872e-06, 1.375871e-06, 1.375883e-06, 1.375888e-06, 
    1.37589e-06, 1.375891e-06, 1.375896e-06, 1.375893e-06, 1.375894e-06, 
    1.375891e-06, 1.375889e-06, 1.37589e-06, 1.375885e-06, 1.375887e-06, 
    1.375876e-06, 1.375881e-06, 1.375869e-06, 1.375872e-06, 1.375868e-06, 
    1.37587e-06, 1.375867e-06, 1.375869e-06, 1.375865e-06, 1.375864e-06, 
    1.375864e-06, 1.375862e-06, 1.37587e-06, 1.375867e-06, 1.37589e-06, 
    1.37589e-06, 1.375889e-06, 1.375892e-06, 1.375892e-06, 1.375895e-06, 
    1.375893e-06, 1.375892e-06, 1.375889e-06, 1.375888e-06, 1.375886e-06, 
    1.375883e-06, 1.37588e-06, 1.375875e-06, 1.375871e-06, 1.375869e-06, 
    1.375871e-06, 1.375869e-06, 1.375871e-06, 1.375871e-06, 1.375864e-06, 
    1.375868e-06, 1.375862e-06, 1.375862e-06, 1.375865e-06, 1.375862e-06, 
    1.37589e-06, 1.375891e-06, 1.375893e-06, 1.375891e-06, 1.375895e-06, 
    1.375893e-06, 1.375892e-06, 1.375887e-06, 1.375886e-06, 1.375885e-06, 
    1.375883e-06, 1.37588e-06, 1.375876e-06, 1.375872e-06, 1.375868e-06, 
    1.375869e-06, 1.375869e-06, 1.375868e-06, 1.37587e-06, 1.375868e-06, 
    1.375867e-06, 1.375868e-06, 1.375862e-06, 1.375864e-06, 1.375862e-06, 
    1.375863e-06, 1.375891e-06, 1.375889e-06, 1.37589e-06, 1.375888e-06, 
    1.375889e-06, 1.375885e-06, 1.375884e-06, 1.375878e-06, 1.37588e-06, 
    1.375876e-06, 1.37588e-06, 1.375879e-06, 1.375876e-06, 1.37588e-06, 
    1.375872e-06, 1.375877e-06, 1.375868e-06, 1.375873e-06, 1.375867e-06, 
    1.375868e-06, 1.375867e-06, 1.375865e-06, 1.375864e-06, 1.37586e-06, 
    1.375861e-06, 1.375858e-06, 1.375887e-06, 1.375885e-06, 1.375886e-06, 
    1.375884e-06, 1.375882e-06, 1.375879e-06, 1.375875e-06, 1.375877e-06, 
    1.375873e-06, 1.375873e-06, 1.375878e-06, 1.375874e-06, 1.375884e-06, 
    1.375883e-06, 1.375884e-06, 1.375887e-06, 1.375876e-06, 1.375882e-06, 
    1.375871e-06, 1.375874e-06, 1.375866e-06, 1.37587e-06, 1.375861e-06, 
    1.375858e-06, 1.375854e-06, 1.37585e-06, 1.375884e-06, 1.375886e-06, 
    1.375883e-06, 1.375881e-06, 1.375878e-06, 1.375874e-06, 1.375874e-06, 
    1.375873e-06, 1.375871e-06, 1.37587e-06, 1.375873e-06, 1.37587e-06, 
    1.375882e-06, 1.375876e-06, 1.375886e-06, 1.375883e-06, 1.375881e-06, 
    1.375882e-06, 1.375877e-06, 1.375876e-06, 1.375871e-06, 1.375873e-06, 
    1.375859e-06, 1.375865e-06, 1.375847e-06, 1.375852e-06, 1.375886e-06, 
    1.375884e-06, 1.375879e-06, 1.375882e-06, 1.375874e-06, 1.375872e-06, 
    1.375871e-06, 1.375869e-06, 1.375868e-06, 1.375867e-06, 1.375869e-06, 
    1.375867e-06, 1.375874e-06, 1.375871e-06, 1.375879e-06, 1.375877e-06, 
    1.375878e-06, 1.375879e-06, 1.375876e-06, 1.375873e-06, 1.375873e-06, 
    1.375872e-06, 1.375869e-06, 1.375874e-06, 1.375858e-06, 1.375868e-06, 
    1.375883e-06, 1.37588e-06, 1.375879e-06, 1.37588e-06, 1.375872e-06, 
    1.375875e-06, 1.375867e-06, 1.375869e-06, 1.375866e-06, 1.375868e-06, 
    1.375868e-06, 1.37587e-06, 1.375872e-06, 1.375875e-06, 1.375878e-06, 
    1.37588e-06, 1.37588e-06, 1.375877e-06, 1.375873e-06, 1.375868e-06, 
    1.375869e-06, 1.375866e-06, 1.375874e-06, 1.375871e-06, 1.375872e-06, 
    1.375869e-06, 1.375877e-06, 1.37587e-06, 1.375878e-06, 1.375877e-06, 
    1.375875e-06, 1.375871e-06, 1.37587e-06, 1.375869e-06, 1.375869e-06, 
    1.375873e-06, 1.375873e-06, 1.375875e-06, 1.375876e-06, 1.375878e-06, 
    1.375879e-06, 1.375878e-06, 1.375876e-06, 1.375873e-06, 1.375869e-06, 
    1.375865e-06, 1.375864e-06, 1.37586e-06, 1.375864e-06, 1.375858e-06, 
    1.375863e-06, 1.375854e-06, 1.37587e-06, 1.375863e-06, 1.375875e-06, 
    1.375874e-06, 1.375871e-06, 1.375866e-06, 1.375869e-06, 1.375865e-06, 
    1.375873e-06, 1.375877e-06, 1.375878e-06, 1.37588e-06, 1.375878e-06, 
    1.375878e-06, 1.375876e-06, 1.375877e-06, 1.375872e-06, 1.375875e-06, 
    1.375868e-06, 1.375866e-06, 1.375858e-06, 1.375854e-06, 1.37585e-06, 
    1.375848e-06, 1.375847e-06, 1.375847e-06 ;

 TOTPFTC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTPFTN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TOTPRODC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTPRODN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTSOMC =
  17.34412, 17.34411, 17.34411, 17.3441, 17.34411, 17.3441, 17.34412, 
    17.34411, 17.34411, 17.34412, 17.34409, 17.3441, 17.34407, 17.34408, 
    17.34406, 17.34407, 17.34406, 17.34406, 17.34405, 17.34405, 17.34404, 
    17.34405, 17.34403, 17.34404, 17.34404, 17.34405, 17.3441, 17.34409, 
    17.3441, 17.3441, 17.3441, 17.34411, 17.34411, 17.34412, 17.34412, 
    17.34411, 17.3441, 17.3441, 17.34409, 17.34409, 17.34408, 17.34408, 
    17.34406, 17.34407, 17.34405, 17.34406, 17.34405, 17.34405, 17.34405, 
    17.34406, 17.34405, 17.34406, 17.34408, 17.34408, 17.3441, 17.34411, 
    17.34412, 17.34412, 17.34412, 17.34412, 17.34411, 17.3441, 17.3441, 
    17.3441, 17.34409, 17.34408, 17.34407, 17.34406, 17.34406, 17.34406, 
    17.34406, 17.34405, 17.34405, 17.34405, 17.34406, 17.34405, 17.34406, 
    17.34406, 17.34409, 17.3441, 17.34411, 17.34411, 17.34412, 17.34411, 
    17.34412, 17.34411, 17.34411, 17.34411, 17.3441, 17.3441, 17.34407, 
    17.34409, 17.34406, 17.34406, 17.34405, 17.34406, 17.34405, 17.34406, 
    17.34405, 17.34404, 17.34405, 17.34404, 17.34406, 17.34405, 17.34411, 
    17.34411, 17.34411, 17.34411, 17.34411, 17.34412, 17.34411, 17.34411, 
    17.34411, 17.3441, 17.3441, 17.34409, 17.34408, 17.34407, 17.34406, 
    17.34406, 17.34406, 17.34406, 17.34406, 17.34406, 17.34404, 17.34405, 
    17.34404, 17.34404, 17.34405, 17.34404, 17.34411, 17.34411, 17.34412, 
    17.34411, 17.34412, 17.34412, 17.34411, 17.3441, 17.3441, 17.3441, 
    17.34409, 17.34408, 17.34407, 17.34406, 17.34406, 17.34406, 17.34406, 
    17.34405, 17.34406, 17.34405, 17.34405, 17.34405, 17.34404, 17.34404, 
    17.34404, 17.34404, 17.34411, 17.34411, 17.34411, 17.3441, 17.34411, 
    17.3441, 17.34409, 17.34408, 17.34408, 17.34407, 17.34408, 17.34408, 
    17.34407, 17.34408, 17.34406, 17.34408, 17.34405, 17.34407, 17.34405, 
    17.34406, 17.34405, 17.34405, 17.34404, 17.34403, 17.34404, 17.34403, 
    17.3441, 17.3441, 17.3441, 17.34409, 17.34409, 17.34408, 17.34407, 
    17.34407, 17.34407, 17.34406, 17.34408, 17.34407, 17.34409, 17.34409, 
    17.34409, 17.3441, 17.34407, 17.34409, 17.34406, 17.34407, 17.34405, 
    17.34406, 17.34404, 17.34403, 17.34402, 17.34401, 17.3441, 17.3441, 
    17.34409, 17.34409, 17.34408, 17.34407, 17.34407, 17.34407, 17.34406, 
    17.34406, 17.34407, 17.34406, 17.34409, 17.34407, 17.3441, 17.34409, 
    17.34409, 17.34409, 17.34408, 17.34407, 17.34406, 17.34407, 17.34403, 
    17.34405, 17.344, 17.34402, 17.3441, 17.3441, 17.34408, 17.34409, 
    17.34407, 17.34406, 17.34406, 17.34406, 17.34406, 17.34405, 17.34406, 
    17.34405, 17.34407, 17.34406, 17.34408, 17.34408, 17.34408, 17.34408, 
    17.34407, 17.34407, 17.34407, 17.34406, 17.34406, 17.34407, 17.34403, 
    17.34405, 17.34409, 17.34408, 17.34408, 17.34408, 17.34406, 17.34407, 
    17.34405, 17.34406, 17.34405, 17.34405, 17.34405, 17.34406, 17.34406, 
    17.34407, 17.34408, 17.34408, 17.34408, 17.34408, 17.34406, 17.34406, 
    17.34406, 17.34405, 17.34407, 17.34406, 17.34406, 17.34406, 17.34407, 
    17.34406, 17.34408, 17.34408, 17.34407, 17.34406, 17.34406, 17.34406, 
    17.34406, 17.34406, 17.34407, 17.34407, 17.34407, 17.34408, 17.34408, 
    17.34408, 17.34407, 17.34406, 17.34406, 17.34405, 17.34405, 17.34403, 
    17.34404, 17.34403, 17.34404, 17.34402, 17.34406, 17.34404, 17.34407, 
    17.34407, 17.34406, 17.34405, 17.34406, 17.34405, 17.34407, 17.34408, 
    17.34408, 17.34408, 17.34408, 17.34408, 17.34407, 17.34408, 17.34406, 
    17.34407, 17.34405, 17.34405, 17.34403, 17.34402, 17.34401, 17.344, 
    17.344, 17.344 ;

 TOTSOMC_1m =
  17.34412, 17.34411, 17.34411, 17.3441, 17.34411, 17.3441, 17.34412, 
    17.34411, 17.34411, 17.34412, 17.34409, 17.3441, 17.34407, 17.34408, 
    17.34406, 17.34407, 17.34406, 17.34406, 17.34405, 17.34405, 17.34404, 
    17.34405, 17.34403, 17.34404, 17.34404, 17.34405, 17.3441, 17.34409, 
    17.3441, 17.3441, 17.3441, 17.34411, 17.34411, 17.34412, 17.34412, 
    17.34411, 17.3441, 17.3441, 17.34409, 17.34409, 17.34408, 17.34408, 
    17.34406, 17.34407, 17.34405, 17.34406, 17.34405, 17.34405, 17.34405, 
    17.34406, 17.34405, 17.34406, 17.34408, 17.34408, 17.3441, 17.34411, 
    17.34412, 17.34412, 17.34412, 17.34412, 17.34411, 17.3441, 17.3441, 
    17.3441, 17.34409, 17.34408, 17.34407, 17.34406, 17.34406, 17.34406, 
    17.34406, 17.34405, 17.34405, 17.34405, 17.34406, 17.34405, 17.34406, 
    17.34406, 17.34409, 17.3441, 17.34411, 17.34411, 17.34412, 17.34411, 
    17.34412, 17.34411, 17.34411, 17.34411, 17.3441, 17.3441, 17.34407, 
    17.34409, 17.34406, 17.34406, 17.34405, 17.34406, 17.34405, 17.34406, 
    17.34405, 17.34404, 17.34405, 17.34404, 17.34406, 17.34405, 17.34411, 
    17.34411, 17.34411, 17.34411, 17.34411, 17.34412, 17.34411, 17.34411, 
    17.34411, 17.3441, 17.3441, 17.34409, 17.34408, 17.34407, 17.34406, 
    17.34406, 17.34406, 17.34406, 17.34406, 17.34406, 17.34404, 17.34405, 
    17.34404, 17.34404, 17.34405, 17.34404, 17.34411, 17.34411, 17.34412, 
    17.34411, 17.34412, 17.34412, 17.34411, 17.3441, 17.3441, 17.3441, 
    17.34409, 17.34408, 17.34407, 17.34406, 17.34406, 17.34406, 17.34406, 
    17.34405, 17.34406, 17.34405, 17.34405, 17.34405, 17.34404, 17.34404, 
    17.34404, 17.34404, 17.34411, 17.34411, 17.34411, 17.3441, 17.34411, 
    17.3441, 17.34409, 17.34408, 17.34408, 17.34407, 17.34408, 17.34408, 
    17.34407, 17.34408, 17.34406, 17.34408, 17.34405, 17.34407, 17.34405, 
    17.34406, 17.34405, 17.34405, 17.34404, 17.34403, 17.34404, 17.34403, 
    17.3441, 17.3441, 17.3441, 17.34409, 17.34409, 17.34408, 17.34407, 
    17.34407, 17.34407, 17.34406, 17.34408, 17.34407, 17.34409, 17.34409, 
    17.34409, 17.3441, 17.34407, 17.34409, 17.34406, 17.34407, 17.34405, 
    17.34406, 17.34404, 17.34403, 17.34402, 17.34401, 17.3441, 17.3441, 
    17.34409, 17.34409, 17.34408, 17.34407, 17.34407, 17.34407, 17.34406, 
    17.34406, 17.34407, 17.34406, 17.34409, 17.34407, 17.3441, 17.34409, 
    17.34409, 17.34409, 17.34408, 17.34407, 17.34406, 17.34407, 17.34403, 
    17.34405, 17.344, 17.34402, 17.3441, 17.3441, 17.34408, 17.34409, 
    17.34407, 17.34406, 17.34406, 17.34406, 17.34406, 17.34405, 17.34406, 
    17.34405, 17.34407, 17.34406, 17.34408, 17.34408, 17.34408, 17.34408, 
    17.34407, 17.34407, 17.34407, 17.34406, 17.34406, 17.34407, 17.34403, 
    17.34405, 17.34409, 17.34408, 17.34408, 17.34408, 17.34406, 17.34407, 
    17.34405, 17.34406, 17.34405, 17.34405, 17.34405, 17.34406, 17.34406, 
    17.34407, 17.34408, 17.34408, 17.34408, 17.34408, 17.34406, 17.34406, 
    17.34406, 17.34405, 17.34407, 17.34406, 17.34406, 17.34406, 17.34407, 
    17.34406, 17.34408, 17.34408, 17.34407, 17.34406, 17.34406, 17.34406, 
    17.34406, 17.34406, 17.34407, 17.34407, 17.34407, 17.34408, 17.34408, 
    17.34408, 17.34407, 17.34406, 17.34406, 17.34405, 17.34405, 17.34403, 
    17.34404, 17.34403, 17.34404, 17.34402, 17.34406, 17.34404, 17.34407, 
    17.34407, 17.34406, 17.34405, 17.34406, 17.34405, 17.34407, 17.34408, 
    17.34408, 17.34408, 17.34408, 17.34408, 17.34407, 17.34408, 17.34406, 
    17.34407, 17.34405, 17.34405, 17.34403, 17.34402, 17.34401, 17.344, 
    17.344, 17.344 ;

 TOTSOMN =
  1.773689, 1.773688, 1.773688, 1.773687, 1.773688, 1.773687, 1.773689, 
    1.773688, 1.773689, 1.773689, 1.773685, 1.773687, 1.773683, 1.773684, 
    1.773681, 1.773683, 1.77368, 1.773681, 1.773679, 1.773679, 1.773677, 
    1.773679, 1.773676, 1.773678, 1.773678, 1.773679, 1.773687, 1.773685, 
    1.773687, 1.773686, 1.773687, 1.773688, 1.773688, 1.773689, 1.773689, 
    1.773688, 1.773686, 1.773687, 1.773685, 1.773685, 1.773683, 1.773684, 
    1.773681, 1.773682, 1.773679, 1.77368, 1.773679, 1.77368, 1.773679, 
    1.77368, 1.77368, 1.773681, 1.773684, 1.773683, 1.773686, 1.773688, 
    1.773689, 1.77369, 1.77369, 1.773689, 1.773688, 1.773687, 1.773686, 
    1.773686, 1.773685, 1.773684, 1.773683, 1.773681, 1.773681, 1.773681, 
    1.77368, 1.773679, 1.773679, 1.773679, 1.773681, 1.773679, 1.773682, 
    1.773681, 1.773685, 1.773687, 1.773687, 1.773688, 1.77369, 1.773689, 
    1.773689, 1.773688, 1.773687, 1.773688, 1.773686, 1.773687, 1.773683, 
    1.773684, 1.77368, 1.773681, 1.77368, 1.773681, 1.773679, 1.77368, 
    1.773679, 1.773678, 1.773679, 1.773678, 1.773681, 1.773679, 1.773688, 
    1.773688, 1.773687, 1.773688, 1.773688, 1.773689, 1.773689, 1.773688, 
    1.773687, 1.773687, 1.773686, 1.773685, 1.773684, 1.773682, 1.773681, 
    1.77368, 1.773681, 1.77368, 1.773681, 1.773681, 1.773679, 1.77368, 
    1.773678, 1.773678, 1.773679, 1.773678, 1.773688, 1.773688, 1.773689, 
    1.773688, 1.77369, 1.773689, 1.773688, 1.773687, 1.773686, 1.773686, 
    1.773685, 1.773684, 1.773683, 1.773681, 1.77368, 1.77368, 1.77368, 
    1.77368, 1.773681, 1.77368, 1.77368, 1.77368, 1.773678, 1.773679, 
    1.773678, 1.773678, 1.773688, 1.773687, 1.773688, 1.773687, 1.773687, 
    1.773686, 1.773685, 1.773683, 1.773684, 1.773683, 1.773684, 1.773684, 
    1.773683, 1.773684, 1.773681, 1.773683, 1.77368, 1.773682, 1.77368, 
    1.77368, 1.773679, 1.773679, 1.773678, 1.773677, 1.773677, 1.773677, 
    1.773687, 1.773686, 1.773686, 1.773685, 1.773685, 1.773684, 1.773682, 
    1.773683, 1.773682, 1.773682, 1.773683, 1.773682, 1.773686, 1.773685, 
    1.773685, 1.773687, 1.773683, 1.773685, 1.773681, 1.773682, 1.773679, 
    1.773681, 1.773678, 1.773676, 1.773675, 1.773674, 1.773686, 1.773686, 
    1.773685, 1.773684, 1.773683, 1.773682, 1.773682, 1.773682, 1.773681, 
    1.773681, 1.773682, 1.77368, 1.773685, 1.773683, 1.773686, 1.773685, 
    1.773684, 1.773685, 1.773683, 1.773683, 1.773681, 1.773682, 1.773677, 
    1.773679, 1.773673, 1.773674, 1.773686, 1.773686, 1.773684, 1.773685, 
    1.773682, 1.773681, 1.773681, 1.77368, 1.77368, 1.77368, 1.77368, 
    1.77368, 1.773682, 1.773681, 1.773684, 1.773683, 1.773684, 1.773684, 
    1.773683, 1.773682, 1.773682, 1.773681, 1.77368, 1.773682, 1.773676, 
    1.77368, 1.773685, 1.773684, 1.773684, 1.773684, 1.773681, 1.773682, 
    1.77368, 1.77368, 1.773679, 1.77368, 1.77368, 1.773681, 1.773681, 
    1.773682, 1.773683, 1.773684, 1.773684, 1.773683, 1.773682, 1.77368, 
    1.77368, 1.773679, 1.773682, 1.773681, 1.773682, 1.77368, 1.773683, 
    1.773681, 1.773684, 1.773683, 1.773682, 1.773681, 1.773681, 1.77368, 
    1.77368, 1.773682, 1.773682, 1.773682, 1.773683, 1.773683, 1.773684, 
    1.773683, 1.773683, 1.773682, 1.77368, 1.773679, 1.773679, 1.773677, 
    1.773678, 1.773676, 1.773678, 1.773675, 1.773681, 1.773678, 1.773682, 
    1.773682, 1.773681, 1.773679, 1.77368, 1.773679, 1.773682, 1.773683, 
    1.773684, 1.773684, 1.773683, 1.773684, 1.773683, 1.773683, 1.773682, 
    1.773682, 1.77368, 1.773679, 1.773677, 1.773675, 1.773674, 1.773673, 
    1.773673, 1.773673 ;

 TOTSOMN_1m =
  1.773689, 1.773688, 1.773688, 1.773687, 1.773688, 1.773687, 1.773689, 
    1.773688, 1.773689, 1.773689, 1.773685, 1.773687, 1.773683, 1.773684, 
    1.773681, 1.773683, 1.77368, 1.773681, 1.773679, 1.773679, 1.773677, 
    1.773679, 1.773676, 1.773678, 1.773678, 1.773679, 1.773687, 1.773685, 
    1.773687, 1.773686, 1.773687, 1.773688, 1.773688, 1.773689, 1.773689, 
    1.773688, 1.773686, 1.773687, 1.773685, 1.773685, 1.773683, 1.773684, 
    1.773681, 1.773682, 1.773679, 1.77368, 1.773679, 1.77368, 1.773679, 
    1.77368, 1.77368, 1.773681, 1.773684, 1.773683, 1.773686, 1.773688, 
    1.773689, 1.77369, 1.77369, 1.773689, 1.773688, 1.773687, 1.773686, 
    1.773686, 1.773685, 1.773684, 1.773683, 1.773681, 1.773681, 1.773681, 
    1.77368, 1.773679, 1.773679, 1.773679, 1.773681, 1.773679, 1.773682, 
    1.773681, 1.773685, 1.773687, 1.773687, 1.773688, 1.77369, 1.773689, 
    1.773689, 1.773688, 1.773687, 1.773688, 1.773686, 1.773687, 1.773683, 
    1.773684, 1.77368, 1.773681, 1.77368, 1.773681, 1.773679, 1.77368, 
    1.773679, 1.773678, 1.773679, 1.773678, 1.773681, 1.773679, 1.773688, 
    1.773688, 1.773687, 1.773688, 1.773688, 1.773689, 1.773689, 1.773688, 
    1.773687, 1.773687, 1.773686, 1.773685, 1.773684, 1.773682, 1.773681, 
    1.77368, 1.773681, 1.77368, 1.773681, 1.773681, 1.773679, 1.77368, 
    1.773678, 1.773678, 1.773679, 1.773678, 1.773688, 1.773688, 1.773689, 
    1.773688, 1.77369, 1.773689, 1.773688, 1.773687, 1.773686, 1.773686, 
    1.773685, 1.773684, 1.773683, 1.773681, 1.77368, 1.77368, 1.77368, 
    1.77368, 1.773681, 1.77368, 1.77368, 1.77368, 1.773678, 1.773679, 
    1.773678, 1.773678, 1.773688, 1.773687, 1.773688, 1.773687, 1.773687, 
    1.773686, 1.773685, 1.773683, 1.773684, 1.773683, 1.773684, 1.773684, 
    1.773683, 1.773684, 1.773681, 1.773683, 1.77368, 1.773682, 1.77368, 
    1.77368, 1.773679, 1.773679, 1.773678, 1.773677, 1.773677, 1.773677, 
    1.773687, 1.773686, 1.773686, 1.773685, 1.773685, 1.773684, 1.773682, 
    1.773683, 1.773682, 1.773682, 1.773683, 1.773682, 1.773686, 1.773685, 
    1.773685, 1.773687, 1.773683, 1.773685, 1.773681, 1.773682, 1.773679, 
    1.773681, 1.773678, 1.773676, 1.773675, 1.773674, 1.773686, 1.773686, 
    1.773685, 1.773684, 1.773683, 1.773682, 1.773682, 1.773682, 1.773681, 
    1.773681, 1.773682, 1.77368, 1.773685, 1.773683, 1.773686, 1.773685, 
    1.773684, 1.773685, 1.773683, 1.773683, 1.773681, 1.773682, 1.773677, 
    1.773679, 1.773673, 1.773674, 1.773686, 1.773686, 1.773684, 1.773685, 
    1.773682, 1.773681, 1.773681, 1.77368, 1.77368, 1.77368, 1.77368, 
    1.77368, 1.773682, 1.773681, 1.773684, 1.773683, 1.773684, 1.773684, 
    1.773683, 1.773682, 1.773682, 1.773681, 1.77368, 1.773682, 1.773676, 
    1.77368, 1.773685, 1.773684, 1.773684, 1.773684, 1.773681, 1.773682, 
    1.77368, 1.77368, 1.773679, 1.77368, 1.77368, 1.773681, 1.773681, 
    1.773682, 1.773683, 1.773684, 1.773684, 1.773683, 1.773682, 1.77368, 
    1.77368, 1.773679, 1.773682, 1.773681, 1.773682, 1.77368, 1.773683, 
    1.773681, 1.773684, 1.773683, 1.773682, 1.773681, 1.773681, 1.77368, 
    1.77368, 1.773682, 1.773682, 1.773682, 1.773683, 1.773683, 1.773684, 
    1.773683, 1.773683, 1.773682, 1.77368, 1.773679, 1.773679, 1.773677, 
    1.773678, 1.773676, 1.773678, 1.773675, 1.773681, 1.773678, 1.773682, 
    1.773682, 1.773681, 1.773679, 1.77368, 1.773679, 1.773682, 1.773683, 
    1.773684, 1.773684, 1.773683, 1.773684, 1.773683, 1.773683, 1.773682, 
    1.773682, 1.77368, 1.773679, 1.773677, 1.773675, 1.773674, 1.773673, 
    1.773673, 1.773673 ;

 TOTVEGC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTVEGN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TREFMNAV =
  249.9921, 249.9923, 249.9923, 249.9925, 249.9924, 249.9925, 249.9921, 
    249.9923, 249.9922, 249.9921, 249.9928, 249.9925, 249.9932, 249.993, 
    249.9936, 249.9932, 249.9937, 249.9936, 249.9939, 249.9938, 249.9941, 
    249.9939, 249.9943, 249.9941, 249.9941, 249.9939, 249.9926, 249.9928, 
    249.9925, 249.9926, 249.9926, 249.9924, 249.9923, 249.9921, 249.9921, 
    249.9922, 249.9926, 249.9925, 249.9928, 249.9928, 249.9931, 249.9929, 
    249.9935, 249.9933, 249.9938, 249.9937, 249.9938, 249.9937, 249.9938, 
    249.9936, 249.9937, 249.9935, 249.993, 249.9931, 249.9926, 249.9923, 
    249.9921, 249.992, 249.992, 249.9921, 249.9922, 249.9924, 249.9926, 
    249.9927, 249.9928, 249.993, 249.9932, 249.9935, 249.9935, 249.9935, 
    249.9937, 249.9938, 249.9938, 249.9939, 249.9935, 249.9937, 249.9934, 
    249.9935, 249.9928, 249.9925, 249.9924, 249.9923, 249.992, 249.9922, 
    249.9921, 249.9923, 249.9924, 249.9924, 249.9927, 249.9926, 249.9932, 
    249.9929, 249.9936, 249.9935, 249.9937, 249.9936, 249.9938, 249.9936, 
    249.9939, 249.9939, 249.9939, 249.9941, 249.9936, 249.9938, 249.9924, 
    249.9924, 249.9924, 249.9922, 249.9922, 249.9921, 249.9922, 249.9923, 
    249.9924, 249.9925, 249.9926, 249.9928, 249.993, 249.9933, 249.9935, 
    249.9936, 249.9935, 249.9936, 249.9935, 249.9935, 249.9939, 249.9937, 
    249.994, 249.994, 249.9939, 249.994, 249.9924, 249.9923, 249.9922, 
    249.9923, 249.9921, 249.9922, 249.9922, 249.9926, 249.9926, 249.9927, 
    249.9928, 249.993, 249.9932, 249.9934, 249.9937, 249.9936, 249.9937, 
    249.9937, 249.9936, 249.9937, 249.9937, 249.9937, 249.994, 249.9939, 
    249.994, 249.994, 249.9923, 249.9924, 249.9924, 249.9924, 249.9924, 
    249.9926, 249.9927, 249.9931, 249.9929, 249.9932, 249.993, 249.993, 
    249.9932, 249.993, 249.9934, 249.9931, 249.9937, 249.9934, 249.9937, 
    249.9937, 249.9938, 249.9938, 249.994, 249.9942, 249.9941, 249.9943, 
    249.9925, 249.9926, 249.9926, 249.9927, 249.9928, 249.993, 249.9933, 
    249.9932, 249.9934, 249.9934, 249.9931, 249.9933, 249.9927, 249.9928, 
    249.9928, 249.9925, 249.9932, 249.9929, 249.9935, 249.9933, 249.9938, 
    249.9936, 249.9941, 249.9943, 249.9945, 249.9948, 249.9927, 249.9926, 
    249.9928, 249.9929, 249.9931, 249.9933, 249.9933, 249.9934, 249.9935, 
    249.9936, 249.9934, 249.9936, 249.9928, 249.9932, 249.9926, 249.9928, 
    249.9929, 249.9929, 249.9932, 249.9932, 249.9935, 249.9934, 249.9942, 
    249.9939, 249.9949, 249.9946, 249.9926, 249.9927, 249.993, 249.9929, 
    249.9933, 249.9934, 249.9935, 249.9936, 249.9937, 249.9937, 249.9936, 
    249.9937, 249.9933, 249.9935, 249.993, 249.9931, 249.9931, 249.993, 
    249.9932, 249.9934, 249.9934, 249.9935, 249.9936, 249.9933, 249.9943, 
    249.9937, 249.9928, 249.993, 249.993, 249.9929, 249.9934, 249.9932, 
    249.9937, 249.9936, 249.9938, 249.9937, 249.9937, 249.9935, 249.9935, 
    249.9933, 249.9931, 249.993, 249.993, 249.9931, 249.9934, 249.9937, 
    249.9936, 249.9938, 249.9933, 249.9935, 249.9934, 249.9936, 249.9932, 
    249.9935, 249.9931, 249.9931, 249.9932, 249.9935, 249.9936, 249.9936, 
    249.9936, 249.9934, 249.9934, 249.9932, 249.9932, 249.9931, 249.993, 
    249.9931, 249.9932, 249.9934, 249.9936, 249.9938, 249.9939, 249.9942, 
    249.9939, 249.9943, 249.994, 249.9945, 249.9936, 249.994, 249.9933, 
    249.9933, 249.9935, 249.9938, 249.9936, 249.9938, 249.9934, 249.9931, 
    249.9931, 249.993, 249.9931, 249.9931, 249.9932, 249.9931, 249.9934, 
    249.9933, 249.9937, 249.9938, 249.9943, 249.9945, 249.9948, 249.9949, 
    249.9949, 249.995 ;

 TREFMNAV_R =
  249.9921, 249.9923, 249.9923, 249.9925, 249.9924, 249.9925, 249.9921, 
    249.9923, 249.9922, 249.9921, 249.9928, 249.9925, 249.9932, 249.993, 
    249.9936, 249.9932, 249.9937, 249.9936, 249.9939, 249.9938, 249.9941, 
    249.9939, 249.9943, 249.9941, 249.9941, 249.9939, 249.9926, 249.9928, 
    249.9925, 249.9926, 249.9926, 249.9924, 249.9923, 249.9921, 249.9921, 
    249.9922, 249.9926, 249.9925, 249.9928, 249.9928, 249.9931, 249.9929, 
    249.9935, 249.9933, 249.9938, 249.9937, 249.9938, 249.9937, 249.9938, 
    249.9936, 249.9937, 249.9935, 249.993, 249.9931, 249.9926, 249.9923, 
    249.9921, 249.992, 249.992, 249.9921, 249.9922, 249.9924, 249.9926, 
    249.9927, 249.9928, 249.993, 249.9932, 249.9935, 249.9935, 249.9935, 
    249.9937, 249.9938, 249.9938, 249.9939, 249.9935, 249.9937, 249.9934, 
    249.9935, 249.9928, 249.9925, 249.9924, 249.9923, 249.992, 249.9922, 
    249.9921, 249.9923, 249.9924, 249.9924, 249.9927, 249.9926, 249.9932, 
    249.9929, 249.9936, 249.9935, 249.9937, 249.9936, 249.9938, 249.9936, 
    249.9939, 249.9939, 249.9939, 249.9941, 249.9936, 249.9938, 249.9924, 
    249.9924, 249.9924, 249.9922, 249.9922, 249.9921, 249.9922, 249.9923, 
    249.9924, 249.9925, 249.9926, 249.9928, 249.993, 249.9933, 249.9935, 
    249.9936, 249.9935, 249.9936, 249.9935, 249.9935, 249.9939, 249.9937, 
    249.994, 249.994, 249.9939, 249.994, 249.9924, 249.9923, 249.9922, 
    249.9923, 249.9921, 249.9922, 249.9922, 249.9926, 249.9926, 249.9927, 
    249.9928, 249.993, 249.9932, 249.9934, 249.9937, 249.9936, 249.9937, 
    249.9937, 249.9936, 249.9937, 249.9937, 249.9937, 249.994, 249.9939, 
    249.994, 249.994, 249.9923, 249.9924, 249.9924, 249.9924, 249.9924, 
    249.9926, 249.9927, 249.9931, 249.9929, 249.9932, 249.993, 249.993, 
    249.9932, 249.993, 249.9934, 249.9931, 249.9937, 249.9934, 249.9937, 
    249.9937, 249.9938, 249.9938, 249.994, 249.9942, 249.9941, 249.9943, 
    249.9925, 249.9926, 249.9926, 249.9927, 249.9928, 249.993, 249.9933, 
    249.9932, 249.9934, 249.9934, 249.9931, 249.9933, 249.9927, 249.9928, 
    249.9928, 249.9925, 249.9932, 249.9929, 249.9935, 249.9933, 249.9938, 
    249.9936, 249.9941, 249.9943, 249.9945, 249.9948, 249.9927, 249.9926, 
    249.9928, 249.9929, 249.9931, 249.9933, 249.9933, 249.9934, 249.9935, 
    249.9936, 249.9934, 249.9936, 249.9928, 249.9932, 249.9926, 249.9928, 
    249.9929, 249.9929, 249.9932, 249.9932, 249.9935, 249.9934, 249.9942, 
    249.9939, 249.9949, 249.9946, 249.9926, 249.9927, 249.993, 249.9929, 
    249.9933, 249.9934, 249.9935, 249.9936, 249.9937, 249.9937, 249.9936, 
    249.9937, 249.9933, 249.9935, 249.993, 249.9931, 249.9931, 249.993, 
    249.9932, 249.9934, 249.9934, 249.9935, 249.9936, 249.9933, 249.9943, 
    249.9937, 249.9928, 249.993, 249.993, 249.9929, 249.9934, 249.9932, 
    249.9937, 249.9936, 249.9938, 249.9937, 249.9937, 249.9935, 249.9935, 
    249.9933, 249.9931, 249.993, 249.993, 249.9931, 249.9934, 249.9937, 
    249.9936, 249.9938, 249.9933, 249.9935, 249.9934, 249.9936, 249.9932, 
    249.9935, 249.9931, 249.9931, 249.9932, 249.9935, 249.9936, 249.9936, 
    249.9936, 249.9934, 249.9934, 249.9932, 249.9932, 249.9931, 249.993, 
    249.9931, 249.9932, 249.9934, 249.9936, 249.9938, 249.9939, 249.9942, 
    249.9939, 249.9943, 249.994, 249.9945, 249.9936, 249.994, 249.9933, 
    249.9933, 249.9935, 249.9938, 249.9936, 249.9938, 249.9934, 249.9931, 
    249.9931, 249.993, 249.9931, 249.9931, 249.9932, 249.9931, 249.9934, 
    249.9933, 249.9937, 249.9938, 249.9943, 249.9945, 249.9948, 249.9949, 
    249.9949, 249.995 ;

 TREFMNAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TREFMXAV =
  258.6147, 258.615, 258.6149, 258.6152, 258.615, 258.6152, 258.6147, 
    258.615, 258.6148, 258.6147, 258.6156, 258.6152, 258.6161, 258.6158, 
    258.6166, 258.6161, 258.6167, 258.6166, 258.617, 258.6169, 258.6173, 
    258.617, 258.6176, 258.6172, 258.6173, 258.617, 258.6153, 258.6156, 
    258.6153, 258.6153, 258.6153, 258.615, 258.6149, 258.6146, 258.6147, 
    258.6149, 258.6153, 258.6152, 258.6155, 258.6155, 258.616, 258.6158, 
    258.6165, 258.6163, 258.6169, 258.6167, 258.6169, 258.6168, 258.6169, 
    258.6166, 258.6167, 258.6165, 258.6158, 258.616, 258.6154, 258.615, 
    258.6147, 258.6146, 258.6146, 258.6146, 258.6149, 258.6151, 258.6153, 
    258.6154, 258.6155, 258.6159, 258.6161, 258.6165, 258.6165, 258.6166, 
    258.6167, 258.6169, 258.6169, 258.617, 258.6166, 258.6168, 258.6164, 
    258.6165, 258.6155, 258.6152, 258.6151, 258.6149, 258.6146, 258.6148, 
    258.6147, 258.615, 258.6151, 258.615, 258.6154, 258.6153, 258.6161, 
    258.6157, 258.6167, 258.6165, 258.6167, 258.6166, 258.6169, 258.6166, 
    258.617, 258.6171, 258.617, 258.6172, 258.6166, 258.6169, 258.615, 
    258.615, 258.6151, 258.6148, 258.6148, 258.6146, 258.6148, 258.6149, 
    258.6151, 258.6152, 258.6153, 258.6155, 258.6158, 258.6162, 258.6165, 
    258.6167, 258.6165, 258.6166, 258.6165, 258.6165, 258.6171, 258.6167, 
    258.6172, 258.6172, 258.617, 258.6172, 258.615, 258.615, 258.6147, 
    258.6149, 258.6146, 258.6148, 258.6149, 258.6153, 258.6154, 258.6154, 
    258.6156, 258.6158, 258.6161, 258.6164, 258.6167, 258.6167, 258.6167, 
    258.6168, 258.6166, 258.6168, 258.6168, 258.6167, 258.6172, 258.6171, 
    258.6172, 258.6171, 258.615, 258.6151, 258.615, 258.6151, 258.6151, 
    258.6154, 258.6155, 258.616, 258.6158, 258.6161, 258.6158, 258.6158, 
    258.6161, 258.6158, 258.6164, 258.616, 258.6168, 258.6163, 258.6168, 
    258.6167, 258.6169, 258.6169, 258.6171, 258.6174, 258.6173, 258.6175, 
    258.6152, 258.6154, 258.6154, 258.6155, 258.6156, 258.6158, 258.6162, 
    258.6161, 258.6163, 258.6164, 258.616, 258.6162, 258.6155, 258.6156, 
    258.6155, 258.6153, 258.6161, 258.6157, 258.6165, 258.6162, 258.6169, 
    258.6166, 258.6173, 258.6176, 258.6178, 258.6181, 258.6154, 258.6154, 
    258.6155, 258.6158, 258.616, 258.6162, 258.6163, 258.6163, 258.6165, 
    258.6166, 258.6164, 258.6166, 258.6156, 258.6161, 258.6153, 258.6156, 
    258.6158, 258.6157, 258.6161, 258.6161, 258.6165, 258.6163, 258.6175, 
    258.617, 258.6184, 258.618, 258.6153, 258.6154, 258.6159, 258.6157, 
    258.6163, 258.6164, 258.6165, 258.6167, 258.6167, 258.6168, 258.6166, 
    258.6168, 258.6162, 258.6165, 258.6158, 258.616, 258.6159, 258.6158, 
    258.6161, 258.6164, 258.6164, 258.6165, 258.6167, 258.6163, 258.6175, 
    258.6167, 258.6156, 258.6158, 258.6159, 258.6158, 258.6164, 258.6162, 
    258.6168, 258.6166, 258.6169, 258.6168, 258.6168, 258.6166, 258.6165, 
    258.6162, 258.616, 258.6158, 258.6158, 258.616, 258.6164, 258.6167, 
    258.6166, 258.6169, 258.6162, 258.6165, 258.6164, 258.6167, 258.6161, 
    258.6166, 258.6159, 258.616, 258.6162, 258.6165, 258.6166, 258.6167, 
    258.6166, 258.6164, 258.6163, 258.6162, 258.6161, 258.616, 258.6159, 
    258.616, 258.6161, 258.6164, 258.6167, 258.6169, 258.617, 258.6174, 
    258.6171, 258.6175, 258.6171, 258.6178, 258.6166, 258.6171, 258.6162, 
    258.6163, 258.6165, 258.6169, 258.6167, 258.6169, 258.6163, 258.616, 
    258.6159, 258.6158, 258.616, 258.6159, 258.6161, 258.616, 258.6164, 
    258.6162, 258.6167, 258.6169, 258.6175, 258.6178, 258.6182, 258.6183, 
    258.6184, 258.6184 ;

 TREFMXAV_R =
  258.6147, 258.615, 258.6149, 258.6152, 258.615, 258.6152, 258.6147, 
    258.615, 258.6148, 258.6147, 258.6156, 258.6152, 258.6161, 258.6158, 
    258.6166, 258.6161, 258.6167, 258.6166, 258.617, 258.6169, 258.6173, 
    258.617, 258.6176, 258.6172, 258.6173, 258.617, 258.6153, 258.6156, 
    258.6153, 258.6153, 258.6153, 258.615, 258.6149, 258.6146, 258.6147, 
    258.6149, 258.6153, 258.6152, 258.6155, 258.6155, 258.616, 258.6158, 
    258.6165, 258.6163, 258.6169, 258.6167, 258.6169, 258.6168, 258.6169, 
    258.6166, 258.6167, 258.6165, 258.6158, 258.616, 258.6154, 258.615, 
    258.6147, 258.6146, 258.6146, 258.6146, 258.6149, 258.6151, 258.6153, 
    258.6154, 258.6155, 258.6159, 258.6161, 258.6165, 258.6165, 258.6166, 
    258.6167, 258.6169, 258.6169, 258.617, 258.6166, 258.6168, 258.6164, 
    258.6165, 258.6155, 258.6152, 258.6151, 258.6149, 258.6146, 258.6148, 
    258.6147, 258.615, 258.6151, 258.615, 258.6154, 258.6153, 258.6161, 
    258.6157, 258.6167, 258.6165, 258.6167, 258.6166, 258.6169, 258.6166, 
    258.617, 258.6171, 258.617, 258.6172, 258.6166, 258.6169, 258.615, 
    258.615, 258.6151, 258.6148, 258.6148, 258.6146, 258.6148, 258.6149, 
    258.6151, 258.6152, 258.6153, 258.6155, 258.6158, 258.6162, 258.6165, 
    258.6167, 258.6165, 258.6166, 258.6165, 258.6165, 258.6171, 258.6167, 
    258.6172, 258.6172, 258.617, 258.6172, 258.615, 258.615, 258.6147, 
    258.6149, 258.6146, 258.6148, 258.6149, 258.6153, 258.6154, 258.6154, 
    258.6156, 258.6158, 258.6161, 258.6164, 258.6167, 258.6167, 258.6167, 
    258.6168, 258.6166, 258.6168, 258.6168, 258.6167, 258.6172, 258.6171, 
    258.6172, 258.6171, 258.615, 258.6151, 258.615, 258.6151, 258.6151, 
    258.6154, 258.6155, 258.616, 258.6158, 258.6161, 258.6158, 258.6158, 
    258.6161, 258.6158, 258.6164, 258.616, 258.6168, 258.6163, 258.6168, 
    258.6167, 258.6169, 258.6169, 258.6171, 258.6174, 258.6173, 258.6175, 
    258.6152, 258.6154, 258.6154, 258.6155, 258.6156, 258.6158, 258.6162, 
    258.6161, 258.6163, 258.6164, 258.616, 258.6162, 258.6155, 258.6156, 
    258.6155, 258.6153, 258.6161, 258.6157, 258.6165, 258.6162, 258.6169, 
    258.6166, 258.6173, 258.6176, 258.6178, 258.6181, 258.6154, 258.6154, 
    258.6155, 258.6158, 258.616, 258.6162, 258.6163, 258.6163, 258.6165, 
    258.6166, 258.6164, 258.6166, 258.6156, 258.6161, 258.6153, 258.6156, 
    258.6158, 258.6157, 258.6161, 258.6161, 258.6165, 258.6163, 258.6175, 
    258.617, 258.6184, 258.618, 258.6153, 258.6154, 258.6159, 258.6157, 
    258.6163, 258.6164, 258.6165, 258.6167, 258.6167, 258.6168, 258.6166, 
    258.6168, 258.6162, 258.6165, 258.6158, 258.616, 258.6159, 258.6158, 
    258.6161, 258.6164, 258.6164, 258.6165, 258.6167, 258.6163, 258.6175, 
    258.6167, 258.6156, 258.6158, 258.6159, 258.6158, 258.6164, 258.6162, 
    258.6168, 258.6166, 258.6169, 258.6168, 258.6168, 258.6166, 258.6165, 
    258.6162, 258.616, 258.6158, 258.6158, 258.616, 258.6164, 258.6167, 
    258.6166, 258.6169, 258.6162, 258.6165, 258.6164, 258.6167, 258.6161, 
    258.6166, 258.6159, 258.616, 258.6162, 258.6165, 258.6166, 258.6167, 
    258.6166, 258.6164, 258.6163, 258.6162, 258.6161, 258.616, 258.6159, 
    258.616, 258.6161, 258.6164, 258.6167, 258.6169, 258.617, 258.6174, 
    258.6171, 258.6175, 258.6171, 258.6178, 258.6166, 258.6171, 258.6162, 
    258.6163, 258.6165, 258.6169, 258.6167, 258.6169, 258.6163, 258.616, 
    258.6159, 258.6158, 258.616, 258.6159, 258.6161, 258.616, 258.6164, 
    258.6162, 258.6167, 258.6169, 258.6175, 258.6178, 258.6182, 258.6183, 
    258.6184, 258.6184 ;

 TREFMXAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSA =
  253.98, 253.9802, 253.9801, 253.9803, 253.9802, 253.9803, 253.98, 253.9802, 
    253.9801, 253.98, 253.9805, 253.9803, 253.9808, 253.9806, 253.981, 
    253.9807, 253.981, 253.981, 253.9812, 253.9811, 253.9814, 253.9812, 
    253.9815, 253.9813, 253.9813, 253.9812, 253.9803, 253.9805, 253.9803, 
    253.9803, 253.9803, 253.9802, 253.9801, 253.98, 253.98, 253.9801, 
    253.9803, 253.9803, 253.9805, 253.9805, 253.9807, 253.9806, 253.9809, 
    253.9808, 253.9811, 253.981, 253.9811, 253.9811, 253.9811, 253.981, 
    253.9811, 253.981, 253.9806, 253.9807, 253.9804, 253.9802, 253.98, 
    253.9799, 253.98, 253.98, 253.9801, 253.9802, 253.9803, 253.9804, 
    253.9805, 253.9806, 253.9807, 253.9809, 253.9809, 253.981, 253.981, 
    253.9812, 253.9811, 253.9812, 253.981, 253.9811, 253.9809, 253.9809, 
    253.9805, 253.9803, 253.9802, 253.9801, 253.98, 253.9801, 253.98, 
    253.9801, 253.9802, 253.9802, 253.9804, 253.9803, 253.9807, 253.9805, 
    253.981, 253.9809, 253.9811, 253.981, 253.9811, 253.981, 253.9812, 
    253.9812, 253.9812, 253.9813, 253.981, 253.9811, 253.9802, 253.9802, 
    253.9802, 253.9801, 253.9801, 253.98, 253.9801, 253.9801, 253.9802, 
    253.9803, 253.9803, 253.9805, 253.9806, 253.9808, 253.9809, 253.981, 
    253.981, 253.981, 253.981, 253.9809, 253.9812, 253.981, 253.9813, 
    253.9813, 253.9812, 253.9813, 253.9802, 253.9802, 253.98, 253.9801, 
    253.98, 253.9801, 253.9801, 253.9803, 253.9803, 253.9804, 253.9805, 
    253.9806, 253.9807, 253.9809, 253.981, 253.981, 253.981, 253.9811, 
    253.981, 253.9811, 253.9811, 253.9811, 253.9813, 253.9812, 253.9813, 
    253.9812, 253.9802, 253.9802, 253.9802, 253.9802, 253.9802, 253.9804, 
    253.9804, 253.9807, 253.9806, 253.9807, 253.9806, 253.9806, 253.9807, 
    253.9806, 253.9809, 253.9807, 253.9811, 253.9809, 253.9811, 253.981, 
    253.9811, 253.9812, 253.9812, 253.9814, 253.9813, 253.9815, 253.9803, 
    253.9804, 253.9804, 253.9804, 253.9805, 253.9806, 253.9808, 253.9807, 
    253.9809, 253.9809, 253.9807, 253.9808, 253.9804, 253.9805, 253.9804, 
    253.9803, 253.9807, 253.9805, 253.9809, 253.9808, 253.9812, 253.981, 
    253.9813, 253.9815, 253.9816, 253.9818, 253.9804, 253.9804, 253.9804, 
    253.9806, 253.9807, 253.9808, 253.9808, 253.9809, 253.9809, 253.981, 
    253.9809, 253.981, 253.9805, 253.9808, 253.9803, 253.9805, 253.9805, 
    253.9805, 253.9807, 253.9808, 253.981, 253.9809, 253.9814, 253.9812, 
    253.9819, 253.9817, 253.9803, 253.9804, 253.9806, 253.9805, 253.9808, 
    253.9809, 253.981, 253.981, 253.981, 253.9811, 253.981, 253.9811, 
    253.9808, 253.9809, 253.9806, 253.9807, 253.9807, 253.9806, 253.9807, 
    253.9809, 253.9809, 253.9809, 253.981, 253.9808, 253.9815, 253.9811, 
    253.9805, 253.9806, 253.9806, 253.9806, 253.9809, 253.9808, 253.9811, 
    253.981, 253.9811, 253.9811, 253.9811, 253.981, 253.9809, 253.9808, 
    253.9807, 253.9806, 253.9806, 253.9807, 253.9809, 253.981, 253.981, 
    253.9811, 253.9808, 253.9809, 253.9809, 253.981, 253.9807, 253.981, 
    253.9807, 253.9807, 253.9808, 253.9809, 253.981, 253.981, 253.981, 
    253.9809, 253.9809, 253.9808, 253.9807, 253.9807, 253.9806, 253.9807, 
    253.9807, 253.9809, 253.981, 253.9812, 253.9812, 253.9814, 253.9812, 
    253.9815, 253.9813, 253.9816, 253.981, 253.9813, 253.9808, 253.9808, 
    253.9809, 253.9811, 253.981, 253.9812, 253.9809, 253.9807, 253.9807, 
    253.9806, 253.9807, 253.9807, 253.9807, 253.9807, 253.9809, 253.9808, 
    253.9811, 253.9812, 253.9814, 253.9816, 253.9818, 253.9819, 253.9819, 
    253.9819 ;

 TSAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 TSA_R =
  253.98, 253.9802, 253.9801, 253.9803, 253.9802, 253.9803, 253.98, 253.9802, 
    253.9801, 253.98, 253.9805, 253.9803, 253.9808, 253.9806, 253.981, 
    253.9807, 253.981, 253.981, 253.9812, 253.9811, 253.9814, 253.9812, 
    253.9815, 253.9813, 253.9813, 253.9812, 253.9803, 253.9805, 253.9803, 
    253.9803, 253.9803, 253.9802, 253.9801, 253.98, 253.98, 253.9801, 
    253.9803, 253.9803, 253.9805, 253.9805, 253.9807, 253.9806, 253.9809, 
    253.9808, 253.9811, 253.981, 253.9811, 253.9811, 253.9811, 253.981, 
    253.9811, 253.981, 253.9806, 253.9807, 253.9804, 253.9802, 253.98, 
    253.9799, 253.98, 253.98, 253.9801, 253.9802, 253.9803, 253.9804, 
    253.9805, 253.9806, 253.9807, 253.9809, 253.9809, 253.981, 253.981, 
    253.9812, 253.9811, 253.9812, 253.981, 253.9811, 253.9809, 253.9809, 
    253.9805, 253.9803, 253.9802, 253.9801, 253.98, 253.9801, 253.98, 
    253.9801, 253.9802, 253.9802, 253.9804, 253.9803, 253.9807, 253.9805, 
    253.981, 253.9809, 253.9811, 253.981, 253.9811, 253.981, 253.9812, 
    253.9812, 253.9812, 253.9813, 253.981, 253.9811, 253.9802, 253.9802, 
    253.9802, 253.9801, 253.9801, 253.98, 253.9801, 253.9801, 253.9802, 
    253.9803, 253.9803, 253.9805, 253.9806, 253.9808, 253.9809, 253.981, 
    253.981, 253.981, 253.981, 253.9809, 253.9812, 253.981, 253.9813, 
    253.9813, 253.9812, 253.9813, 253.9802, 253.9802, 253.98, 253.9801, 
    253.98, 253.9801, 253.9801, 253.9803, 253.9803, 253.9804, 253.9805, 
    253.9806, 253.9807, 253.9809, 253.981, 253.981, 253.981, 253.9811, 
    253.981, 253.9811, 253.9811, 253.9811, 253.9813, 253.9812, 253.9813, 
    253.9812, 253.9802, 253.9802, 253.9802, 253.9802, 253.9802, 253.9804, 
    253.9804, 253.9807, 253.9806, 253.9807, 253.9806, 253.9806, 253.9807, 
    253.9806, 253.9809, 253.9807, 253.9811, 253.9809, 253.9811, 253.981, 
    253.9811, 253.9812, 253.9812, 253.9814, 253.9813, 253.9815, 253.9803, 
    253.9804, 253.9804, 253.9804, 253.9805, 253.9806, 253.9808, 253.9807, 
    253.9809, 253.9809, 253.9807, 253.9808, 253.9804, 253.9805, 253.9804, 
    253.9803, 253.9807, 253.9805, 253.9809, 253.9808, 253.9812, 253.981, 
    253.9813, 253.9815, 253.9816, 253.9818, 253.9804, 253.9804, 253.9804, 
    253.9806, 253.9807, 253.9808, 253.9808, 253.9809, 253.9809, 253.981, 
    253.9809, 253.981, 253.9805, 253.9808, 253.9803, 253.9805, 253.9805, 
    253.9805, 253.9807, 253.9808, 253.981, 253.9809, 253.9814, 253.9812, 
    253.9819, 253.9817, 253.9803, 253.9804, 253.9806, 253.9805, 253.9808, 
    253.9809, 253.981, 253.981, 253.981, 253.9811, 253.981, 253.9811, 
    253.9808, 253.9809, 253.9806, 253.9807, 253.9807, 253.9806, 253.9807, 
    253.9809, 253.9809, 253.9809, 253.981, 253.9808, 253.9815, 253.9811, 
    253.9805, 253.9806, 253.9806, 253.9806, 253.9809, 253.9808, 253.9811, 
    253.981, 253.9811, 253.9811, 253.9811, 253.981, 253.9809, 253.9808, 
    253.9807, 253.9806, 253.9806, 253.9807, 253.9809, 253.981, 253.981, 
    253.9811, 253.9808, 253.9809, 253.9809, 253.981, 253.9807, 253.981, 
    253.9807, 253.9807, 253.9808, 253.9809, 253.981, 253.981, 253.981, 
    253.9809, 253.9809, 253.9808, 253.9807, 253.9807, 253.9806, 253.9807, 
    253.9807, 253.9809, 253.981, 253.9812, 253.9812, 253.9814, 253.9812, 
    253.9815, 253.9813, 253.9816, 253.981, 253.9813, 253.9808, 253.9808, 
    253.9809, 253.9811, 253.981, 253.9812, 253.9809, 253.9807, 253.9807, 
    253.9806, 253.9807, 253.9807, 253.9807, 253.9807, 253.9809, 253.9808, 
    253.9811, 253.9812, 253.9814, 253.9816, 253.9818, 253.9819, 253.9819, 
    253.9819 ;

 TSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSOI =
  254.5829, 254.5844, 254.5841, 254.5853, 254.5846, 254.5854, 254.5832, 
    254.5844, 254.5836, 254.583, 254.5875, 254.5853, 254.5899, 254.5885, 
    254.5921, 254.5897, 254.5926, 254.5921, 254.5938, 254.5933, 254.5954, 
    254.594, 254.5966, 254.5951, 254.5953, 254.594, 254.5858, 254.5872, 
    254.5857, 254.5859, 254.5858, 254.5846, 254.584, 254.5828, 254.583, 
    254.5839, 254.586, 254.5853, 254.5871, 254.5871, 254.5891, 254.5882, 
    254.5915, 254.5906, 254.5933, 254.5926, 254.5933, 254.5931, 254.5933, 
    254.5923, 254.5927, 254.5918, 254.5883, 254.5893, 254.5863, 254.5844, 
    254.5833, 254.5824, 254.5825, 254.5827, 254.5839, 254.5851, 254.5859, 
    254.5865, 254.5871, 254.5887, 254.5896, 254.5917, 254.5913, 254.5919, 
    254.5926, 254.5936, 254.5934, 254.5938, 254.5919, 254.5932, 254.5911, 
    254.5917, 254.5871, 254.5855, 254.5847, 254.5841, 254.5826, 254.5837, 
    254.5832, 254.5843, 254.5849, 254.5846, 254.5865, 254.5858, 254.5897, 
    254.588, 254.5925, 254.5914, 254.5927, 254.5921, 254.5932, 254.5922, 
    254.594, 254.5944, 254.5941, 254.5952, 254.5921, 254.5933, 254.5846, 
    254.5846, 254.5849, 254.5838, 254.5837, 254.5828, 254.5836, 254.584, 
    254.5849, 254.5855, 254.586, 254.5871, 254.5884, 254.5902, 254.5915, 
    254.5924, 254.5918, 254.5923, 254.5918, 254.5915, 254.5942, 254.5927, 
    254.595, 254.5949, 254.5938, 254.5949, 254.5847, 254.5844, 254.5833, 
    254.5841, 254.5827, 254.5835, 254.5839, 254.5857, 254.5862, 254.5865, 
    254.5873, 254.5882, 254.5898, 254.5913, 254.5926, 254.5925, 254.5925, 
    254.5928, 254.5921, 254.5929, 254.5931, 254.5927, 254.5949, 254.5943, 
    254.5949, 254.5945, 254.5845, 254.5849, 254.5847, 254.5852, 254.5848, 
    254.5864, 254.5868, 254.5891, 254.5882, 254.5896, 254.5883, 254.5885, 
    254.5896, 254.5884, 254.5912, 254.5892, 254.5928, 254.5909, 254.593, 
    254.5926, 254.5932, 254.5937, 254.5944, 254.5957, 254.5954, 254.5965, 
    254.5857, 254.5863, 254.5863, 254.5869, 254.5874, 254.5885, 254.5902, 
    254.5896, 254.5908, 254.591, 254.5892, 254.5903, 254.5867, 254.5873, 
    254.587, 254.5857, 254.5897, 254.5877, 254.5915, 254.5904, 254.5937, 
    254.592, 254.5952, 254.5966, 254.5979, 254.5994, 254.5867, 254.5862, 
    254.587, 254.5881, 254.5891, 254.5904, 254.5906, 254.5908, 254.5915, 
    254.592, 254.5909, 254.5922, 254.5874, 254.5899, 254.5861, 254.5872, 
    254.588, 254.5877, 254.5895, 254.59, 254.5917, 254.5908, 254.5962, 
    254.5938, 254.6006, 254.5986, 254.5861, 254.5867, 254.5887, 254.5877, 
    254.5905, 254.5912, 254.5918, 254.5925, 254.5926, 254.593, 254.5923, 
    254.593, 254.5905, 254.5916, 254.5885, 254.5892, 254.5889, 254.5885, 
    254.5897, 254.5909, 254.591, 254.5914, 254.5924, 254.5906, 254.5965, 
    254.5927, 254.5873, 254.5884, 254.5886, 254.5882, 254.5912, 254.5901, 
    254.593, 254.5922, 254.5935, 254.5929, 254.5928, 254.5919, 254.5914, 
    254.5901, 254.5891, 254.5882, 254.5884, 254.5893, 254.591, 254.5926, 
    254.5922, 254.5934, 254.5903, 254.5916, 254.5911, 254.5924, 254.5896, 
    254.5919, 254.589, 254.5892, 254.5901, 254.5917, 254.5921, 254.5925, 
    254.5922, 254.591, 254.5909, 254.59, 254.5898, 254.5892, 254.5887, 
    254.5891, 254.5896, 254.591, 254.5923, 254.5937, 254.5941, 254.5957, 
    254.5943, 254.5965, 254.5946, 254.5979, 254.5921, 254.5946, 254.5901, 
    254.5906, 254.5914, 254.5935, 254.5924, 254.5937, 254.5909, 254.5894, 
    254.589, 254.5883, 254.589, 254.589, 254.5897, 254.5894, 254.5911, 
    254.5902, 254.5928, 254.5937, 254.5963, 254.5979, 254.5996, 254.6004, 
    254.6006, 254.6007,
  255.718, 255.7195, 255.7192, 255.7205, 255.7198, 255.7206, 255.7183, 
    255.7196, 255.7188, 255.7182, 255.7228, 255.7205, 255.7254, 255.7239, 
    255.7276, 255.7251, 255.7282, 255.7276, 255.7294, 255.7289, 255.7311, 
    255.7296, 255.7323, 255.7308, 255.731, 255.7296, 255.721, 255.7225, 
    255.7209, 255.7211, 255.7211, 255.7198, 255.7192, 255.7179, 255.7181, 
    255.7191, 255.7212, 255.7205, 255.7224, 255.7224, 255.7244, 255.7235, 
    255.727, 255.726, 255.7289, 255.7282, 255.7289, 255.7287, 255.7289, 
    255.7278, 255.7282, 255.7273, 255.7236, 255.7247, 255.7215, 255.7196, 
    255.7184, 255.7175, 255.7176, 255.7178, 255.7191, 255.7203, 255.7212, 
    255.7218, 255.7224, 255.7241, 255.725, 255.7272, 255.7268, 255.7274, 
    255.7281, 255.7291, 255.729, 255.7294, 255.7274, 255.7287, 255.7266, 
    255.7272, 255.7224, 255.7207, 255.7199, 255.7193, 255.7177, 255.7188, 
    255.7184, 255.7194, 255.7201, 255.7198, 255.7218, 255.721, 255.7251, 
    255.7233, 255.728, 255.7269, 255.7283, 255.7276, 255.7288, 255.7277, 
    255.7296, 255.73, 255.7297, 255.7308, 255.7276, 255.7289, 255.7197, 
    255.7198, 255.72, 255.7189, 255.7189, 255.7179, 255.7188, 255.7191, 
    255.7201, 255.7207, 255.7212, 255.7224, 255.7237, 255.7256, 255.727, 
    255.7279, 255.7273, 255.7278, 255.7273, 255.727, 255.7298, 255.7282, 
    255.7307, 255.7305, 255.7294, 255.7305, 255.7198, 255.7195, 255.7185, 
    255.7193, 255.7178, 255.7186, 255.7191, 255.721, 255.7214, 255.7218, 
    255.7226, 255.7235, 255.7252, 255.7267, 255.7281, 255.728, 255.7281, 
    255.7284, 255.7276, 255.7285, 255.7286, 255.7283, 255.7305, 255.7299, 
    255.7305, 255.7301, 255.7196, 255.7201, 255.7199, 255.7204, 255.72, 
    255.7216, 255.7221, 255.7244, 255.7235, 255.725, 255.7237, 255.7239, 
    255.725, 255.7238, 255.7266, 255.7246, 255.7284, 255.7263, 255.7285, 
    255.7281, 255.7288, 255.7293, 255.7301, 255.7314, 255.7311, 255.7322, 
    255.7209, 255.7216, 255.7215, 255.7222, 255.7227, 255.7239, 255.7257, 
    255.725, 255.7263, 255.7265, 255.7246, 255.7258, 255.722, 255.7226, 
    255.7223, 255.7209, 255.7251, 255.723, 255.727, 255.7258, 255.7292, 
    255.7275, 255.7309, 255.7323, 255.7337, 255.7352, 255.7219, 255.7215, 
    255.7223, 255.7234, 255.7245, 255.7259, 255.726, 255.7263, 255.727, 
    255.7276, 255.7263, 255.7277, 255.7227, 255.7253, 255.7213, 255.7225, 
    255.7234, 255.723, 255.7249, 255.7254, 255.7272, 255.7263, 255.7319, 
    255.7294, 255.7365, 255.7345, 255.7213, 255.722, 255.7241, 255.7231, 
    255.726, 255.7267, 255.7273, 255.728, 255.7281, 255.7286, 255.7278, 
    255.7285, 255.7259, 255.7271, 255.7238, 255.7246, 255.7243, 255.7239, 
    255.7251, 255.7264, 255.7264, 255.7268, 255.7279, 255.726, 255.7322, 
    255.7283, 255.7226, 255.7238, 255.724, 255.7235, 255.7266, 255.7255, 
    255.7286, 255.7277, 255.7291, 255.7284, 255.7283, 255.7274, 255.7269, 
    255.7255, 255.7244, 255.7236, 255.7238, 255.7247, 255.7265, 255.7281, 
    255.7278, 255.729, 255.7258, 255.7271, 255.7266, 255.728, 255.725, 
    255.7274, 255.7243, 255.7246, 255.7255, 255.7272, 255.7276, 255.728, 
    255.7278, 255.7265, 255.7263, 255.7255, 255.7252, 255.7246, 255.724, 
    255.7245, 255.725, 255.7265, 255.7279, 255.7293, 255.7297, 255.7314, 
    255.73, 255.7322, 255.7302, 255.7337, 255.7276, 255.7302, 255.7255, 
    255.726, 255.7269, 255.7291, 255.728, 255.7293, 255.7263, 255.7247, 
    255.7244, 255.7236, 255.7244, 255.7243, 255.7251, 255.7248, 255.7266, 
    255.7256, 255.7283, 255.7293, 255.732, 255.7337, 255.7355, 255.7363, 
    255.7365, 255.7366,
  257.2901, 257.2917, 257.2914, 257.2928, 257.292, 257.2929, 257.2904, 
    257.2918, 257.2909, 257.2902, 257.2953, 257.2928, 257.2981, 257.2964, 
    257.3006, 257.2978, 257.3011, 257.3005, 257.3025, 257.3019, 257.3044, 
    257.3027, 257.3056, 257.304, 257.3042, 257.3027, 257.2934, 257.295, 
    257.2932, 257.2935, 257.2934, 257.292, 257.2914, 257.2899, 257.2902, 
    257.2912, 257.2936, 257.2928, 257.2949, 257.2948, 257.2971, 257.2961, 
    257.2999, 257.2988, 257.3019, 257.3011, 257.3019, 257.3017, 257.3019, 
    257.3007, 257.3012, 257.3002, 257.2962, 257.2974, 257.2939, 257.2918, 
    257.2905, 257.2895, 257.2896, 257.2899, 257.2912, 257.2925, 257.2935, 
    257.2942, 257.2948, 257.2967, 257.2977, 257.3001, 257.2997, 257.3004, 
    257.3011, 257.3022, 257.302, 257.3025, 257.3004, 257.3018, 257.2994, 
    257.3001, 257.2949, 257.293, 257.2922, 257.2915, 257.2898, 257.291, 
    257.2905, 257.2916, 257.2923, 257.292, 257.2942, 257.2933, 257.2978, 
    257.2959, 257.301, 257.2997, 257.3013, 257.3005, 257.3018, 257.3006, 
    257.3027, 257.3031, 257.3029, 257.304, 257.3006, 257.3019, 257.292, 
    257.292, 257.2923, 257.2911, 257.291, 257.2899, 257.2909, 257.2913, 
    257.2924, 257.293, 257.2936, 257.2949, 257.2963, 257.2983, 257.2998, 
    257.3008, 257.3002, 257.3008, 257.3002, 257.2999, 257.303, 257.3012, 
    257.3039, 257.3037, 257.3025, 257.3037, 257.2921, 257.2917, 257.2906, 
    257.2915, 257.2898, 257.2907, 257.2913, 257.2933, 257.2938, 257.2942, 
    257.295, 257.2961, 257.2979, 257.2996, 257.3011, 257.301, 257.301, 
    257.3014, 257.3005, 257.3015, 257.3017, 257.3012, 257.3037, 257.303, 
    257.3037, 257.3033, 257.2918, 257.2924, 257.2921, 257.2927, 257.2923, 
    257.294, 257.2946, 257.2971, 257.2961, 257.2977, 257.2962, 257.2965, 
    257.2977, 257.2963, 257.2995, 257.2973, 257.3014, 257.2992, 257.3015, 
    257.3011, 257.3018, 257.3024, 257.3032, 257.3046, 257.3043, 257.3055, 
    257.2932, 257.2939, 257.2939, 257.2946, 257.2952, 257.2964, 257.2984, 
    257.2977, 257.2991, 257.2993, 257.2973, 257.2985, 257.2944, 257.2951, 
    257.2947, 257.2933, 257.2979, 257.2955, 257.2999, 257.2986, 257.3023, 
    257.3004, 257.3041, 257.3057, 257.3072, 257.3089, 257.2943, 257.2939, 
    257.2948, 257.296, 257.2971, 257.2986, 257.2988, 257.2991, 257.2998, 
    257.3005, 257.2992, 257.3006, 257.2952, 257.298, 257.2937, 257.295, 
    257.2959, 257.2955, 257.2976, 257.2981, 257.3001, 257.2991, 257.3053, 
    257.3025, 257.3102, 257.308, 257.2937, 257.2944, 257.2967, 257.2956, 
    257.2988, 257.2995, 257.3002, 257.301, 257.3011, 257.3016, 257.3008, 
    257.3015, 257.2986, 257.3, 257.2964, 257.2973, 257.2969, 257.2964, 
    257.2978, 257.2992, 257.2993, 257.2997, 257.3009, 257.2988, 257.3056, 
    257.3013, 257.2951, 257.2964, 257.2966, 257.2961, 257.2995, 257.2982, 
    257.3016, 257.3007, 257.3022, 257.3014, 257.3013, 257.3004, 257.2998, 
    257.2983, 257.2971, 257.2961, 257.2964, 257.2974, 257.2993, 257.3011, 
    257.3007, 257.302, 257.2985, 257.3, 257.2994, 257.3009, 257.2977, 
    257.3004, 257.297, 257.2973, 257.2982, 257.3, 257.3005, 257.301, 
    257.3007, 257.2993, 257.2991, 257.2982, 257.2979, 257.2972, 257.2966, 
    257.2971, 257.2977, 257.2993, 257.3008, 257.3024, 257.3028, 257.3046, 
    257.3031, 257.3056, 257.3034, 257.3072, 257.3005, 257.3034, 257.2982, 
    257.2988, 257.2998, 257.3021, 257.3009, 257.3023, 257.2991, 257.2974, 
    257.297, 257.2962, 257.297, 257.297, 257.2978, 257.2975, 257.2994, 
    257.2984, 257.3013, 257.3023, 257.3054, 257.3072, 257.3092, 257.31, 
    257.3103, 257.3104,
  259.3257, 259.3275, 259.3271, 259.3285, 259.3277, 259.3286, 259.3261, 
    259.3275, 259.3266, 259.3259, 259.3311, 259.3286, 259.3339, 259.3322, 
    259.3365, 259.3336, 259.337, 259.3364, 259.3384, 259.3378, 259.3403, 
    259.3386, 259.3416, 259.3399, 259.3402, 259.3386, 259.3291, 259.3308, 
    259.329, 259.3292, 259.3291, 259.3278, 259.3271, 259.3256, 259.3259, 
    259.3269, 259.3293, 259.3286, 259.3306, 259.3306, 259.3329, 259.3318, 
    259.3357, 259.3346, 259.3378, 259.337, 259.3378, 259.3376, 259.3378, 
    259.3366, 259.3371, 259.3361, 259.332, 259.3332, 259.3297, 259.3275, 
    259.3262, 259.3252, 259.3253, 259.3256, 259.3269, 259.3282, 259.3292, 
    259.3299, 259.3306, 259.3325, 259.3336, 259.3359, 259.3355, 259.3362, 
    259.3369, 259.3381, 259.3379, 259.3384, 259.3362, 259.3377, 259.3353, 
    259.3359, 259.3307, 259.3288, 259.3279, 259.3272, 259.3254, 259.3266, 
    259.3262, 259.3273, 259.328, 259.3277, 259.3299, 259.329, 259.3336, 
    259.3316, 259.3369, 259.3356, 259.3372, 259.3364, 259.3377, 259.3365, 
    259.3386, 259.3391, 259.3388, 259.34, 259.3364, 259.3378, 259.3277, 
    259.3277, 259.328, 259.3268, 259.3267, 259.3256, 259.3266, 259.327, 
    259.3281, 259.3287, 259.3293, 259.3306, 259.3321, 259.3342, 259.3357, 
    259.3367, 259.3361, 259.3366, 259.336, 259.3357, 259.3389, 259.3371, 
    259.3398, 259.3397, 259.3384, 259.3397, 259.3278, 259.3274, 259.3263, 
    259.3272, 259.3255, 259.3264, 259.327, 259.329, 259.3295, 259.33, 
    259.3308, 259.3319, 259.3338, 259.3354, 259.337, 259.3369, 259.3369, 
    259.3372, 259.3364, 259.3374, 259.3376, 259.3371, 259.3396, 259.3389, 
    259.3397, 259.3392, 259.3275, 259.3281, 259.3278, 259.3284, 259.328, 
    259.3298, 259.3303, 259.3329, 259.3318, 259.3335, 259.332, 259.3323, 
    259.3336, 259.3321, 259.3353, 259.3331, 259.3372, 259.335, 259.3374, 
    259.337, 259.3377, 259.3383, 259.3391, 259.3406, 259.3402, 259.3415, 
    259.329, 259.3297, 259.3297, 259.3304, 259.331, 259.3322, 259.3343, 
    259.3335, 259.3349, 259.3352, 259.3331, 259.3344, 259.3302, 259.3308, 
    259.3305, 259.329, 259.3336, 259.3313, 259.3357, 259.3344, 259.3382, 
    259.3363, 259.3401, 259.3416, 259.3432, 259.3449, 259.3301, 259.3296, 
    259.3305, 259.3318, 259.3329, 259.3345, 259.3347, 259.3349, 259.3357, 
    259.3363, 259.335, 259.3365, 259.331, 259.3339, 259.3294, 259.3307, 
    259.3317, 259.3313, 259.3334, 259.3339, 259.336, 259.3349, 259.3412, 
    259.3384, 259.3463, 259.3441, 259.3294, 259.3301, 259.3325, 259.3314, 
    259.3346, 259.3354, 259.3361, 259.3369, 259.337, 259.3375, 259.3367, 
    259.3374, 259.3345, 259.3358, 259.3322, 259.3331, 259.3327, 259.3322, 
    259.3336, 259.3351, 259.3351, 259.3355, 259.3368, 259.3346, 259.3416, 
    259.3372, 259.3309, 259.3322, 259.3324, 259.3318, 259.3353, 259.334, 
    259.3375, 259.3365, 259.338, 259.3373, 259.3372, 259.3362, 259.3356, 
    259.3341, 259.3329, 259.3319, 259.3322, 259.3332, 259.3351, 259.337, 
    259.3366, 259.3379, 259.3344, 259.3358, 259.3353, 259.3368, 259.3335, 
    259.3362, 259.3328, 259.3331, 259.334, 259.3359, 259.3364, 259.3368, 
    259.3365, 259.3352, 259.335, 259.334, 259.3337, 259.333, 259.3324, 
    259.3329, 259.3335, 259.3352, 259.3367, 259.3383, 259.3387, 259.3406, 
    259.3391, 259.3416, 259.3394, 259.3432, 259.3364, 259.3394, 259.3341, 
    259.3347, 259.3357, 259.338, 259.3368, 259.3383, 259.335, 259.3332, 
    259.3328, 259.332, 259.3328, 259.3328, 259.3336, 259.3333, 259.3352, 
    259.3342, 259.3372, 259.3383, 259.3414, 259.3433, 259.3452, 259.3461, 
    259.3463, 259.3465,
  261.4341, 261.4354, 261.4351, 261.4362, 261.4356, 261.4362, 261.4343, 
    261.4354, 261.4347, 261.4342, 261.4382, 261.4362, 261.4403, 261.439, 
    261.4423, 261.4401, 261.4427, 261.4422, 261.4437, 261.4433, 261.4452, 
    261.4439, 261.4463, 261.4449, 261.4451, 261.4439, 261.4366, 261.438, 
    261.4365, 261.4367, 261.4366, 261.4356, 261.4351, 261.434, 261.4342, 
    261.435, 261.4368, 261.4362, 261.4378, 261.4377, 261.4395, 261.4387, 
    261.4417, 261.4409, 261.4433, 261.4427, 261.4433, 261.4431, 261.4433, 
    261.4424, 261.4428, 261.442, 261.4388, 261.4398, 261.437, 261.4354, 
    261.4344, 261.4336, 261.4337, 261.4339, 261.435, 261.436, 261.4367, 
    261.4372, 261.4377, 261.4392, 261.4401, 261.4419, 261.4416, 261.4421, 
    261.4426, 261.4435, 261.4434, 261.4438, 261.4421, 261.4432, 261.4414, 
    261.4419, 261.4378, 261.4364, 261.4357, 261.4352, 261.4338, 261.4347, 
    261.4344, 261.4352, 261.4358, 261.4355, 261.4373, 261.4366, 261.4401, 
    261.4386, 261.4426, 261.4416, 261.4428, 261.4422, 261.4432, 261.4423, 
    261.4439, 261.4443, 261.444, 261.445, 261.4423, 261.4433, 261.4355, 
    261.4356, 261.4358, 261.4348, 261.4348, 261.434, 261.4347, 261.435, 
    261.4359, 261.4363, 261.4368, 261.4378, 261.4389, 261.4405, 261.4417, 
    261.4424, 261.442, 261.4424, 261.4419, 261.4417, 261.4442, 261.4428, 
    261.4448, 261.4447, 261.4438, 261.4447, 261.4356, 261.4353, 261.4344, 
    261.4352, 261.4339, 261.4346, 261.435, 261.4366, 261.437, 261.4373, 
    261.4379, 261.4388, 261.4402, 261.4415, 261.4427, 261.4426, 261.4426, 
    261.4429, 261.4422, 261.443, 261.4431, 261.4428, 261.4447, 261.4442, 
    261.4447, 261.4444, 261.4354, 261.4359, 261.4356, 261.4361, 261.4358, 
    261.4371, 261.4376, 261.4395, 261.4387, 261.44, 261.4389, 261.4391, 
    261.44, 261.4389, 261.4414, 261.4397, 261.4429, 261.4412, 261.443, 
    261.4427, 261.4432, 261.4437, 261.4443, 261.4454, 261.4452, 261.4461, 
    261.4365, 261.4371, 261.437, 261.4376, 261.4381, 261.439, 261.4406, 
    261.44, 261.4411, 261.4413, 261.4397, 261.4406, 261.4375, 261.438, 
    261.4377, 261.4366, 261.4401, 261.4383, 261.4417, 261.4407, 261.4436, 
    261.4422, 261.445, 261.4463, 261.4474, 261.4488, 261.4374, 261.437, 
    261.4377, 261.4387, 261.4395, 261.4408, 261.4409, 261.4411, 261.4417, 
    261.4422, 261.4412, 261.4423, 261.4381, 261.4403, 261.4369, 261.4379, 
    261.4386, 261.4383, 261.4399, 261.4403, 261.4419, 261.4411, 261.446, 
    261.4438, 261.4499, 261.4482, 261.4369, 261.4374, 261.4392, 261.4384, 
    261.4408, 261.4414, 261.442, 261.4426, 261.4427, 261.4431, 261.4424, 
    261.443, 261.4408, 261.4418, 261.439, 261.4397, 261.4394, 261.439, 
    261.4401, 261.4412, 261.4412, 261.4416, 261.4425, 261.4409, 261.4462, 
    261.4429, 261.438, 261.439, 261.4391, 261.4387, 261.4414, 261.4404, 
    261.443, 261.4423, 261.4435, 261.4429, 261.4428, 261.4421, 261.4416, 
    261.4405, 261.4395, 261.4388, 261.439, 261.4398, 261.4413, 261.4427, 
    261.4424, 261.4434, 261.4406, 261.4418, 261.4413, 261.4425, 261.44, 
    261.4421, 261.4394, 261.4397, 261.4404, 261.4419, 261.4422, 261.4426, 
    261.4424, 261.4413, 261.4411, 261.4404, 261.4402, 261.4396, 261.4391, 
    261.4396, 261.44, 261.4413, 261.4424, 261.4437, 261.444, 261.4455, 
    261.4443, 261.4462, 261.4445, 261.4475, 261.4423, 261.4445, 261.4404, 
    261.4409, 261.4417, 261.4435, 261.4425, 261.4437, 261.4411, 261.4398, 
    261.4395, 261.4388, 261.4395, 261.4394, 261.44, 261.4398, 261.4413, 
    261.4405, 261.4428, 261.4437, 261.446, 261.4475, 261.449, 261.4497, 
    261.4499, 261.45,
  262.7637, 262.7643, 262.7642, 262.7646, 262.7643, 262.7646, 262.7638, 
    262.7643, 262.764, 262.7638, 262.7654, 262.7646, 262.7662, 262.7657, 
    262.767, 262.7661, 262.7672, 262.767, 262.7675, 262.7674, 262.7682, 
    262.7676, 262.7686, 262.768, 262.7681, 262.7676, 262.7647, 262.7653, 
    262.7647, 262.7648, 262.7647, 262.7643, 262.7641, 262.7637, 262.7638, 
    262.7641, 262.7648, 262.7646, 262.7652, 262.7652, 262.7659, 262.7656, 
    262.7668, 262.7664, 262.7674, 262.7672, 262.7674, 262.7673, 262.7674, 
    262.767, 262.7672, 262.7668, 262.7656, 262.766, 262.7649, 262.7643, 
    262.7639, 262.7635, 262.7636, 262.7637, 262.7641, 262.7645, 262.7648, 
    262.765, 262.7652, 262.7658, 262.7661, 262.7668, 262.7667, 262.7669, 
    262.7671, 262.7675, 262.7674, 262.7676, 262.7669, 262.7673, 262.7666, 
    262.7668, 262.7652, 262.7646, 262.7644, 262.7642, 262.7636, 262.764, 
    262.7639, 262.7642, 262.7644, 262.7643, 262.765, 262.7647, 262.7661, 
    262.7655, 262.7671, 262.7667, 262.7672, 262.7669, 262.7674, 262.767, 
    262.7676, 262.7678, 262.7677, 262.768, 262.767, 262.7674, 262.7643, 
    262.7643, 262.7644, 262.764, 262.764, 262.7637, 262.764, 262.7641, 
    262.7644, 262.7646, 262.7648, 262.7652, 262.7657, 262.7663, 262.7667, 
    262.7671, 262.7668, 262.767, 262.7668, 262.7668, 262.7677, 262.7672, 
    262.768, 262.7679, 262.7676, 262.7679, 262.7643, 262.7643, 262.7639, 
    262.7642, 262.7637, 262.7639, 262.7641, 262.7647, 262.7649, 262.765, 
    262.7653, 262.7656, 262.7662, 262.7667, 262.7671, 262.7671, 262.7671, 
    262.7672, 262.767, 262.7672, 262.7673, 262.7672, 262.7679, 262.7677, 
    262.7679, 262.7678, 262.7643, 262.7644, 262.7643, 262.7645, 262.7644, 
    262.765, 262.7651, 262.7659, 262.7656, 262.7661, 262.7656, 262.7657, 
    262.7661, 262.7657, 262.7666, 262.766, 262.7672, 262.7665, 262.7673, 
    262.7671, 262.7673, 262.7675, 262.7678, 262.7682, 262.7681, 262.7685, 
    262.7647, 262.7649, 262.7649, 262.7651, 262.7653, 262.7657, 262.7663, 
    262.7661, 262.7665, 262.7666, 262.7659, 262.7663, 262.7651, 262.7653, 
    262.7652, 262.7647, 262.7661, 262.7654, 262.7668, 262.7664, 262.7675, 
    262.7669, 262.7681, 262.7686, 262.769, 262.7696, 262.765, 262.7649, 
    262.7652, 262.7655, 262.7659, 262.7664, 262.7664, 262.7665, 262.7668, 
    262.7669, 262.7665, 262.767, 262.7653, 262.7662, 262.7648, 262.7652, 
    262.7655, 262.7654, 262.7661, 262.7662, 262.7668, 262.7665, 262.7684, 
    262.7676, 262.77, 262.7693, 262.7648, 262.765, 262.7658, 262.7654, 
    262.7664, 262.7667, 262.7668, 262.7671, 262.7671, 262.7673, 262.767, 
    262.7673, 262.7664, 262.7668, 262.7657, 262.766, 262.7658, 262.7657, 
    262.7661, 262.7665, 262.7665, 262.7667, 262.7671, 262.7664, 262.7686, 
    262.7672, 262.7653, 262.7657, 262.7657, 262.7656, 262.7666, 262.7662, 
    262.7673, 262.767, 262.7675, 262.7672, 262.7672, 262.7669, 262.7667, 
    262.7663, 262.7659, 262.7656, 262.7657, 262.766, 262.7666, 262.7671, 
    262.767, 262.7674, 262.7663, 262.7668, 262.7666, 262.7671, 262.7661, 
    262.7669, 262.7658, 262.766, 262.7662, 262.7668, 262.7669, 262.7671, 
    262.767, 262.7666, 262.7665, 262.7662, 262.7661, 262.7659, 262.7657, 
    262.7659, 262.7661, 262.7666, 262.767, 262.7675, 262.7677, 262.7682, 
    262.7678, 262.7686, 262.7679, 262.769, 262.767, 262.7679, 262.7662, 
    262.7664, 262.7667, 262.7675, 262.7671, 262.7675, 262.7665, 262.766, 
    262.7659, 262.7656, 262.7659, 262.7658, 262.7661, 262.766, 262.7666, 
    262.7663, 262.7672, 262.7675, 262.7685, 262.769, 262.7697, 262.7699, 
    262.77, 262.77,
  263.1172, 263.1173, 263.1172, 263.1173, 263.1173, 263.1173, 263.1172, 
    263.1173, 263.1172, 263.1172, 263.1174, 263.1173, 263.1176, 263.1175, 
    263.1177, 263.1176, 263.1177, 263.1177, 263.1178, 263.1177, 263.1179, 
    263.1178, 263.1179, 263.1178, 263.1179, 263.1178, 263.1173, 263.1174, 
    263.1173, 263.1174, 263.1173, 263.1173, 263.1172, 263.1172, 263.1172, 
    263.1172, 263.1174, 263.1173, 263.1174, 263.1174, 263.1175, 263.1175, 
    263.1176, 263.1176, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1175, 263.1175, 263.1174, 263.1173, 
    263.1172, 263.1172, 263.1172, 263.1172, 263.1172, 263.1173, 263.1174, 
    263.1174, 263.1174, 263.1175, 263.1176, 263.1176, 263.1176, 263.1177, 
    263.1177, 263.1178, 263.1177, 263.1178, 263.1177, 263.1177, 263.1176, 
    263.1176, 263.1174, 263.1173, 263.1173, 263.1173, 263.1172, 263.1172, 
    263.1172, 263.1173, 263.1173, 263.1173, 263.1174, 263.1173, 263.1176, 
    263.1175, 263.1177, 263.1176, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 263.1177, 263.1173, 
    263.1173, 263.1173, 263.1172, 263.1172, 263.1172, 263.1172, 263.1172, 
    263.1173, 263.1173, 263.1174, 263.1174, 263.1175, 263.1176, 263.1176, 
    263.1177, 263.1177, 263.1177, 263.1176, 263.1176, 263.1178, 263.1177, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1173, 263.1173, 263.1172, 
    263.1173, 263.1172, 263.1172, 263.1172, 263.1173, 263.1174, 263.1174, 
    263.1174, 263.1175, 263.1176, 263.1176, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1173, 263.1173, 263.1173, 263.1173, 263.1173, 
    263.1174, 263.1174, 263.1175, 263.1175, 263.1176, 263.1175, 263.1175, 
    263.1176, 263.1175, 263.1176, 263.1175, 263.1177, 263.1176, 263.1177, 
    263.1177, 263.1177, 263.1178, 263.1178, 263.1179, 263.1179, 263.1179, 
    263.1173, 263.1174, 263.1174, 263.1174, 263.1174, 263.1175, 263.1176, 
    263.1176, 263.1176, 263.1176, 263.1175, 263.1176, 263.1174, 263.1174, 
    263.1174, 263.1173, 263.1176, 263.1175, 263.1176, 263.1176, 263.1178, 
    263.1177, 263.1178, 263.1179, 263.118, 263.1181, 263.1174, 263.1174, 
    263.1174, 263.1175, 263.1175, 263.1176, 263.1176, 263.1176, 263.1176, 
    263.1177, 263.1176, 263.1177, 263.1174, 263.1176, 263.1174, 263.1174, 
    263.1175, 263.1175, 263.1176, 263.1176, 263.1176, 263.1176, 263.1179, 
    263.1178, 263.1181, 263.118, 263.1174, 263.1174, 263.1175, 263.1175, 
    263.1176, 263.1176, 263.1176, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1176, 263.1176, 263.1175, 263.1175, 263.1175, 263.1175, 
    263.1176, 263.1176, 263.1176, 263.1176, 263.1177, 263.1176, 263.1179, 
    263.1177, 263.1174, 263.1175, 263.1175, 263.1175, 263.1176, 263.1176, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1176, 
    263.1176, 263.1175, 263.1175, 263.1175, 263.1175, 263.1176, 263.1177, 
    263.1177, 263.1177, 263.1176, 263.1176, 263.1176, 263.1177, 263.1176, 
    263.1177, 263.1175, 263.1175, 263.1176, 263.1176, 263.1177, 263.1177, 
    263.1177, 263.1176, 263.1176, 263.1176, 263.1176, 263.1175, 263.1175, 
    263.1175, 263.1176, 263.1176, 263.1177, 263.1178, 263.1178, 263.1179, 
    263.1178, 263.1179, 263.1178, 263.118, 263.1177, 263.1178, 263.1176, 
    263.1176, 263.1176, 263.1177, 263.1177, 263.1178, 263.1176, 263.1175, 
    263.1175, 263.1175, 263.1175, 263.1175, 263.1176, 263.1175, 263.1176, 
    263.1176, 263.1177, 263.1178, 263.1179, 263.118, 263.1181, 263.1181, 
    263.1181, 263.1181,
  263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15 ;

 TSOI_10CM =
  263.7267, 263.7377, 263.7356, 263.7444, 263.7395, 263.7453, 263.729, 
    263.7381, 263.7323, 263.7278, 263.7614, 263.7448, 263.7787, 263.7681, 
    263.7947, 263.777, 263.7983, 263.7943, 263.8065, 263.803, 263.8186, 
    263.8081, 263.8267, 263.8161, 263.8178, 263.8078, 263.7482, 263.7594, 
    263.7475, 263.7491, 263.7484, 263.7396, 263.7352, 263.7259, 263.7276, 
    263.7344, 263.7498, 263.7446, 263.7578, 263.7575, 263.772, 263.7655, 
    263.79, 263.783, 263.8032, 263.7981, 263.8029, 263.8015, 263.8029, 
    263.7955, 263.7987, 263.7921, 263.7667, 263.7742, 263.7519, 263.7383, 
    263.7294, 263.723, 263.7239, 263.7256, 263.7344, 263.7427, 263.7491, 
    263.7533, 263.7574, 263.7699, 263.7765, 263.7914, 263.7887, 263.7932, 
    263.7976, 263.8048, 263.8036, 263.8069, 263.7932, 263.8022, 263.7872, 
    263.7913, 263.7585, 263.746, 263.7406, 263.736, 263.7246, 263.7325, 
    263.7294, 263.7368, 263.7414, 263.7391, 263.7534, 263.7478, 263.7769, 
    263.7645, 263.7971, 263.7893, 263.799, 263.794, 263.8025, 263.7949, 
    263.808, 263.8109, 263.809, 263.8165, 263.7944, 263.8029, 263.739, 
    263.7394, 263.7412, 263.7334, 263.733, 263.7259, 263.7322, 263.7349, 
    263.7417, 263.7457, 263.7495, 263.758, 263.7673, 263.7804, 263.7898, 
    263.7961, 263.7922, 263.7956, 263.7918, 263.79, 263.8098, 263.7987, 
    263.8154, 263.8145, 263.8069, 263.8146, 263.7397, 263.7375, 263.7299, 
    263.7359, 263.7251, 263.7311, 263.7346, 263.748, 263.7509, 263.7536, 
    263.759, 263.7658, 263.7778, 263.7883, 263.7979, 263.7971, 263.7974, 
    263.7995, 263.7943, 263.8004, 263.8014, 263.7987, 263.8144, 263.8099, 
    263.8145, 263.8116, 263.7382, 263.7419, 263.7399, 263.7436, 263.741, 
    263.7526, 263.7561, 263.7723, 263.7657, 263.7762, 263.7668, 263.7684, 
    263.7766, 263.7672, 263.7877, 263.7738, 263.7996, 263.7857, 263.8005, 
    263.7978, 263.8022, 263.8062, 263.8111, 263.8203, 263.8182, 263.8258, 
    263.7473, 263.752, 263.7516, 263.7566, 263.7603, 263.7681, 263.7808, 
    263.776, 263.7848, 263.7866, 263.7733, 263.7814, 263.7552, 263.7595, 
    263.757, 263.7477, 263.7771, 263.7621, 263.7899, 263.7817, 263.8056, 
    263.7937, 263.817, 263.8269, 263.8363, 263.8471, 263.7546, 263.7514, 
    263.7572, 263.7651, 263.7725, 263.7823, 263.7833, 263.7851, 263.7898, 
    263.7938, 263.7856, 263.7948, 263.7604, 263.7784, 263.7502, 263.7587, 
    263.7647, 263.7621, 263.7755, 263.7787, 263.7916, 263.7849, 263.8244, 
    263.807, 263.8554, 263.8419, 263.7503, 263.7546, 263.7696, 263.7625, 
    263.7829, 263.7879, 263.792, 263.7972, 263.7978, 263.8009, 263.7958, 
    263.8007, 263.7823, 263.7905, 263.7679, 263.7734, 263.7709, 263.7681, 
    263.7767, 263.7858, 263.786, 263.7889, 263.7971, 263.783, 263.8267, 
    263.7997, 263.7594, 263.7676, 263.7688, 263.7657, 263.7874, 263.7795, 
    263.8008, 263.7951, 263.8045, 263.7998, 263.7991, 263.7931, 263.7893, 
    263.7799, 263.7722, 263.7661, 263.7675, 263.7742, 263.7863, 263.7978, 
    263.7953, 263.8038, 263.7814, 263.7908, 263.7872, 263.7966, 263.7759, 
    263.7935, 263.7714, 263.7733, 263.7794, 263.7914, 263.7941, 263.7969, 
    263.7952, 263.7867, 263.7852, 263.7792, 263.7775, 263.7729, 263.7691, 
    263.7726, 263.7762, 263.7867, 263.796, 263.8062, 263.8087, 263.8206, 
    263.8109, 263.8268, 263.8132, 263.8367, 263.7945, 263.8129, 263.7796, 
    263.7832, 263.7897, 263.8046, 263.7966, 263.8059, 263.7852, 263.7744, 
    263.7716, 263.7665, 263.7718, 263.7713, 263.7764, 263.7748, 263.787, 
    263.7805, 263.7991, 263.8059, 263.825, 263.8367, 263.8487, 263.8539, 
    263.8555, 263.8562 ;

 TSOI_ICE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TV =
  254.0113, 254.0121, 254.012, 254.0126, 254.0123, 254.0127, 254.0115, 
    254.0122, 254.0117, 254.0114, 254.0139, 254.0127, 254.0152, 254.0144, 
    254.0164, 254.015, 254.0166, 254.0163, 254.0173, 254.017, 254.0181, 
    254.0174, 254.0188, 254.018, 254.0181, 254.0173, 254.0129, 254.0137, 
    254.0129, 254.013, 254.0129, 254.0123, 254.0119, 254.0113, 254.0114, 
    254.0119, 254.013, 254.0126, 254.0136, 254.0136, 254.0147, 254.0142, 
    254.016, 254.0155, 254.017, 254.0166, 254.017, 254.0169, 254.017, 
    254.0164, 254.0167, 254.0162, 254.0143, 254.0148, 254.0132, 254.0122, 
    254.0115, 254.0111, 254.0111, 254.0112, 254.0119, 254.0125, 254.013, 
    254.0133, 254.0136, 254.0145, 254.015, 254.0161, 254.0159, 254.0163, 
    254.0166, 254.0171, 254.017, 254.0173, 254.0163, 254.0169, 254.0158, 
    254.0161, 254.0136, 254.0128, 254.0123, 254.012, 254.0112, 254.0117, 
    254.0115, 254.0121, 254.0124, 254.0123, 254.0133, 254.0129, 254.015, 
    254.0141, 254.0166, 254.016, 254.0167, 254.0163, 254.017, 254.0164, 
    254.0174, 254.0176, 254.0174, 254.018, 254.0164, 254.017, 254.0123, 
    254.0123, 254.0124, 254.0118, 254.0118, 254.0113, 254.0117, 254.0119, 
    254.0125, 254.0127, 254.013, 254.0136, 254.0143, 254.0153, 254.016, 
    254.0165, 254.0162, 254.0164, 254.0162, 254.016, 254.0175, 254.0167, 
    254.0179, 254.0179, 254.0173, 254.0179, 254.0123, 254.0121, 254.0116, 
    254.012, 254.0112, 254.0117, 254.0119, 254.0129, 254.0131, 254.0133, 
    254.0137, 254.0142, 254.0151, 254.0159, 254.0166, 254.0166, 254.0166, 
    254.0167, 254.0163, 254.0168, 254.0169, 254.0167, 254.0179, 254.0175, 
    254.0179, 254.0176, 254.0122, 254.0125, 254.0123, 254.0126, 254.0124, 
    254.0132, 254.0135, 254.0147, 254.0142, 254.015, 254.0143, 254.0144, 
    254.015, 254.0143, 254.0158, 254.0148, 254.0167, 254.0157, 254.0168, 
    254.0166, 254.0169, 254.0172, 254.0176, 254.0183, 254.0181, 254.0187, 
    254.0129, 254.0132, 254.0132, 254.0135, 254.0138, 254.0144, 254.0153, 
    254.015, 254.0156, 254.0158, 254.0148, 254.0154, 254.0134, 254.0137, 
    254.0136, 254.0129, 254.015, 254.0139, 254.016, 254.0154, 254.0172, 
    254.0163, 254.018, 254.0188, 254.0195, 254.0203, 254.0134, 254.0132, 
    254.0136, 254.0142, 254.0147, 254.0154, 254.0155, 254.0157, 254.016, 
    254.0163, 254.0157, 254.0164, 254.0138, 254.0152, 254.0131, 254.0137, 
    254.0141, 254.0139, 254.015, 254.0152, 254.0161, 254.0157, 254.0186, 
    254.0173, 254.0209, 254.0199, 254.0131, 254.0134, 254.0145, 254.014, 
    254.0155, 254.0159, 254.0162, 254.0166, 254.0166, 254.0168, 254.0165, 
    254.0168, 254.0154, 254.0161, 254.0144, 254.0148, 254.0146, 254.0144, 
    254.015, 254.0157, 254.0157, 254.0159, 254.0165, 254.0155, 254.0187, 
    254.0167, 254.0137, 254.0143, 254.0145, 254.0142, 254.0158, 254.0152, 
    254.0168, 254.0164, 254.0171, 254.0168, 254.0167, 254.0163, 254.016, 
    254.0153, 254.0147, 254.0143, 254.0144, 254.0148, 254.0157, 254.0166, 
    254.0164, 254.0171, 254.0154, 254.0161, 254.0158, 254.0165, 254.015, 
    254.0162, 254.0146, 254.0148, 254.0152, 254.0161, 254.0163, 254.0165, 
    254.0164, 254.0158, 254.0157, 254.0152, 254.0151, 254.0148, 254.0145, 
    254.0147, 254.015, 254.0158, 254.0165, 254.0172, 254.0174, 254.0183, 
    254.0176, 254.0187, 254.0177, 254.0195, 254.0163, 254.0177, 254.0153, 
    254.0155, 254.016, 254.0171, 254.0165, 254.0172, 254.0157, 254.0148, 
    254.0147, 254.0143, 254.0147, 254.0146, 254.015, 254.0149, 254.0158, 
    254.0153, 254.0167, 254.0172, 254.0186, 254.0195, 254.0204, 254.0208, 
    254.021, 254.021 ;

 TWS =
  NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, NaNf, 
    NaNf, NaNf ;

 T_SCALAR =
  0.1411014, 0.1411097, 0.1411081, 0.1411147, 0.1411111, 0.1411154, 
    0.1411031, 0.1411099, 0.1411056, 0.1411022, 0.1411274, 0.141115, 
    0.141141, 0.141133, 0.1411534, 0.1411396, 0.1411562, 0.1411532, 
    0.1411627, 0.14116, 0.1411718, 0.141164, 0.1411783, 0.1411701, 0.1411713, 
    0.1411637, 0.1411177, 0.1411258, 0.1411172, 0.1411183, 0.1411179, 
    0.1411111, 0.1411076, 0.1411008, 0.1411021, 0.1411072, 0.1411189, 
    0.141115, 0.1411251, 0.1411249, 0.141136, 0.141131, 0.1411499, 0.1411445, 
    0.1411601, 0.1411562, 0.1411599, 0.1411588, 0.1411599, 0.1411541, 
    0.1411566, 0.1411516, 0.1411319, 0.1411376, 0.1411205, 0.1411099, 
    0.1411034, 0.1410986, 0.1410993, 0.1411005, 0.1411072, 0.1411136, 
    0.1411184, 0.1411216, 0.1411248, 0.141134, 0.1411393, 0.1411508, 
    0.1411489, 0.1411523, 0.1411558, 0.1411614, 0.1411605, 0.1411629, 
    0.1411523, 0.1411593, 0.1411478, 0.1411509, 0.1411251, 0.1411161, 
    0.1411117, 0.1411084, 0.1410998, 0.1411057, 0.1411033, 0.141109, 
    0.1411126, 0.1411109, 0.1411217, 0.1411175, 0.1411396, 0.1411301, 
    0.1411554, 0.1411493, 0.1411568, 0.141153, 0.1411595, 0.1411537, 
    0.1411639, 0.141166, 0.1411645, 0.1411704, 0.1411534, 0.1411598, 
    0.1411108, 0.1411111, 0.1411124, 0.1411064, 0.1411061, 0.1411008, 
    0.1411056, 0.1411075, 0.1411128, 0.1411159, 0.1411188, 0.1411252, 
    0.1411323, 0.1411424, 0.1411497, 0.1411546, 0.1411517, 0.1411543, 
    0.1411513, 0.14115, 0.1411652, 0.1411566, 0.1411696, 0.1411689, 
    0.1411629, 0.141169, 0.1411113, 0.1411096, 0.1411038, 0.1411084, 
    0.1411002, 0.1411047, 0.1411072, 0.1411174, 0.1411198, 0.1411218, 
    0.141126, 0.1411312, 0.1411404, 0.1411485, 0.141156, 0.1411555, 
    0.1411556, 0.1411573, 0.1411532, 0.1411579, 0.1411587, 0.1411566, 
    0.1411688, 0.1411653, 0.1411689, 0.1411666, 0.1411102, 0.1411129, 
    0.1411114, 0.1411142, 0.1411122, 0.141121, 0.1411236, 0.1411361, 
    0.1411311, 0.1411392, 0.141132, 0.1411332, 0.1411392, 0.1411324, 
    0.1411479, 0.1411372, 0.1411573, 0.1411463, 0.141158, 0.141156, 
    0.1411594, 0.1411624, 0.1411663, 0.1411733, 0.1411717, 0.1411777, 
    0.1411171, 0.1411206, 0.1411204, 0.1411242, 0.1411269, 0.1411331, 
    0.1411428, 0.1411392, 0.1411459, 0.1411472, 0.141137, 0.1411432, 
    0.141123, 0.1411262, 0.1411244, 0.1411173, 0.1411398, 0.1411282, 
    0.1411498, 0.1411435, 0.1411619, 0.1411527, 0.1411708, 0.1411783, 
    0.1411859, 0.1411941, 0.1411227, 0.1411203, 0.1411247, 0.1411305, 
    0.1411363, 0.1411439, 0.1411447, 0.1411461, 0.1411498, 0.1411529, 
    0.1411464, 0.1411537, 0.1411267, 0.1411409, 0.1411192, 0.1411256, 
    0.1411302, 0.1411283, 0.1411388, 0.1411412, 0.141151, 0.141146, 
    0.1411763, 0.1411629, 0.1412008, 0.1411901, 0.1411194, 0.1411227, 
    0.1411341, 0.1411287, 0.1411445, 0.1411483, 0.1411515, 0.1411554, 
    0.1411559, 0.1411583, 0.1411544, 0.1411582, 0.1411439, 0.1411503, 
    0.1411329, 0.1411371, 0.1411352, 0.1411331, 0.1411397, 0.1411465, 
    0.1411468, 0.141149, 0.1411548, 0.1411445, 0.1411777, 0.1411569, 
    0.1411263, 0.1411324, 0.1411336, 0.1411311, 0.1411479, 0.1411418, 
    0.1411583, 0.1411538, 0.1411611, 0.1411575, 0.1411569, 0.1411523, 
    0.1411494, 0.141142, 0.1411361, 0.1411315, 0.1411326, 0.1411376, 
    0.141147, 0.1411559, 0.1411539, 0.1411606, 0.1411433, 0.1411504, 
    0.1411476, 0.141155, 0.141139, 0.1411521, 0.1411356, 0.1411371, 
    0.1411417, 0.1411508, 0.1411531, 0.1411552, 0.1411539, 0.1411472, 
    0.1411462, 0.1411416, 0.1411402, 0.1411368, 0.1411339, 0.1411365, 
    0.1411392, 0.1411473, 0.1411545, 0.1411624, 0.1411644, 0.1411732, 
    0.1411658, 0.1411778, 0.1411672, 0.1411858, 0.1411531, 0.1411673, 
    0.1411419, 0.1411447, 0.1411495, 0.141161, 0.141155, 0.1411621, 
    0.1411462, 0.1411377, 0.1411358, 0.1411317, 0.1411359, 0.1411355, 
    0.1411395, 0.1411382, 0.1411476, 0.1411426, 0.1411569, 0.1411621, 
    0.141177, 0.1411861, 0.1411956, 0.1411997, 0.141201, 0.1412015,
  0.1476997, 0.1477089, 0.1477071, 0.1477145, 0.1477105, 0.1477152, 
    0.1477017, 0.1477092, 0.1477044, 0.1477007, 0.1477284, 0.1477148, 
    0.1477434, 0.1477345, 0.147757, 0.1477419, 0.1477601, 0.1477568, 
    0.1477673, 0.1477643, 0.1477774, 0.1477687, 0.1477845, 0.1477754, 
    0.1477768, 0.1477684, 0.1477177, 0.1477267, 0.1477171, 0.1477184, 
    0.1477179, 0.1477105, 0.1477066, 0.1476992, 0.1477005, 0.1477061, 
    0.147719, 0.1477147, 0.1477258, 0.1477256, 0.1477379, 0.1477323, 
    0.1477531, 0.1477472, 0.1477644, 0.1477601, 0.1477642, 0.147763, 
    0.1477642, 0.1477578, 0.1477606, 0.147755, 0.1477333, 0.1477396, 
    0.1477208, 0.1477092, 0.147702, 0.1476967, 0.1476975, 0.1476988, 
    0.1477062, 0.1477132, 0.1477185, 0.147722, 0.1477256, 0.1477357, 
    0.1477415, 0.1477542, 0.1477521, 0.1477558, 0.1477597, 0.1477658, 
    0.1477648, 0.1477675, 0.1477559, 0.1477636, 0.1477508, 0.1477543, 
    0.1477259, 0.1477159, 0.1477112, 0.1477075, 0.147698, 0.1477045, 
    0.1477019, 0.1477082, 0.1477121, 0.1477102, 0.1477221, 0.1477175, 
    0.1477419, 0.1477313, 0.1477592, 0.1477526, 0.1477608, 0.1477566, 
    0.1477638, 0.1477574, 0.1477686, 0.147771, 0.1477693, 0.1477758, 
    0.147757, 0.1477641, 0.1477101, 0.1477104, 0.1477119, 0.1477053, 
    0.1477049, 0.1476991, 0.1477043, 0.1477065, 0.1477123, 0.1477157, 
    0.1477189, 0.1477259, 0.1477337, 0.1477449, 0.147753, 0.1477584, 
    0.1477551, 0.147758, 0.1477547, 0.1477533, 0.14777, 0.1477606, 0.1477749, 
    0.1477741, 0.1477676, 0.1477742, 0.1477106, 0.1477088, 0.1477025, 
    0.1477075, 0.1476985, 0.1477034, 0.1477062, 0.1477174, 0.14772, 
    0.1477223, 0.1477268, 0.1477326, 0.1477427, 0.1477516, 0.1477599, 
    0.1477593, 0.1477595, 0.1477613, 0.1477568, 0.147762, 0.1477629, 
    0.1477606, 0.147774, 0.1477702, 0.1477741, 0.1477716, 0.1477094, 
    0.1477125, 0.1477108, 0.1477139, 0.1477117, 0.1477213, 0.1477242, 
    0.147738, 0.1477325, 0.1477414, 0.1477334, 0.1477348, 0.1477414, 
    0.1477339, 0.147751, 0.1477392, 0.1477614, 0.1477492, 0.1477621, 
    0.1477599, 0.1477636, 0.147767, 0.1477713, 0.147779, 0.1477773, 
    0.1477839, 0.147717, 0.1477209, 0.1477207, 0.1477248, 0.1477279, 
    0.1477346, 0.1477453, 0.1477413, 0.1477488, 0.1477502, 0.147739, 
    0.1477458, 0.1477236, 0.1477271, 0.1477251, 0.1477173, 0.1477421, 
    0.1477293, 0.1477531, 0.1477461, 0.1477665, 0.1477562, 0.1477763, 
    0.1477845, 0.1477929, 0.1478021, 0.1477232, 0.1477205, 0.1477254, 
    0.1477319, 0.1477382, 0.1477465, 0.1477475, 0.147749, 0.1477531, 
    0.1477565, 0.1477493, 0.1477573, 0.1477276, 0.1477433, 0.1477194, 
    0.1477264, 0.1477315, 0.1477294, 0.1477409, 0.1477436, 0.1477544, 
    0.1477489, 0.1477824, 0.1477675, 0.1478095, 0.1477976, 0.1477195, 
    0.1477232, 0.1477358, 0.1477298, 0.1477472, 0.1477514, 0.1477549, 
    0.1477593, 0.1477598, 0.1477624, 0.1477582, 0.1477623, 0.1477466, 
    0.1477536, 0.1477345, 0.147739, 0.147737, 0.1477346, 0.1477419, 
    0.1477494, 0.1477498, 0.1477522, 0.1477586, 0.1477472, 0.147784, 
    0.1477609, 0.1477272, 0.147734, 0.1477352, 0.1477325, 0.147751, 
    0.1477442, 0.1477624, 0.1477575, 0.1477656, 0.1477616, 0.1477609, 
    0.1477558, 0.1477526, 0.1477445, 0.147738, 0.1477329, 0.1477341, 
    0.1477397, 0.1477499, 0.1477598, 0.1477576, 0.147765, 0.1477459, 
    0.1477538, 0.1477507, 0.1477588, 0.1477412, 0.1477556, 0.1477374, 
    0.1477391, 0.1477441, 0.1477542, 0.1477567, 0.1477591, 0.1477576, 
    0.1477502, 0.1477491, 0.147744, 0.1477425, 0.1477387, 0.1477355, 
    0.1477384, 0.1477414, 0.1477503, 0.1477582, 0.147767, 0.1477692, 
    0.147779, 0.1477708, 0.1477841, 0.1477724, 0.1477929, 0.1477568, 
    0.1477724, 0.1477444, 0.1477474, 0.1477528, 0.1477654, 0.1477588, 
    0.1477666, 0.1477491, 0.1477398, 0.1477376, 0.1477332, 0.1477377, 
    0.1477373, 0.1477417, 0.1477403, 0.1477506, 0.1477451, 0.1477609, 
    0.1477666, 0.1477831, 0.1477931, 0.1478037, 0.1478082, 0.1478096, 
    0.1478102,
  0.1573442, 0.1573547, 0.1573527, 0.1573611, 0.1573565, 0.157362, 0.1573464, 
    0.1573551, 0.1573496, 0.1573452, 0.1573773, 0.1573615, 0.1573945, 
    0.1573843, 0.1574103, 0.1573928, 0.1574139, 0.15741, 0.1574221, 
    0.1574187, 0.1574339, 0.1574237, 0.1574421, 0.1574316, 0.1574332, 
    0.1574234, 0.1573649, 0.1573753, 0.1573642, 0.1573657, 0.1573651, 
    0.1573565, 0.1573522, 0.1573435, 0.1573451, 0.1573515, 0.1573664, 
    0.1573614, 0.1573742, 0.1573739, 0.1573881, 0.1573817, 0.1574057, 
    0.1573989, 0.1574188, 0.1574138, 0.1574185, 0.1574171, 0.1574185, 
    0.1574112, 0.1574143, 0.1574079, 0.1573829, 0.1573902, 0.1573684, 
    0.1573551, 0.1573467, 0.1573407, 0.1573415, 0.1573431, 0.1573516, 
    0.1573596, 0.1573658, 0.1573698, 0.1573739, 0.1573858, 0.1573924, 
    0.157407, 0.1574045, 0.1574089, 0.1574133, 0.1574204, 0.1574193, 
    0.1574224, 0.1574089, 0.1574178, 0.1574031, 0.1574071, 0.1573744, 
    0.1573628, 0.1573574, 0.1573531, 0.1573422, 0.1573497, 0.1573467, 
    0.1573539, 0.1573584, 0.1573562, 0.15737, 0.1573646, 0.1573928, 
    0.1573806, 0.1574128, 0.1574051, 0.1574146, 0.1574098, 0.1574181, 
    0.1574106, 0.1574236, 0.1574264, 0.1574245, 0.157432, 0.1574102, 
    0.1574185, 0.1573561, 0.1573564, 0.1573581, 0.1573506, 0.1573502, 
    0.1573434, 0.1573495, 0.157352, 0.1573587, 0.1573625, 0.1573662, 
    0.1573744, 0.1573834, 0.1573962, 0.1574056, 0.1574118, 0.157408, 
    0.1574114, 0.1574076, 0.1574059, 0.1574253, 0.1574143, 0.1574309, 
    0.15743, 0.1574225, 0.1574301, 0.1573567, 0.1573546, 0.1573473, 0.157353, 
    0.1573427, 0.1573484, 0.1573517, 0.1573646, 0.1573675, 0.1573701, 
    0.1573754, 0.157382, 0.1573938, 0.157404, 0.1574136, 0.1574129, 
    0.1574131, 0.1574152, 0.15741, 0.157416, 0.157417, 0.1574144, 0.1574299, 
    0.1574255, 0.15743, 0.1574271, 0.1573553, 0.1573588, 0.1573569, 
    0.1573604, 0.1573579, 0.157369, 0.1573724, 0.1573883, 0.1573819, 
    0.1573922, 0.157383, 0.1573846, 0.1573923, 0.1573835, 0.1574034, 
    0.1573897, 0.1574153, 0.1574013, 0.1574161, 0.1574135, 0.1574179, 
    0.1574217, 0.1574267, 0.1574357, 0.1574337, 0.1574413, 0.1573641, 
    0.1573686, 0.1573683, 0.1573731, 0.1573766, 0.1573844, 0.1573967, 
    0.1573921, 0.1574007, 0.1574024, 0.1573894, 0.1573973, 0.1573717, 
    0.1573757, 0.1573734, 0.1573644, 0.157393, 0.1573782, 0.1574057, 
    0.1573977, 0.1574212, 0.1574094, 0.1574325, 0.1574422, 0.1574518, 
    0.1574625, 0.1573711, 0.1573681, 0.1573737, 0.1573812, 0.1573886, 
    0.1573981, 0.1573992, 0.157401, 0.1574057, 0.1574096, 0.1574014, 
    0.1574106, 0.1573764, 0.1573943, 0.1573668, 0.1573749, 0.1573808, 
    0.1573783, 0.1573916, 0.1573947, 0.1574073, 0.1574008, 0.1574397, 
    0.1574224, 0.157471, 0.1574573, 0.157367, 0.1573712, 0.1573857, 
    0.1573788, 0.1573988, 0.1574037, 0.1574078, 0.1574129, 0.1574135, 
    0.1574165, 0.1574116, 0.1574163, 0.1573982, 0.1574063, 0.1573842, 
    0.1573895, 0.1573871, 0.1573844, 0.1573927, 0.1574015, 0.1574019, 
    0.1574047, 0.1574122, 0.1573989, 0.1574416, 0.1574149, 0.1573758, 
    0.1573837, 0.157385, 0.1573819, 0.1574032, 0.1573955, 0.1574164, 
    0.1574108, 0.1574201, 0.1574155, 0.1574148, 0.1574089, 0.1574051, 
    0.1573958, 0.1573882, 0.1573824, 0.1573837, 0.1573902, 0.1574021, 
    0.1574135, 0.1574109, 0.1574194, 0.1573974, 0.1574065, 0.1574029, 
    0.1574123, 0.157392, 0.1574088, 0.1573876, 0.1573895, 0.1573953, 
    0.157407, 0.1574099, 0.1574126, 0.1574109, 0.1574024, 0.1574011, 
    0.1573952, 0.1573935, 0.1573891, 0.1573853, 0.1573887, 0.1573922, 
    0.1574025, 0.1574117, 0.1574218, 0.1574243, 0.1574357, 0.1574262, 
    0.1574417, 0.1574282, 0.1574518, 0.15741, 0.1574281, 0.1573956, 
    0.1573992, 0.1574054, 0.15742, 0.1574123, 0.1574214, 0.1574011, 
    0.1573904, 0.1573878, 0.1573827, 0.1573879, 0.1573875, 0.1573925, 
    0.1573909, 0.1574028, 0.1573964, 0.1574147, 0.1574214, 0.1574404, 
    0.1574521, 0.1574643, 0.1574695, 0.1574712, 0.1574718,
  0.1706327, 0.1706441, 0.1706419, 0.1706511, 0.1706461, 0.1706521, 0.170635, 
    0.1706445, 0.1706385, 0.1706338, 0.1706689, 0.1706516, 0.1706876, 
    0.1706764, 0.1707048, 0.1706858, 0.1707087, 0.1707044, 0.1707177, 
    0.1707139, 0.1707306, 0.1707194, 0.1707396, 0.170728, 0.1707298, 
    0.170719, 0.1706552, 0.1706667, 0.1706545, 0.1706561, 0.1706554, 
    0.1706461, 0.1706414, 0.1706319, 0.1706336, 0.1706407, 0.1706569, 
    0.1706514, 0.1706654, 0.1706651, 0.1706806, 0.1706735, 0.1706998, 
    0.1706923, 0.170714, 0.1707085, 0.1707137, 0.1707122, 0.1707138, 
    0.1707057, 0.1707092, 0.1707021, 0.1706748, 0.1706828, 0.170659, 
    0.1706447, 0.1706354, 0.1706288, 0.1706298, 0.1706315, 0.1706407, 
    0.1706495, 0.1706561, 0.1706606, 0.170665, 0.1706781, 0.1706853, 
    0.1707012, 0.1706985, 0.1707032, 0.170708, 0.1707158, 0.1707146, 
    0.170718, 0.1707032, 0.170713, 0.1706969, 0.1707012, 0.1706658, 
    0.1706529, 0.1706471, 0.1706423, 0.1706305, 0.1706386, 0.1706354, 
    0.1706432, 0.1706481, 0.1706457, 0.1706607, 0.1706548, 0.1706857, 
    0.1706724, 0.1707074, 0.170699, 0.1707095, 0.1707042, 0.1707132, 
    0.1707051, 0.1707193, 0.1707224, 0.1707203, 0.1707285, 0.1707046, 
    0.1707137, 0.1706456, 0.170646, 0.1706478, 0.1706397, 0.1706392, 
    0.1706318, 0.1706384, 0.1706412, 0.1706484, 0.1706526, 0.1706567, 
    0.1706655, 0.1706754, 0.1706894, 0.1706996, 0.1707064, 0.1707022, 
    0.1707059, 0.1707018, 0.1706999, 0.1707212, 0.1707092, 0.1707273, 
    0.1707263, 0.1707181, 0.1707264, 0.1706463, 0.170644, 0.1706361, 
    0.1706423, 0.170631, 0.1706373, 0.1706408, 0.1706549, 0.1706581, 
    0.1706609, 0.1706666, 0.1706739, 0.1706867, 0.1706979, 0.1707083, 
    0.1707075, 0.1707078, 0.1707101, 0.1707044, 0.170711, 0.1707121, 
    0.1707092, 0.1707262, 0.1707213, 0.1707263, 0.1707231, 0.1706448, 
    0.1706486, 0.1706465, 0.1706504, 0.1706476, 0.1706598, 0.1706635, 
    0.1706807, 0.1706737, 0.170685, 0.1706749, 0.1706767, 0.1706852, 
    0.1706755, 0.1706972, 0.1706823, 0.1707101, 0.1706951, 0.1707111, 
    0.1707082, 0.170713, 0.1707173, 0.1707227, 0.1707326, 0.1707303, 
    0.1707387, 0.1706543, 0.1706592, 0.1706589, 0.1706641, 0.170668, 
    0.1706764, 0.1706899, 0.1706849, 0.1706943, 0.1706961, 0.1706819, 
    0.1706906, 0.1706626, 0.170667, 0.1706644, 0.1706547, 0.1706859, 
    0.1706698, 0.1706997, 0.170691, 0.1707166, 0.1707038, 0.170729, 
    0.1707397, 0.1707501, 0.1707619, 0.170662, 0.1706587, 0.1706648, 
    0.1706731, 0.170681, 0.1706915, 0.1706926, 0.1706945, 0.1706997, 
    0.1707039, 0.1706951, 0.170705, 0.1706679, 0.1706874, 0.1706573, 
    0.1706662, 0.1706726, 0.1706699, 0.1706843, 0.1706877, 0.1707014, 
    0.1706944, 0.170737, 0.170718, 0.1707712, 0.1707562, 0.1706575, 0.170662, 
    0.1706779, 0.1706704, 0.1706922, 0.1706976, 0.170702, 0.1707076, 
    0.1707082, 0.1707115, 0.1707061, 0.1707113, 0.1706915, 0.1707004, 
    0.1706762, 0.170682, 0.1706794, 0.1706764, 0.1706856, 0.1706952, 
    0.1706955, 0.1706986, 0.1707071, 0.1706923, 0.1707392, 0.17071, 0.170667, 
    0.1706757, 0.1706771, 0.1706737, 0.170697, 0.1706886, 0.1707115, 
    0.1707053, 0.1707155, 0.1707104, 0.1707096, 0.1707032, 0.1706991, 
    0.1706889, 0.1706807, 0.1706742, 0.1706758, 0.1706828, 0.1706958, 
    0.1707082, 0.1707055, 0.1707147, 0.1706906, 0.1707006, 0.1706967, 
    0.1707069, 0.1706847, 0.1707032, 0.1706799, 0.170682, 0.1706884, 
    0.1707012, 0.1707043, 0.1707073, 0.1707054, 0.1706962, 0.1706947, 
    0.1706883, 0.1706864, 0.1706816, 0.1706775, 0.1706812, 0.1706851, 
    0.1706962, 0.1707063, 0.1707173, 0.1707201, 0.1707327, 0.1707222, 
    0.1707393, 0.1707245, 0.1707503, 0.1707045, 0.1707243, 0.1706887, 
    0.1706926, 0.1706994, 0.1707154, 0.1707069, 0.1707169, 0.1706947, 
    0.170683, 0.1706802, 0.1706746, 0.1706803, 0.1706798, 0.1706853, 
    0.1706835, 0.1706966, 0.1706896, 0.1707096, 0.1707169, 0.1707377, 
    0.1707505, 0.1707637, 0.1707696, 0.1707713, 0.1707721,
  0.1854227, 0.1854323, 0.1854304, 0.1854381, 0.1854339, 0.1854389, 
    0.1854247, 0.1854326, 0.1854276, 0.1854236, 0.185453, 0.1854385, 
    0.1854685, 0.1854591, 0.1854828, 0.185467, 0.185486, 0.1854824, 
    0.1854935, 0.1854903, 0.1855043, 0.1854949, 0.1855118, 0.1855021, 
    0.1855036, 0.1854946, 0.1854414, 0.1854511, 0.1854409, 0.1854422, 
    0.1854416, 0.1854339, 0.18543, 0.1854221, 0.1854235, 0.1854294, 
    0.1854428, 0.1854383, 0.1854499, 0.1854496, 0.1854625, 0.1854567, 
    0.1854786, 0.1854724, 0.1854904, 0.1854859, 0.1854902, 0.1854889, 
    0.1854902, 0.1854835, 0.1854864, 0.1854805, 0.1854578, 0.1854644, 
    0.1854447, 0.1854328, 0.185425, 0.1854195, 0.1854203, 0.1854218, 
    0.1854294, 0.1854367, 0.1854422, 0.1854459, 0.1854496, 0.1854606, 
    0.1854665, 0.1854798, 0.1854775, 0.1854815, 0.1854854, 0.1854919, 
    0.1854909, 0.1854938, 0.1854814, 0.1854896, 0.1854761, 0.1854798, 
    0.1854504, 0.1854396, 0.1854348, 0.1854308, 0.1854209, 0.1854277, 
    0.185425, 0.1854315, 0.1854355, 0.1854335, 0.185446, 0.1854412, 
    0.1854669, 0.1854558, 0.1854849, 0.1854779, 0.1854866, 0.1854822, 
    0.1854898, 0.185483, 0.1854948, 0.1854974, 0.1854956, 0.1855025, 
    0.1854826, 0.1854902, 0.1854335, 0.1854338, 0.1854353, 0.1854286, 
    0.1854281, 0.185422, 0.1854275, 0.1854298, 0.1854358, 0.1854393, 
    0.1854427, 0.18545, 0.1854583, 0.1854699, 0.1854784, 0.1854841, 
    0.1854806, 0.1854836, 0.1854802, 0.1854786, 0.1854964, 0.1854864, 
    0.1855015, 0.1855007, 0.1854938, 0.1855008, 0.185434, 0.1854322, 
    0.1854255, 0.1854307, 0.1854213, 0.1854265, 0.1854295, 0.1854412, 
    0.1854438, 0.1854462, 0.185451, 0.185457, 0.1854677, 0.185477, 0.1854856, 
    0.185485, 0.1854852, 0.1854872, 0.1854824, 0.1854879, 0.1854888, 
    0.1854864, 0.1855006, 0.1854965, 0.1855007, 0.185498, 0.1854328, 
    0.1854359, 0.1854342, 0.1854374, 0.1854352, 0.1854453, 0.1854484, 
    0.1854627, 0.1854569, 0.1854663, 0.1854579, 0.1854593, 0.1854665, 
    0.1854583, 0.1854765, 0.1854641, 0.1854872, 0.1854747, 0.185488, 
    0.1854856, 0.1854896, 0.1854931, 0.1854977, 0.1855059, 0.185504, 
    0.185511, 0.1854407, 0.1854448, 0.1854445, 0.1854489, 0.1854521, 
    0.1854591, 0.1854704, 0.1854661, 0.185474, 0.1854755, 0.1854637, 
    0.1854709, 0.1854476, 0.1854513, 0.1854492, 0.185441, 0.185467, 
    0.1854536, 0.1854785, 0.1854712, 0.1854926, 0.1854819, 0.185503, 
    0.1855119, 0.1855206, 0.1855305, 0.1854471, 0.1854443, 0.1854494, 
    0.1854563, 0.1854629, 0.1854717, 0.1854726, 0.1854742, 0.1854785, 
    0.185482, 0.1854747, 0.1854829, 0.1854521, 0.1854682, 0.1854432, 
    0.1854507, 0.1854559, 0.1854537, 0.1854657, 0.1854685, 0.18548, 
    0.1854741, 0.1855097, 0.1854938, 0.1855382, 0.1855257, 0.1854433, 
    0.1854471, 0.1854604, 0.1854541, 0.1854723, 0.1854767, 0.1854804, 
    0.1854851, 0.1854856, 0.1854884, 0.1854838, 0.1854882, 0.1854717, 
    0.185479, 0.1854589, 0.1854638, 0.1854616, 0.1854591, 0.1854667, 
    0.1854748, 0.185475, 0.1854776, 0.1854848, 0.1854724, 0.1855116, 
    0.1854872, 0.1854513, 0.1854586, 0.1854597, 0.1854569, 0.1854763, 
    0.1854692, 0.1854883, 0.1854832, 0.1854916, 0.1854874, 0.1854868, 
    0.1854814, 0.185478, 0.1854695, 0.1854627, 0.1854573, 0.1854585, 
    0.1854645, 0.1854753, 0.1854856, 0.1854834, 0.185491, 0.1854709, 
    0.1854793, 0.185476, 0.1854845, 0.185466, 0.1854816, 0.185462, 0.1854638, 
    0.1854691, 0.1854798, 0.1854823, 0.1854848, 0.1854833, 0.1854756, 
    0.1854744, 0.185469, 0.1854675, 0.1854634, 0.18546, 0.1854631, 0.1854663, 
    0.1854756, 0.185484, 0.1854932, 0.1854955, 0.1855061, 0.1854973, 
    0.1855117, 0.1854994, 0.1855208, 0.1854826, 0.1854991, 0.1854693, 
    0.1854725, 0.1854783, 0.1854916, 0.1854845, 0.1854929, 0.1854743, 
    0.1854646, 0.1854622, 0.1854576, 0.1854623, 0.185462, 0.1854665, 
    0.185465, 0.1854759, 0.1854701, 0.1854867, 0.1854928, 0.1855102, 
    0.1855209, 0.185532, 0.1855368, 0.1855383, 0.1855389,
  0.1954593, 0.1954633, 0.1954626, 0.1954658, 0.195464, 0.1954661, 0.1954601, 
    0.1954635, 0.1954613, 0.1954597, 0.1954721, 0.195466, 0.1954786, 
    0.1954747, 0.1954847, 0.195478, 0.1954861, 0.1954845, 0.1954892, 
    0.1954879, 0.1954938, 0.1954898, 0.195497, 0.1954929, 0.1954935, 
    0.1954897, 0.1954672, 0.1954713, 0.195467, 0.1954675, 0.1954673, 
    0.195464, 0.1954624, 0.195459, 0.1954596, 0.1954621, 0.1954678, 
    0.1954659, 0.1954708, 0.1954707, 0.1954761, 0.1954737, 0.1954829, 
    0.1954803, 0.1954879, 0.195486, 0.1954878, 0.1954873, 0.1954878, 
    0.195485, 0.1954862, 0.1954837, 0.1954741, 0.1954769, 0.1954686, 
    0.1954636, 0.1954603, 0.195458, 0.1954583, 0.1954589, 0.1954621, 
    0.1954652, 0.1954675, 0.1954691, 0.1954706, 0.1954753, 0.1954778, 
    0.1954834, 0.1954824, 0.1954841, 0.1954858, 0.1954886, 0.1954881, 
    0.1954893, 0.1954841, 0.1954876, 0.1954819, 0.1954834, 0.195471, 
    0.1954664, 0.1954644, 0.1954627, 0.1954585, 0.1954614, 0.1954603, 
    0.195463, 0.1954647, 0.1954639, 0.1954691, 0.1954671, 0.1954779, 
    0.1954733, 0.1954856, 0.1954826, 0.1954863, 0.1954844, 0.1954876, 
    0.1954848, 0.1954898, 0.1954909, 0.1954901, 0.195493, 0.1954846, 
    0.1954878, 0.1954638, 0.195464, 0.1954646, 0.1954618, 0.1954616, 
    0.195459, 0.1954613, 0.1954623, 0.1954648, 0.1954663, 0.1954677, 
    0.1954708, 0.1954743, 0.1954792, 0.1954828, 0.1954852, 0.1954838, 
    0.195485, 0.1954836, 0.1954829, 0.1954905, 0.1954862, 0.1954926, 
    0.1954923, 0.1954894, 0.1954923, 0.1954641, 0.1954633, 0.1954605, 
    0.1954627, 0.1954587, 0.1954609, 0.1954622, 0.1954671, 0.1954682, 
    0.1954692, 0.1954712, 0.1954738, 0.1954783, 0.1954822, 0.1954859, 
    0.1954856, 0.1954857, 0.1954865, 0.1954845, 0.1954869, 0.1954872, 
    0.1954862, 0.1954922, 0.1954905, 0.1954923, 0.1954911, 0.1954635, 
    0.1954649, 0.1954641, 0.1954655, 0.1954646, 0.1954688, 0.1954701, 
    0.1954762, 0.1954737, 0.1954777, 0.1954741, 0.1954748, 0.1954778, 
    0.1954743, 0.195482, 0.1954768, 0.1954865, 0.1954813, 0.1954869, 
    0.1954859, 0.1954876, 0.1954891, 0.195491, 0.1954945, 0.1954937, 
    0.1954966, 0.1954669, 0.1954686, 0.1954685, 0.1954703, 0.1954717, 
    0.1954747, 0.1954794, 0.1954776, 0.1954809, 0.1954816, 0.1954766, 
    0.1954796, 0.1954698, 0.1954714, 0.1954705, 0.195467, 0.195478, 
    0.1954724, 0.1954829, 0.1954798, 0.1954888, 0.1954843, 0.1954932, 
    0.195497, 0.1955007, 0.1955049, 0.1954696, 0.1954684, 0.1954706, 
    0.1954735, 0.1954763, 0.19548, 0.1954804, 0.195481, 0.1954829, 0.1954844, 
    0.1954813, 0.1954847, 0.1954717, 0.1954785, 0.195468, 0.1954711, 
    0.1954733, 0.1954724, 0.1954774, 0.1954786, 0.1954835, 0.195481, 
    0.1954961, 0.1954894, 0.1955082, 0.1955029, 0.195468, 0.1954696, 
    0.1954752, 0.1954725, 0.1954802, 0.1954821, 0.1954837, 0.1954857, 
    0.1954859, 0.195487, 0.1954851, 0.195487, 0.19548, 0.1954831, 0.1954746, 
    0.1954766, 0.1954757, 0.1954747, 0.1954779, 0.1954813, 0.1954814, 
    0.1954825, 0.1954855, 0.1954803, 0.1954969, 0.1954866, 0.1954714, 
    0.1954744, 0.1954749, 0.1954737, 0.1954819, 0.1954789, 0.195487, 
    0.1954848, 0.1954884, 0.1954866, 0.1954864, 0.1954841, 0.1954827, 
    0.1954791, 0.1954762, 0.1954739, 0.1954744, 0.1954769, 0.1954815, 
    0.1954859, 0.1954849, 0.1954881, 0.1954797, 0.1954832, 0.1954818, 
    0.1954854, 0.1954776, 0.1954842, 0.1954759, 0.1954766, 0.1954789, 
    0.1954834, 0.1954845, 0.1954855, 0.1954849, 0.1954816, 0.1954811, 
    0.1954788, 0.1954782, 0.1954765, 0.195475, 0.1954763, 0.1954777, 
    0.1954816, 0.1954852, 0.1954891, 0.19549, 0.1954946, 0.1954909, 0.195497, 
    0.1954917, 0.1955008, 0.1954846, 0.1954916, 0.195479, 0.1954803, 
    0.1954828, 0.1954884, 0.1954854, 0.195489, 0.1954811, 0.195477, 0.195476, 
    0.195474, 0.195476, 0.1954759, 0.1954778, 0.1954772, 0.1954818, 
    0.1954793, 0.1954864, 0.1954889, 0.1954963, 0.1955009, 0.1955055, 
    0.1955076, 0.1955082, 0.1955085,
  0.1982588, 0.1982594, 0.1982593, 0.1982598, 0.1982595, 0.1982598, 
    0.1982589, 0.1982594, 0.1982591, 0.1982588, 0.1982607, 0.1982598, 
    0.1982617, 0.1982611, 0.1982626, 0.1982616, 0.1982628, 0.1982626, 
    0.1982633, 0.1982631, 0.198264, 0.1982634, 0.1982645, 0.1982639, 
    0.198264, 0.1982634, 0.19826, 0.1982606, 0.1982599, 0.19826, 0.19826, 
    0.1982595, 0.1982592, 0.1982587, 0.1982588, 0.1982592, 0.1982601, 
    0.1982598, 0.1982605, 0.1982605, 0.1982613, 0.1982609, 0.1982623, 
    0.1982619, 0.1982631, 0.1982628, 0.1982631, 0.198263, 0.1982631, 
    0.1982627, 0.1982629, 0.1982625, 0.198261, 0.1982614, 0.1982602, 
    0.1982594, 0.1982589, 0.1982586, 0.1982586, 0.1982587, 0.1982592, 
    0.1982597, 0.19826, 0.1982603, 0.1982605, 0.1982612, 0.1982616, 
    0.1982624, 0.1982623, 0.1982625, 0.1982628, 0.1982632, 0.1982631, 
    0.1982633, 0.1982625, 0.198263, 0.1982622, 0.1982624, 0.1982605, 
    0.1982599, 0.1982596, 0.1982593, 0.1982587, 0.1982591, 0.1982589, 
    0.1982593, 0.1982596, 0.1982595, 0.1982603, 0.19826, 0.1982616, 
    0.1982609, 0.1982628, 0.1982623, 0.1982629, 0.1982626, 0.1982631, 
    0.1982626, 0.1982634, 0.1982636, 0.1982635, 0.1982639, 0.1982626, 
    0.1982631, 0.1982595, 0.1982595, 0.1982596, 0.1982592, 0.1982591, 
    0.1982587, 0.1982591, 0.1982592, 0.1982596, 0.1982598, 0.1982601, 
    0.1982605, 0.1982611, 0.1982618, 0.1982623, 0.1982627, 0.1982625, 
    0.1982627, 0.1982625, 0.1982623, 0.1982635, 0.1982629, 0.1982638, 
    0.1982638, 0.1982633, 0.1982638, 0.1982595, 0.1982594, 0.198259, 
    0.1982593, 0.1982587, 0.198259, 0.1982592, 0.19826, 0.1982601, 0.1982603, 
    0.1982606, 0.198261, 0.1982616, 0.1982622, 0.1982628, 0.1982628, 
    0.1982628, 0.1982629, 0.1982626, 0.1982629, 0.198263, 0.1982629, 
    0.1982638, 0.1982635, 0.1982638, 0.1982636, 0.1982594, 0.1982596, 
    0.1982595, 0.1982597, 0.1982596, 0.1982602, 0.1982604, 0.1982613, 
    0.198261, 0.1982616, 0.198261, 0.1982611, 0.1982616, 0.1982611, 
    0.1982622, 0.1982614, 0.1982629, 0.1982621, 0.198263, 0.1982628, 
    0.198263, 0.1982633, 0.1982636, 0.1982641, 0.198264, 0.1982644, 
    0.1982599, 0.1982602, 0.1982602, 0.1982604, 0.1982607, 0.1982611, 
    0.1982618, 0.1982615, 0.1982621, 0.1982622, 0.1982614, 0.1982619, 
    0.1982604, 0.1982606, 0.1982605, 0.1982599, 0.1982616, 0.1982608, 
    0.1982623, 0.1982619, 0.1982633, 0.1982626, 0.1982639, 0.1982645, 
    0.1982651, 0.1982657, 0.1982603, 0.1982602, 0.1982605, 0.1982609, 
    0.1982614, 0.1982619, 0.198262, 0.1982621, 0.1982623, 0.1982626, 
    0.1982621, 0.1982626, 0.1982607, 0.1982617, 0.1982601, 0.1982606, 
    0.1982609, 0.1982608, 0.1982615, 0.1982617, 0.1982624, 0.1982621, 
    0.1982644, 0.1982633, 0.1982662, 0.1982654, 0.1982601, 0.1982603, 
    0.1982612, 0.1982608, 0.1982619, 0.1982622, 0.1982625, 0.1982628, 
    0.1982628, 0.198263, 0.1982627, 0.198263, 0.1982619, 0.1982624, 
    0.1982611, 0.1982614, 0.1982613, 0.1982611, 0.1982616, 0.1982621, 
    0.1982621, 0.1982623, 0.1982628, 0.1982619, 0.1982645, 0.1982629, 
    0.1982606, 0.1982611, 0.1982611, 0.198261, 0.1982622, 0.1982618, 
    0.198263, 0.1982626, 0.1982632, 0.1982629, 0.1982629, 0.1982625, 
    0.1982623, 0.1982618, 0.1982613, 0.198261, 0.1982611, 0.1982614, 
    0.1982621, 0.1982628, 0.1982627, 0.1982631, 0.1982619, 0.1982624, 
    0.1982622, 0.1982627, 0.1982615, 0.1982625, 0.1982613, 0.1982614, 
    0.1982617, 0.1982624, 0.1982626, 0.1982628, 0.1982626, 0.1982622, 
    0.1982621, 0.1982617, 0.1982616, 0.1982614, 0.1982612, 0.1982614, 
    0.1982616, 0.1982622, 0.1982627, 0.1982633, 0.1982634, 0.1982641, 
    0.1982636, 0.1982645, 0.1982637, 0.1982651, 0.1982626, 0.1982637, 
    0.1982618, 0.198262, 0.1982623, 0.1982632, 0.1982627, 0.1982633, 
    0.1982621, 0.1982615, 0.1982613, 0.198261, 0.1982613, 0.1982613, 
    0.1982616, 0.1982615, 0.1982622, 0.1982618, 0.1982629, 0.1982633, 
    0.1982644, 0.1982651, 0.1982658, 0.1982661, 0.1982662, 0.1982663,
  0.1985152, 0.1985152, 0.1985152, 0.1985152, 0.1985152, 0.1985152, 
    0.1985152, 0.1985152, 0.1985152, 0.1985152, 0.1985153, 0.1985152, 
    0.1985153, 0.1985153, 0.1985154, 0.1985153, 0.1985154, 0.1985154, 
    0.1985154, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 
    0.1985154, 0.1985154, 0.1985152, 0.1985153, 0.1985152, 0.1985152, 
    0.1985152, 0.1985152, 0.1985152, 0.1985151, 0.1985152, 0.1985152, 
    0.1985152, 0.1985152, 0.1985152, 0.1985152, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 
    0.1985154, 0.1985154, 0.1985154, 0.1985153, 0.1985153, 0.1985153, 
    0.1985152, 0.1985152, 0.1985152, 0.1985151, 0.1985151, 0.1985151, 
    0.1985152, 0.1985152, 0.1985152, 0.1985152, 0.1985152, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985154, 0.1985154, 
    0.1985154, 0.1985154, 0.1985153, 0.1985154, 0.1985153, 0.1985153, 
    0.1985153, 0.1985152, 0.1985152, 0.1985152, 0.1985151, 0.1985152, 
    0.1985152, 0.1985152, 0.1985152, 0.1985152, 0.1985152, 0.1985152, 
    0.1985153, 0.1985153, 0.1985154, 0.1985153, 0.1985154, 0.1985153, 
    0.1985154, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 
    0.1985154, 0.1985154, 0.1985152, 0.1985152, 0.1985152, 0.1985152, 
    0.1985152, 0.1985151, 0.1985152, 0.1985152, 0.1985152, 0.1985152, 
    0.1985152, 0.1985152, 0.1985153, 0.1985153, 0.1985153, 0.1985154, 
    0.1985153, 0.1985154, 0.1985153, 0.1985153, 0.1985154, 0.1985154, 
    0.1985154, 0.1985154, 0.1985154, 0.1985154, 0.1985152, 0.1985152, 
    0.1985152, 0.1985152, 0.1985151, 0.1985152, 0.1985152, 0.1985152, 
    0.1985152, 0.1985152, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985154, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 
    0.1985154, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 
    0.1985152, 0.1985152, 0.1985152, 0.1985152, 0.1985152, 0.1985152, 
    0.1985152, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985154, 0.1985153, 
    0.1985154, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 
    0.1985154, 0.1985154, 0.1985152, 0.1985152, 0.1985152, 0.1985152, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985152, 0.1985153, 0.1985152, 0.1985152, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985154, 0.1985153, 
    0.1985154, 0.1985154, 0.1985155, 0.1985155, 0.1985152, 0.1985152, 
    0.1985152, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985154, 0.1985153, 0.1985153, 
    0.1985152, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985154, 0.1985154, 0.1985155, 0.1985155, 
    0.1985152, 0.1985152, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985154, 0.1985153, 
    0.1985154, 0.1985154, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 
    0.1985154, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985154, 0.1985154, 0.1985154, 
    0.1985153, 0.1985153, 0.1985153, 0.1985154, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985154, 
    0.1985154, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985154, 0.1985154, 
    0.1985154, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 0.1985155, 
    0.1985154, 0.1985154, 0.1985153, 0.1985153, 0.1985153, 0.1985154, 
    0.1985154, 0.1985154, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985154, 0.1985154, 0.1985154, 0.1985155, 0.1985155, 0.1985155, 
    0.1985155, 0.1985155,
  0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 U10 =
  8.609481, 8.609554, 8.60954, 8.609598, 8.609567, 8.609604, 8.609496, 
    8.609556, 8.609518, 8.609488, 8.609708, 8.609601, 8.609828, 8.609756, 
    8.609936, 8.609816, 8.609961, 8.609934, 8.610017, 8.609993, 8.610095, 
    8.610027, 8.61015, 8.61008, 8.61009, 8.610025, 8.609624, 8.609694, 
    8.609619, 8.60963, 8.609625, 8.609567, 8.609536, 8.609476, 8.609488, 
    8.609531, 8.609634, 8.6096, 8.609688, 8.609686, 8.609784, 8.609738, 
    8.609905, 8.609859, 8.609994, 8.609961, 8.609992, 8.609982, 8.609993, 
    8.609942, 8.609963, 8.609921, 8.609746, 8.609797, 8.609648, 8.609556, 
    8.609499, 8.609457, 8.609463, 8.609473, 8.609532, 8.609589, 8.609631, 
    8.609658, 8.609686, 8.609766, 8.609813, 8.609914, 8.609898, 8.609927, 
    8.609957, 8.610005, 8.609998, 8.610019, 8.609927, 8.609987, 8.609887, 
    8.609915, 8.609688, 8.60961, 8.609571, 8.609543, 8.609468, 8.609519, 
    8.609498, 8.609549, 8.609579, 8.609565, 8.609659, 8.609622, 8.609816, 
    8.609731, 8.609953, 8.6099, 8.609966, 8.609933, 8.609989, 8.609939, 
    8.610026, 8.610045, 8.610032, 8.610084, 8.609936, 8.609992, 8.609564, 
    8.609566, 8.609578, 8.609526, 8.609523, 8.609476, 8.609518, 8.609535, 
    8.609582, 8.609608, 8.609633, 8.609689, 8.60975, 8.609839, 8.609904, 
    8.609947, 8.609921, 8.609943, 8.609919, 8.609906, 8.610038, 8.609963, 
    8.610076, 8.61007, 8.610019, 8.61007, 8.609568, 8.609553, 8.609503, 
    8.609543, 8.60947, 8.60951, 8.609532, 8.609622, 8.609642, 8.60966, 
    8.609695, 8.609741, 8.609822, 8.609894, 8.609959, 8.609954, 8.609956, 
    8.60997, 8.609934, 8.609976, 8.609982, 8.609964, 8.610069, 8.61004, 
    8.61007, 8.61005, 8.609558, 8.609583, 8.60957, 8.609593, 8.609576, 
    8.609653, 8.609674, 8.609784, 8.609739, 8.609812, 8.609747, 8.609758, 
    8.609812, 8.609751, 8.609889, 8.609794, 8.60997, 8.609875, 8.609976, 
    8.609959, 8.609988, 8.610014, 8.610047, 8.610108, 8.610094, 8.610146, 
    8.609618, 8.609649, 8.609648, 8.60968, 8.609704, 8.609757, 8.609843, 
    8.609812, 8.609871, 8.609882, 8.609793, 8.609847, 8.609671, 8.609697, 
    8.609682, 8.60962, 8.609818, 8.609715, 8.609905, 8.60985, 8.61001, 
    8.60993, 8.610086, 8.61015, 8.610215, 8.610286, 8.609667, 8.609646, 
    8.609684, 8.609735, 8.609787, 8.609853, 8.60986, 8.609873, 8.609905, 
    8.609932, 8.609876, 8.609939, 8.609701, 8.609827, 8.609637, 8.609693, 
    8.609733, 8.609715, 8.609808, 8.60983, 8.609916, 8.609872, 8.610134, 
    8.610018, 8.610342, 8.610251, 8.609638, 8.609667, 8.609767, 8.609719, 
    8.609859, 8.609892, 8.60992, 8.609954, 8.609959, 8.609979, 8.609945, 
    8.609978, 8.609854, 8.609909, 8.609756, 8.609794, 8.609776, 8.609757, 
    8.609816, 8.609876, 8.609879, 8.609898, 8.609948, 8.609859, 8.610146, 
    8.609966, 8.609698, 8.609752, 8.609762, 8.60974, 8.609888, 8.609835, 
    8.609979, 8.60994, 8.610003, 8.609972, 8.609967, 8.609927, 8.609901, 
    8.609837, 8.609785, 8.609743, 8.609753, 8.609798, 8.60988, 8.609958, 
    8.609941, 8.609999, 8.609848, 8.60991, 8.609886, 8.60995, 8.609811, 
    8.609924, 8.60978, 8.609794, 8.609834, 8.609914, 8.609934, 8.609952, 
    8.609941, 8.609882, 8.609874, 8.609833, 8.609821, 8.609791, 8.609764, 
    8.609788, 8.609813, 8.609883, 8.609945, 8.610014, 8.610031, 8.610107, 
    8.610044, 8.610147, 8.610056, 8.610214, 8.609934, 8.610056, 8.609837, 
    8.60986, 8.609902, 8.610002, 8.60995, 8.610011, 8.609874, 8.609799, 
    8.609781, 8.609745, 8.609782, 8.609779, 8.609815, 8.609803, 8.609885, 
    8.609841, 8.609966, 8.610011, 8.61014, 8.610217, 8.610298, 8.610332, 
    8.610343, 8.610348 ;

 URBAN_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 URBAN_HEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 VOCFLXT =
  4.009859e-15, 4.010252e-15, 4.010181e-15, 4.010481e-15, 4.010317e-15, 
    4.010512e-15, 4.009954e-15, 4.010264e-15, 4.010068e-15, 4.009899e-15, 
    4.011055e-15, 4.010496e-15, 4.011673e-15, 4.01131e-15, 4.012234e-15, 
    4.011612e-15, 4.012361e-15, 4.012224e-15, 4.012656e-15, 4.012533e-15, 
    4.013069e-15, 4.012714e-15, 4.013362e-15, 4.012989e-15, 4.013044e-15, 
    4.0127e-15, 4.010616e-15, 4.010983e-15, 4.010593e-15, 4.010645e-15, 
    4.010624e-15, 4.010318e-15, 4.010159e-15, 4.009837e-15, 4.009894e-15, 
    4.010137e-15, 4.010669e-15, 4.010494e-15, 4.010952e-15, 4.010942e-15, 
    4.011447e-15, 4.011218e-15, 4.012074e-15, 4.011833e-15, 4.012538e-15, 
    4.012359e-15, 4.012528e-15, 4.012479e-15, 4.012529e-15, 4.012268e-15, 
    4.012379e-15, 4.012152e-15, 4.011259e-15, 4.011519e-15, 4.010742e-15, 
    4.010264e-15, 4.009966e-15, 4.009735e-15, 4.009766e-15, 4.009823e-15, 
    4.010139e-15, 4.01043e-15, 4.010649e-15, 4.010795e-15, 4.01094e-15, 
    4.011357e-15, 4.011597e-15, 4.012119e-15, 4.012032e-15, 4.012185e-15, 
    4.012342e-15, 4.012596e-15, 4.012555e-15, 4.012665e-15, 4.012186e-15, 
    4.012502e-15, 4.01198e-15, 4.012122e-15, 4.010951e-15, 4.010543e-15, 
    4.010345e-15, 4.010193e-15, 4.009789e-15, 4.010071e-15, 4.009965e-15, 
    4.010223e-15, 4.010384e-15, 4.010306e-15, 4.010799e-15, 4.010606e-15, 
    4.011611e-15, 4.011177e-15, 4.012324e-15, 4.01205e-15, 4.01239e-15, 
    4.012218e-15, 4.012511e-15, 4.012248e-15, 4.012709e-15, 4.012806e-15, 
    4.012739e-15, 4.013006e-15, 4.012232e-15, 4.012526e-15, 4.010302e-15, 
    4.010315e-15, 4.010377e-15, 4.010104e-15, 4.010089e-15, 4.009834e-15, 
    4.010065e-15, 4.010155e-15, 4.010395e-15, 4.010532e-15, 4.010665e-15, 
    4.010956e-15, 4.011277e-15, 4.011734e-15, 4.012068e-15, 4.01229e-15, 
    4.012156e-15, 4.012274e-15, 4.012141e-15, 4.012079e-15, 4.012768e-15, 
    4.012379e-15, 4.012968e-15, 4.012936e-15, 4.012667e-15, 4.01294e-15, 
    4.010324e-15, 4.010251e-15, 4.009987e-15, 4.010194e-15, 4.009807e-15, 
    4.010026e-15, 4.010142e-15, 4.010604e-15, 4.010712e-15, 4.010804e-15, 
    4.010992e-15, 4.01123e-15, 4.011646e-15, 4.012013e-15, 4.012352e-15, 
    4.012328e-15, 4.012336e-15, 4.012409e-15, 4.012225e-15, 4.01244e-15, 
    4.012473e-15, 4.012382e-15, 4.012932e-15, 4.012775e-15, 4.012935e-15, 
    4.012834e-15, 4.010275e-15, 4.0104e-15, 4.010332e-15, 4.010458e-15, 
    4.010367e-15, 4.010764e-15, 4.010883e-15, 4.011449e-15, 4.011224e-15, 
    4.01159e-15, 4.011263e-15, 4.01132e-15, 4.01159e-15, 4.011283e-15, 
    4.011987e-15, 4.011499e-15, 4.012412e-15, 4.011913e-15, 4.012443e-15, 
    4.012351e-15, 4.012506e-15, 4.012642e-15, 4.012819e-15, 4.013136e-15, 
    4.013064e-15, 4.013334e-15, 4.010589e-15, 4.010748e-15, 4.010739e-15, 
    4.01091e-15, 4.011035e-15, 4.011313e-15, 4.011753e-15, 4.011589e-15, 
    4.011896e-15, 4.011955e-15, 4.011493e-15, 4.011772e-15, 4.010859e-15, 
    4.011e-15, 4.01092e-15, 4.010598e-15, 4.01162e-15, 4.011091e-15, 
    4.012072e-15, 4.011787e-15, 4.012622e-15, 4.012201e-15, 4.013023e-15, 
    4.013361e-15, 4.013705e-15, 4.014078e-15, 4.010841e-15, 4.010732e-15, 
    4.010931e-15, 4.011199e-15, 4.011462e-15, 4.011803e-15, 4.011841e-15, 
    4.011904e-15, 4.012072e-15, 4.012211e-15, 4.011919e-15, 4.012246e-15, 
    4.011023e-15, 4.011668e-15, 4.010686e-15, 4.010974e-15, 4.011185e-15, 
    4.011098e-15, 4.011572e-15, 4.011682e-15, 4.012127e-15, 4.0119e-15, 
    4.013273e-15, 4.012664e-15, 4.014381e-15, 4.013896e-15, 4.010693e-15, 
    4.010843e-15, 4.01136e-15, 4.011114e-15, 4.011829e-15, 4.012003e-15, 
    4.012149e-15, 4.012327e-15, 4.01235e-15, 4.012456e-15, 4.012282e-15, 
    4.012451e-15, 4.011804e-15, 4.012094e-15, 4.011307e-15, 4.011495e-15, 
    4.01141e-15, 4.011313e-15, 4.011612e-15, 4.011922e-15, 4.011937e-15, 
    4.012035e-15, 4.012296e-15, 4.011832e-15, 4.013336e-15, 4.012391e-15, 
    4.011006e-15, 4.011285e-15, 4.011335e-15, 4.011225e-15, 4.011985e-15, 
    4.011709e-15, 4.012455e-15, 4.012254e-15, 4.012585e-15, 4.01242e-15, 
    4.012395e-15, 4.012186e-15, 4.012053e-15, 4.01172e-15, 4.011451e-15, 
    4.011242e-15, 4.011292e-15, 4.011521e-15, 4.011943e-15, 4.012348e-15, 
    4.012258e-15, 4.01256e-15, 4.011777e-15, 4.0121e-15, 4.011972e-15, 
    4.012308e-15, 4.011583e-15, 4.012174e-15, 4.011429e-15, 4.011496e-15, 
    4.011703e-15, 4.012117e-15, 4.012221e-15, 4.012317e-15, 4.01226e-15, 
    4.011955e-15, 4.011909e-15, 4.0117e-15, 4.011638e-15, 4.011482e-15, 
    4.011349e-15, 4.011468e-15, 4.011593e-15, 4.011958e-15, 4.012284e-15, 
    4.012643e-15, 4.012734e-15, 4.013132e-15, 4.012796e-15, 4.01334e-15, 
    4.01286e-15, 4.0137e-15, 4.012221e-15, 4.012863e-15, 4.011715e-15, 
    4.011841e-15, 4.012059e-15, 4.012578e-15, 4.012306e-15, 4.012628e-15, 
    4.011908e-15, 4.011525e-15, 4.011436e-15, 4.011253e-15, 4.01144e-15, 
    4.011426e-15, 4.011604e-15, 4.011547e-15, 4.011971e-15, 4.011743e-15, 
    4.012393e-15, 4.012627e-15, 4.013303e-15, 4.013712e-15, 4.014144e-15, 
    4.01433e-15, 4.014388e-15, 4.014411e-15 ;

 VOLR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WA =
  4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000 ;

 WASTEHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WF =
  11.11574, 11.16004, 11.15141, 11.18721, 11.16734, 11.19079, 11.12471, 
    11.1618, 11.13811, 11.11972, 11.25687, 11.1888, 11.32778, 11.28419, 
    11.39385, 11.321, 11.40857, 11.39174, 11.44242, 11.42789, 11.49287, 
    11.44913, 11.52662, 11.48241, 11.48933, 11.44769, 11.20247, 11.24838, 
    11.19976, 11.2063, 11.20336, 11.16775, 11.14984, 11.11235, 11.11915, 
    11.14668, 11.20924, 11.18798, 11.24159, 11.24038, 11.30024, 11.27323, 
    11.37411, 11.34538, 11.42849, 11.40756, 11.42751, 11.42146, 11.42759, 
    11.3969, 11.41004, 11.38306, 11.27829, 11.30902, 11.2175, 11.16268, 
    11.12633, 11.10059, 11.10423, 11.11116, 11.14684, 11.18044, 11.20609, 
    11.22327, 11.2402, 11.29158, 11.31881, 11.37993, 11.36888, 11.38759, 
    11.40548, 11.43556, 11.4306, 11.44386, 11.38709, 11.42481, 11.36259, 
    11.37959, 11.24484, 11.19371, 11.17204, 11.15307, 11.10702, 11.13881, 
    11.12628, 11.15611, 11.1751, 11.1657, 11.22374, 11.20116, 11.32043, 
    11.26896, 11.40339, 11.37114, 11.41113, 11.39071, 11.42571, 11.39421, 
    11.4488, 11.46071, 11.45257, 11.48384, 11.39247, 11.42752, 11.16544, 
    11.16697, 11.17411, 11.14277, 11.14085, 11.11216, 11.13768, 11.14856, 
    11.17619, 11.19256, 11.20813, 11.24241, 11.28078, 11.33453, 11.37323, 
    11.39922, 11.38328, 11.39735, 11.38162, 11.37425, 11.45625, 11.41017, 
    11.47934, 11.47551, 11.44418, 11.47594, 11.16805, 11.15924, 11.12868, 
    11.15259, 11.10904, 11.13341, 11.14744, 11.20163, 11.21355, 11.22462, 
    11.2465, 11.27461, 11.32402, 11.36711, 11.40652, 11.40363, 11.40465, 
    11.41346, 11.39164, 11.41705, 11.42132, 11.41016, 11.47499, 11.45645, 
    11.47542, 11.46335, 11.1621, 11.17693, 11.16891, 11.18399, 11.17337, 
    11.22065, 11.23485, 11.30141, 11.27406, 11.3176, 11.27847, 11.2854, 
    11.31903, 11.28059, 11.36474, 11.30766, 11.41381, 11.35668, 11.41739, 
    11.40635, 11.42463, 11.44103, 11.46166, 11.4998, 11.49096, 11.52289, 
    11.19906, 11.21834, 11.21664, 11.23683, 11.25177, 11.2842, 11.33633, 
    11.31671, 11.35274, 11.35998, 11.30525, 11.33884, 11.23125, 11.2486, 
    11.23826, 11.20058, 11.32124, 11.25923, 11.37387, 11.34017, 11.43869, 
    11.38964, 11.4861, 11.52748, 11.56648, 11.61217, 11.22886, 11.21576, 
    11.23923, 11.27176, 11.30198, 11.34223, 11.34634, 11.3539, 11.37347, 
    11.38994, 11.35629, 11.39407, 11.25264, 11.32662, 11.21081, 11.24562, 
    11.26984, 11.2592, 11.31447, 11.32752, 11.38063, 11.35315, 11.51726, 
    11.4445, 11.64701, 11.59023, 11.21118, 11.22882, 11.29033, 11.26104, 
    11.34491, 11.36561, 11.38245, 11.40401, 11.40633, 11.41912, 11.39817, 
    11.41829, 11.34231, 11.37623, 11.28328, 11.30587, 11.29547, 11.28408, 
    11.31926, 11.35682, 11.35762, 11.36968, 11.40372, 11.34525, 11.52669, 
    11.41447, 11.24807, 11.28213, 11.28699, 11.27379, 11.36354, 11.33097, 
    11.4188, 11.39503, 11.434, 11.41462, 11.41177, 11.38692, 11.37146, 
    11.33247, 11.30079, 11.2757, 11.28153, 11.3091, 11.35912, 11.40655, 
    11.39615, 11.43103, 11.33882, 11.37744, 11.36251, 11.40146, 11.31619, 
    11.38881, 11.29767, 11.30564, 11.33033, 11.38007, 11.39108, 11.40285, 
    11.39558, 11.36039, 11.35463, 11.32972, 11.32286, 11.30391, 11.28824, 
    11.30256, 11.31761, 11.3604, 11.39905, 11.44126, 11.4516, 11.50108, 
    11.46081, 11.52732, 11.47078, 11.56874, 11.39301, 11.4691, 11.33145, 
    11.34623, 11.373, 11.43453, 11.40128, 11.44016, 11.3544, 11.31005, 
    11.29859, 11.27722, 11.29907, 11.2973, 11.31822, 11.3115, 11.36182, 
    11.33477, 11.41171, 11.43985, 11.51954, 11.56855, 11.61853, 11.64064, 
    11.64737, 11.65018 ;

 WIND =
  8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267 ;

 WOODC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 WOODC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOODC_LOSS =
  1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11 ;

 WOOD_HARVESTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOOD_HARVESTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WTGQ =
  2.972229e-09, 2.937783e-09, 2.944407e-09, 2.917149e-09, 2.932198e-09, 
    2.914454e-09, 2.965171e-09, 2.936433e-09, 2.954704e-09, 2.969092e-09, 
    2.865886e-09, 2.915947e-09, 2.815969e-09, 2.846382e-09, 2.771391e-09, 
    2.820649e-09, 2.7617e-09, 2.772788e-09, 2.739733e-09, 2.749109e-09, 
    2.707804e-09, 2.73543e-09, 2.686958e-09, 2.714345e-09, 2.710016e-09, 
    2.736352e-09, 2.905714e-09, 2.872008e-09, 2.907738e-09, 2.902868e-09, 
    2.905052e-09, 2.931884e-09, 2.945624e-09, 2.974903e-09, 2.969538e-09, 
    2.948059e-09, 2.900685e-09, 2.916569e-09, 2.876926e-09, 2.877808e-09, 
    2.835087e-09, 2.854165e-09, 2.784521e-09, 2.803912e-09, 2.748717e-09, 
    2.762359e-09, 2.749353e-09, 2.753282e-09, 2.749302e-09, 2.769374e-09, 
    2.760733e-09, 2.77855e-09, 2.850568e-09, 2.828954e-09, 2.894573e-09, 
    2.935763e-09, 2.963896e-09, 2.984242e-09, 2.981346e-09, 2.975842e-09, 
    2.947934e-09, 2.922249e-09, 2.90302e-09, 2.890321e-09, 2.877934e-09, 
    2.841171e-09, 2.822159e-09, 2.780636e-09, 2.788028e-09, 2.775534e-09, 
    2.763725e-09, 2.744152e-09, 2.747352e-09, 2.738807e-09, 2.775865e-09, 
    2.751106e-09, 2.792258e-09, 2.780861e-09, 2.874574e-09, 2.912264e-09, 
    2.928624e-09, 2.943131e-09, 2.979123e-09, 2.954158e-09, 2.963941e-09, 
    2.940793e-09, 2.926299e-09, 2.933447e-09, 2.889975e-09, 2.906696e-09, 
    2.821042e-09, 2.857208e-09, 2.765096e-09, 2.786507e-09, 2.760021e-09, 
    2.773464e-09, 2.750522e-09, 2.77115e-09, 2.735643e-09, 2.728049e-09, 
    2.733233e-09, 2.713449e-09, 2.772303e-09, 2.749352e-09, 2.933648e-09, 
    2.932479e-09, 2.927049e-09, 2.951092e-09, 2.952578e-09, 2.97505e-09, 
    2.955036e-09, 2.946608e-09, 2.925466e-09, 2.913123e-09, 2.901503e-09, 
    2.876329e-09, 2.848805e-09, 2.81133e-09, 2.785107e-09, 2.767844e-09, 
    2.778401e-09, 2.769076e-09, 2.779505e-09, 2.784425e-09, 2.730888e-09, 
    2.760651e-09, 2.716274e-09, 2.718687e-09, 2.738604e-09, 2.718415e-09, 
    2.931659e-09, 2.938395e-09, 2.96206e-09, 2.943503e-09, 2.977522e-09, 
    2.958365e-09, 2.947479e-09, 2.906342e-09, 2.897485e-09, 2.889324e-09, 
    2.873366e-09, 2.853181e-09, 2.818556e-09, 2.789214e-09, 2.763042e-09, 
    2.76494e-09, 2.764271e-09, 2.758495e-09, 2.772853e-09, 2.756154e-09, 
    2.753373e-09, 2.760657e-09, 2.71901e-09, 2.730759e-09, 2.718738e-09, 
    2.726373e-09, 2.936202e-09, 2.924908e-09, 2.930998e-09, 2.91957e-09, 
    2.927609e-09, 2.892249e-09, 2.88184e-09, 2.834271e-09, 2.853574e-09, 
    2.822999e-09, 2.850435e-09, 2.845527e-09, 2.822008e-09, 2.848937e-09, 
    2.79081e-09, 2.829908e-09, 2.758271e-09, 2.796249e-09, 2.755931e-09, 
    2.763154e-09, 2.75122e-09, 2.740631e-09, 2.727445e-09, 2.703493e-09, 
    2.708997e-09, 2.689246e-09, 2.90826e-09, 2.893951e-09, 2.895207e-09, 
    2.880394e-09, 2.869551e-09, 2.846376e-09, 2.810097e-09, 2.823614e-09, 
    2.798916e-09, 2.794017e-09, 2.831587e-09, 2.80838e-09, 2.884468e-09, 
    2.871848e-09, 2.879349e-09, 2.907124e-09, 2.820482e-09, 2.864183e-09, 
    2.784678e-09, 2.807469e-09, 2.742135e-09, 2.774178e-09, 2.712037e-09, 
    2.686436e-09, 2.662858e-09, 2.635889e-09, 2.886214e-09, 2.895858e-09, 
    2.878645e-09, 2.855214e-09, 2.833874e-09, 2.806066e-09, 2.803258e-09, 
    2.79813e-09, 2.78495e-09, 2.773979e-09, 2.79651e-09, 2.771244e-09, 
    2.868935e-09, 2.816762e-09, 2.899521e-09, 2.874006e-09, 2.856584e-09, 
    2.864199e-09, 2.825169e-09, 2.816148e-09, 2.780167e-09, 2.798634e-09, 
    2.6927e-09, 2.738403e-09, 2.615782e-09, 2.648756e-09, 2.899244e-09, 
    2.886248e-09, 2.84205e-09, 2.862882e-09, 2.804234e-09, 2.79022e-09, 
    2.778951e-09, 2.764692e-09, 2.763165e-09, 2.754808e-09, 2.768533e-09, 
    2.755348e-09, 2.806007e-09, 2.783104e-09, 2.847026e-09, 2.831153e-09, 
    2.83843e-09, 2.846461e-09, 2.821844e-09, 2.796152e-09, 2.795613e-09, 
    2.787492e-09, 2.764891e-09, 2.804002e-09, 2.686922e-09, 2.757845e-09, 
    2.87223e-09, 2.847846e-09, 2.844407e-09, 2.853768e-09, 2.791618e-09, 
    2.813771e-09, 2.755012e-09, 2.770611e-09, 2.745159e-09, 2.757738e-09, 
    2.7596e-09, 2.77598e-09, 2.786292e-09, 2.812745e-09, 2.834705e-09, 
    2.852407e-09, 2.848268e-09, 2.828902e-09, 2.794599e-09, 2.763025e-09, 
    2.76987e-09, 2.747074e-09, 2.808392e-09, 2.782295e-09, 2.792313e-09, 
    2.766365e-09, 2.823974e-09, 2.774731e-09, 2.836887e-09, 2.831309e-09, 
    2.814215e-09, 2.780542e-09, 2.773225e-09, 2.765453e-09, 2.770243e-09, 
    2.793741e-09, 2.797637e-09, 2.814628e-09, 2.81936e-09, 2.832522e-09, 
    2.843525e-09, 2.833467e-09, 2.822992e-09, 2.793733e-09, 2.767959e-09, 
    2.74048e-09, 2.733853e-09, 2.702699e-09, 2.727991e-09, 2.686538e-09, 
    2.721678e-09, 2.661509e-09, 2.771945e-09, 2.722736e-09, 2.813444e-09, 
    2.803336e-09, 2.785262e-09, 2.744818e-09, 2.766486e-09, 2.741186e-09, 
    2.79779e-09, 2.828238e-09, 2.836247e-09, 2.851322e-09, 2.835904e-09, 
    2.837151e-09, 2.822563e-09, 2.827232e-09, 2.792774e-09, 2.811161e-09, 
    2.759646e-09, 2.741385e-09, 2.691299e-09, 2.661624e-09, 2.632188e-09, 
    2.619429e-09, 2.615574e-09, 2.613966e-09 ;

 W_SCALAR =
  0.6401832, 0.6417798, 0.6414695, 0.6427562, 0.6420426, 0.6428849, 0.640507, 
    0.6418432, 0.6409903, 0.640327, 0.6452495, 0.6428136, 0.6477738, 
    0.6462242, 0.6501127, 0.6475329, 0.6506321, 0.6500382, 0.6518245, 
    0.6513131, 0.6535952, 0.6520605, 0.6547761, 0.6532288, 0.6534711, 
    0.6520099, 0.643304, 0.6449465, 0.6432067, 0.643441, 0.6433358, 
    0.6420574, 0.6414127, 0.640061, 0.6403065, 0.6412992, 0.6435464, 
    0.6427839, 0.6447043, 0.6446609, 0.6467955, 0.6458336, 0.6494153, 
    0.6483984, 0.6513344, 0.6505968, 0.6512998, 0.6510866, 0.6513026, 
    0.6502206, 0.6506843, 0.6497316, 0.6460138, 0.6471077, 0.6438422, 
    0.6418747, 0.6405657, 0.6396361, 0.6397675, 0.6400182, 0.641305, 
    0.6425135, 0.6434337, 0.6440489, 0.6446547, 0.6464871, 0.6474554, 
    0.649621, 0.6492302, 0.6498919, 0.6505234, 0.651583, 0.6514086, 
    0.6518753, 0.6498743, 0.6512046, 0.6490077, 0.649609, 0.64482, 0.6429896, 
    0.6422113, 0.6415292, 0.6398686, 0.6410156, 0.6405636, 0.6416386, 
    0.6423213, 0.6419837, 0.6440657, 0.6432567, 0.6475128, 0.6456814, 
    0.6504497, 0.6493105, 0.6507226, 0.6500022, 0.6512364, 0.6501257, 
    0.6520488, 0.6524672, 0.6521813, 0.6532789, 0.6500641, 0.6512998, 
    0.6419743, 0.6420293, 0.6422858, 0.641158, 0.641089, 0.6400543, 
    0.6409749, 0.6413668, 0.6423609, 0.6429486, 0.6435069, 0.6447337, 
    0.6461023, 0.6480134, 0.6493843, 0.6503024, 0.6497395, 0.6502365, 
    0.6496809, 0.6494204, 0.6523105, 0.6506886, 0.6531211, 0.6529866, 
    0.6518863, 0.6530018, 0.642068, 0.6417511, 0.6406503, 0.6415119, 
    0.6399416, 0.6408209, 0.6413262, 0.6432738, 0.6437011, 0.6440974, 
    0.6448796, 0.6458828, 0.6476406, 0.6491678, 0.6505601, 0.6504581, 
    0.650494, 0.6508049, 0.6500347, 0.6509312, 0.6510817, 0.6506884, 
    0.6529686, 0.6523176, 0.6529838, 0.6525599, 0.6418541, 0.6423873, 
    0.6420992, 0.6426409, 0.6422593, 0.6439551, 0.6444631, 0.6468369, 
    0.6458631, 0.6474124, 0.6460205, 0.6462673, 0.6474631, 0.6460958, 
    0.6490837, 0.647059, 0.650817, 0.6487983, 0.6509433, 0.6505541, 
    0.6511984, 0.6517754, 0.6525006, 0.6538378, 0.6535283, 0.6546455, 
    0.6431816, 0.6438724, 0.6438115, 0.6445339, 0.645068, 0.6462246, 
    0.6480772, 0.6473809, 0.6486589, 0.6489154, 0.6469735, 0.6481662, 
    0.6443344, 0.6449544, 0.6445853, 0.6432362, 0.6475415, 0.645334, 
    0.649407, 0.6482135, 0.6516932, 0.6499641, 0.6533579, 0.6548058, 
    0.6561664, 0.6577547, 0.6442491, 0.6437799, 0.6446198, 0.645781, 
    0.6468571, 0.6482864, 0.6484324, 0.6487, 0.6493927, 0.6499748, 0.6487847, 
    0.6501206, 0.6450984, 0.6477329, 0.6436026, 0.644848, 0.6457126, 
    0.6453332, 0.6473013, 0.6477646, 0.6496458, 0.6486737, 0.6544487, 
    0.6518974, 0.6589622, 0.6569926, 0.643616, 0.6442475, 0.6464427, 
    0.6453987, 0.6483817, 0.6491148, 0.6497104, 0.6504714, 0.6505534, 
    0.651004, 0.6502655, 0.6509748, 0.6482894, 0.6494902, 0.6461918, 
    0.6469956, 0.6466259, 0.6462203, 0.6474716, 0.6488035, 0.6488317, 
    0.6492585, 0.6504606, 0.6483938, 0.654778, 0.6508398, 0.6449357, 
    0.6461505, 0.6463237, 0.6458534, 0.6490414, 0.6478872, 0.650993, 
    0.6501545, 0.6515281, 0.6508457, 0.6507453, 0.6498682, 0.6493218, 
    0.6479402, 0.6468149, 0.6459216, 0.6461294, 0.6471103, 0.6488849, 
    0.6505609, 0.650194, 0.6514238, 0.6481656, 0.649533, 0.6490048, 
    0.6503816, 0.6473624, 0.6499345, 0.6467041, 0.6469877, 0.6478643, 
    0.6496258, 0.6500149, 0.6504306, 0.6501741, 0.6489298, 0.6487258, 
    0.647843, 0.6475992, 0.6469259, 0.6463683, 0.6468778, 0.6474127, 
    0.6489303, 0.6502963, 0.6517836, 0.6521472, 0.6538825, 0.6524704, 
    0.6547999, 0.6528201, 0.6562449, 0.6500831, 0.6527614, 0.6479042, 
    0.6484284, 0.6493762, 0.6515466, 0.6503752, 0.651745, 0.6487178, 
    0.6471443, 0.6467366, 0.6459759, 0.646754, 0.6466907, 0.6474348, 
    0.6471957, 0.6489806, 0.6480222, 0.6507428, 0.6517341, 0.6545286, 
    0.6562383, 0.6579756, 0.6587418, 0.6589748, 0.6590723,
  0.6386675, 0.6403092, 0.6399902, 0.6413131, 0.6405793, 0.6414454, 
    0.6390004, 0.6403744, 0.6394974, 0.6388153, 0.6438766, 0.6413721, 
    0.6464719, 0.6448788, 0.6488765, 0.6462243, 0.6494105, 0.6487998, 
    0.6506363, 0.6501105, 0.6524565, 0.6508788, 0.6536704, 0.6520798, 
    0.6523289, 0.6508268, 0.6418763, 0.6435651, 0.6417763, 0.6420172, 
    0.6419091, 0.6405946, 0.6399317, 0.6385418, 0.6387942, 0.639815, 
    0.6421255, 0.6413416, 0.6433161, 0.6432715, 0.6454661, 0.6444771, 
    0.6481595, 0.647114, 0.6501324, 0.6493741, 0.6500968, 0.6498777, 
    0.6500997, 0.6489873, 0.6494641, 0.6484846, 0.6446624, 0.6457871, 
    0.6424297, 0.6404067, 0.6390608, 0.6381049, 0.6382401, 0.6384978, 
    0.6398209, 0.6410636, 0.6420097, 0.6426422, 0.6432651, 0.6451491, 
    0.6461446, 0.6483709, 0.6479692, 0.6486494, 0.6492986, 0.6503879, 
    0.6502087, 0.6506884, 0.6486314, 0.649999, 0.6477405, 0.6483586, 
    0.643435, 0.6415531, 0.6407529, 0.6400515, 0.638344, 0.6395234, 
    0.6390586, 0.640164, 0.640866, 0.6405188, 0.6426595, 0.6418278, 
    0.6462035, 0.6443207, 0.6492229, 0.6480517, 0.6495034, 0.6487628, 
    0.6500316, 0.6488898, 0.6508668, 0.6512969, 0.6510031, 0.6521314, 
    0.6488265, 0.6500969, 0.6405091, 0.6405658, 0.6408295, 0.6396698, 
    0.6395988, 0.638535, 0.6394816, 0.6398845, 0.6409066, 0.6415108, 
    0.642085, 0.6433463, 0.6447535, 0.6467182, 0.6481277, 0.6490715, 
    0.6484928, 0.6490037, 0.6484326, 0.6481647, 0.6511359, 0.6494685, 
    0.6519691, 0.6518309, 0.6506998, 0.6518465, 0.6406055, 0.6402797, 
    0.6391478, 0.6400337, 0.638419, 0.6393231, 0.6398427, 0.6418453, 
    0.6422846, 0.6426921, 0.6434963, 0.6445277, 0.6463349, 0.647905, 
    0.6493363, 0.6492315, 0.6492684, 0.649588, 0.6487963, 0.6497179, 
    0.6498726, 0.6494682, 0.6518124, 0.6511432, 0.651828, 0.6513923, 
    0.6403856, 0.6409338, 0.6406376, 0.6411945, 0.6408022, 0.6425458, 
    0.6430681, 0.6455087, 0.6445075, 0.6461003, 0.6446694, 0.644923, 
    0.6461525, 0.6447467, 0.6478186, 0.6457371, 0.6496004, 0.6475252, 
    0.6497304, 0.6493301, 0.6499926, 0.6505857, 0.6513313, 0.6527059, 
    0.6523877, 0.6535362, 0.6417505, 0.6424608, 0.6423981, 0.6431409, 
    0.64369, 0.6448791, 0.6467839, 0.6460679, 0.6473818, 0.6476455, 
    0.6456491, 0.6468754, 0.6429358, 0.6435733, 0.6431937, 0.6418066, 
    0.6462331, 0.6439635, 0.648151, 0.646924, 0.6505012, 0.6487237, 
    0.6522126, 0.6537011, 0.6550996, 0.6567324, 0.6428481, 0.6423657, 
    0.6432292, 0.6444231, 0.6455294, 0.6469989, 0.647149, 0.6474241, 
    0.6481362, 0.6487346, 0.6475112, 0.6488846, 0.6437213, 0.6464298, 
    0.6421834, 0.6434639, 0.6443527, 0.6439627, 0.6459861, 0.6464624, 
    0.6483964, 0.647397, 0.653334, 0.6507111, 0.6579735, 0.6559489, 
    0.6421971, 0.6428464, 0.6451034, 0.64403, 0.6470968, 0.6478506, 
    0.6484628, 0.6492451, 0.6493295, 0.6497928, 0.6490335, 0.6497627, 
    0.647002, 0.6482365, 0.6448455, 0.6456718, 0.6452917, 0.6448748, 
    0.6461613, 0.6475305, 0.6475595, 0.6479983, 0.6492341, 0.6471092, 
    0.6536724, 0.6496239, 0.643554, 0.644803, 0.6449811, 0.6444975, 0.647775, 
    0.6465886, 0.6497815, 0.6489193, 0.6503315, 0.64963, 0.6495268, 
    0.6486251, 0.6480634, 0.646643, 0.645486, 0.6445677, 0.6447812, 
    0.6457898, 0.6476142, 0.6493372, 0.6489601, 0.6502243, 0.6468747, 
    0.6482806, 0.6477374, 0.6491529, 0.646049, 0.6486933, 0.6453722, 
    0.6456637, 0.646565, 0.6483759, 0.6487759, 0.6492032, 0.6489395, 
    0.6476604, 0.6474506, 0.646543, 0.6462924, 0.6456002, 0.6450269, 
    0.6455507, 0.6461007, 0.6476609, 0.6490651, 0.6505942, 0.650968, 
    0.6527518, 0.6513002, 0.6536949, 0.6516597, 0.6551803, 0.648846, 
    0.6515994, 0.6466059, 0.6471449, 0.6481192, 0.6503506, 0.6491463, 
    0.6505544, 0.6474424, 0.6458247, 0.6454055, 0.6446235, 0.6454234, 
    0.6453584, 0.6461233, 0.6458775, 0.6477126, 0.6467273, 0.6495242, 
    0.6505433, 0.653416, 0.6551735, 0.6569594, 0.657747, 0.6579865, 0.6580867,
  0.6424639, 0.6441357, 0.6438108, 0.6451582, 0.6444108, 0.645293, 0.642803, 
    0.6442021, 0.643309, 0.6426144, 0.6477698, 0.6452183, 0.6504147, 
    0.648791, 0.6528661, 0.6501623, 0.6534106, 0.652788, 0.6546607, 
    0.6541244, 0.6565174, 0.6549081, 0.6577559, 0.6561331, 0.6563872, 
    0.654855, 0.6457319, 0.6474525, 0.64563, 0.6458755, 0.6457653, 0.6444263, 
    0.6437513, 0.642336, 0.642593, 0.6436324, 0.6459858, 0.6451873, 
    0.6471987, 0.6471533, 0.6493896, 0.6483817, 0.6521351, 0.6510693, 
    0.6541468, 0.6533735, 0.6541106, 0.6538871, 0.6541135, 0.6529791, 
    0.6534652, 0.6524666, 0.6485705, 0.6497167, 0.6462957, 0.6442351, 
    0.6428643, 0.6418911, 0.6420287, 0.6422911, 0.6436385, 0.644904, 
    0.6458678, 0.6465122, 0.6471468, 0.6490664, 0.650081, 0.6523506, 
    0.6519411, 0.6526346, 0.6532965, 0.6544074, 0.6542246, 0.6547139, 
    0.6526162, 0.6540107, 0.6517079, 0.6523381, 0.6473199, 0.6454027, 
    0.6445876, 0.6438733, 0.6421345, 0.6433355, 0.6428622, 0.6439879, 
    0.6447028, 0.6443492, 0.6465298, 0.6456825, 0.6501412, 0.6482223, 
    0.6532193, 0.6520252, 0.6535054, 0.6527503, 0.654044, 0.6528797, 
    0.6548958, 0.6553345, 0.6550348, 0.6561857, 0.6528151, 0.6541106, 
    0.6443393, 0.644397, 0.6446656, 0.6434846, 0.6434123, 0.6423289, 
    0.6432929, 0.6437032, 0.6447442, 0.6453597, 0.6459445, 0.6472294, 
    0.6486633, 0.6506658, 0.6521026, 0.653065, 0.6524749, 0.6529958, 
    0.6524135, 0.6521404, 0.6551702, 0.6534698, 0.6560202, 0.6558792, 
    0.6547255, 0.6558951, 0.6444375, 0.6441056, 0.6429529, 0.6438551, 
    0.6422109, 0.6431316, 0.6436607, 0.6457003, 0.6461479, 0.646563, 
    0.6473824, 0.6484333, 0.6502751, 0.6518756, 0.653335, 0.6532281, 
    0.6532658, 0.6535916, 0.6527843, 0.6537241, 0.6538818, 0.6534696, 
    0.6558603, 0.6551777, 0.6558762, 0.6554318, 0.6442135, 0.6447718, 
    0.6444702, 0.6450374, 0.6446379, 0.6464139, 0.646946, 0.649433, 
    0.6484126, 0.650036, 0.6485776, 0.6488361, 0.6500891, 0.6486564, 
    0.6517875, 0.6496657, 0.6536043, 0.6514884, 0.6537368, 0.6533287, 
    0.6540043, 0.6546091, 0.6553696, 0.6567718, 0.6564472, 0.6576189, 
    0.6456038, 0.6463273, 0.6462635, 0.6470203, 0.6475797, 0.6487914, 
    0.6507328, 0.650003, 0.6513423, 0.6516111, 0.6495761, 0.650826, 
    0.6468112, 0.6474608, 0.647074, 0.6456609, 0.6501713, 0.6478584, 
    0.6521264, 0.6508755, 0.654523, 0.6527103, 0.6562685, 0.6577871, 
    0.6592143, 0.6608809, 0.6467219, 0.6462305, 0.6471102, 0.6483267, 
    0.6494542, 0.6509519, 0.651105, 0.6513854, 0.6521114, 0.6527215, 
    0.6514741, 0.6528744, 0.6476116, 0.6503718, 0.6460447, 0.6473492, 
    0.6482549, 0.6478576, 0.6499195, 0.6504051, 0.6523767, 0.6513578, 
    0.6574126, 0.6547371, 0.662148, 0.6600811, 0.6460587, 0.6467202, 0.64902, 
    0.6479262, 0.6510518, 0.6518201, 0.6524443, 0.6532421, 0.6533281, 
    0.6538004, 0.6530263, 0.6537699, 0.6509551, 0.6522136, 0.6487571, 
    0.6495993, 0.6492119, 0.6487869, 0.6500981, 0.6514938, 0.6515234, 
    0.6519707, 0.6532307, 0.6510644, 0.6577579, 0.6536283, 0.6474411, 
    0.6487138, 0.6488953, 0.6484025, 0.6517431, 0.6505336, 0.6537889, 
    0.6529098, 0.6543499, 0.6536345, 0.6535292, 0.6526098, 0.6520371, 
    0.6505891, 0.6494099, 0.648474, 0.6486917, 0.6497195, 0.6515791, 
    0.6533359, 0.6529513, 0.6542405, 0.6508253, 0.6522585, 0.6517048, 
    0.653148, 0.6499836, 0.6526793, 0.6492938, 0.649591, 0.6505096, 
    0.6523558, 0.6527636, 0.6531993, 0.6529304, 0.6516262, 0.6514124, 
    0.6504872, 0.6502318, 0.6495262, 0.6489419, 0.6494759, 0.6500364, 
    0.6516267, 0.6530585, 0.6546178, 0.654999, 0.6568187, 0.6553379, 
    0.6577809, 0.6557045, 0.6592966, 0.6528351, 0.655643, 0.6505513, 
    0.6511007, 0.6520941, 0.6543693, 0.6531412, 0.6545773, 0.651404, 
    0.6497551, 0.6493279, 0.648531, 0.6493461, 0.6492798, 0.6500595, 
    0.6498089, 0.6516795, 0.650675, 0.6535266, 0.6545659, 0.6574963, 
    0.6592897, 0.6611126, 0.6619167, 0.6621613, 0.6622636,
  0.6480097, 0.649733, 0.649398, 0.6507874, 0.6500167, 0.6509264, 0.6483591, 
    0.6498015, 0.6488808, 0.6481648, 0.6534818, 0.6508494, 0.6562126, 
    0.6545359, 0.6587454, 0.6559519, 0.6593083, 0.6586647, 0.6606008, 
    0.6600463, 0.6625215, 0.6608567, 0.6638032, 0.6621239, 0.6623868, 
    0.6608018, 0.6513792, 0.6531543, 0.651274, 0.6515272, 0.6514136, 
    0.6500327, 0.6493367, 0.6478779, 0.6481428, 0.6492141, 0.6516411, 
    0.6508173, 0.6528924, 0.6528456, 0.6551539, 0.6541134, 0.65799, 
    0.6568887, 0.6600695, 0.6592699, 0.6600319, 0.6598009, 0.660035, 
    0.6588623, 0.6593648, 0.6583326, 0.6543084, 0.6554918, 0.6519607, 
    0.6498355, 0.6484224, 0.6474194, 0.6475613, 0.6478316, 0.6492204, 
    0.6505253, 0.6515193, 0.6521841, 0.6528388, 0.6548203, 0.655868, 
    0.6582127, 0.6577895, 0.6585062, 0.6591904, 0.6603389, 0.6601499, 
    0.6606558, 0.6584871, 0.6599287, 0.6575485, 0.6581998, 0.6530175, 
    0.6510396, 0.6501989, 0.6494625, 0.6476703, 0.6489081, 0.6484202, 
    0.6495806, 0.6503178, 0.6499532, 0.6522022, 0.6513281, 0.6559301, 
    0.6539489, 0.6591106, 0.6578764, 0.6594063, 0.6586257, 0.6599631, 
    0.6587595, 0.660844, 0.6612977, 0.6609877, 0.6621783, 0.6586928, 
    0.660032, 0.649943, 0.6500025, 0.6502794, 0.6490617, 0.6489872, 
    0.6478706, 0.6488642, 0.6492872, 0.6503605, 0.6509952, 0.6515984, 
    0.6529242, 0.6544041, 0.656472, 0.6579564, 0.658951, 0.6583411, 
    0.6588796, 0.6582777, 0.6579955, 0.6611278, 0.6593695, 0.6620071, 
    0.6618612, 0.6606678, 0.6618776, 0.6500442, 0.649702, 0.6485137, 
    0.6494437, 0.647749, 0.6486978, 0.6492433, 0.6513465, 0.6518083, 
    0.6522365, 0.653082, 0.6541667, 0.6560684, 0.6577218, 0.6592302, 
    0.6591197, 0.6591586, 0.6594955, 0.6586609, 0.6596324, 0.6597955, 
    0.6593692, 0.6618416, 0.6611356, 0.6618581, 0.6613984, 0.6498132, 
    0.650389, 0.6500779, 0.6506628, 0.6502508, 0.6520827, 0.6526317, 
    0.6551988, 0.6541454, 0.6558214, 0.6543157, 0.6545826, 0.6558764, 
    0.654397, 0.6576308, 0.6554391, 0.6595086, 0.6573218, 0.6596456, 
    0.6592236, 0.6599221, 0.6605475, 0.661334, 0.6627847, 0.6624488, 
    0.6636615, 0.651247, 0.6519933, 0.6519275, 0.6527083, 0.6532856, 
    0.6545363, 0.6565411, 0.6557873, 0.6571708, 0.6574485, 0.6553466, 
    0.6566374, 0.6524926, 0.6531629, 0.6527637, 0.6513059, 0.6559612, 
    0.6535733, 0.657981, 0.6566886, 0.6604584, 0.6585844, 0.6622639, 
    0.6638355, 0.6653132, 0.6670395, 0.6524004, 0.6518934, 0.6528011, 
    0.6540566, 0.6552206, 0.6567675, 0.6569256, 0.6572153, 0.6579654, 
    0.658596, 0.657307, 0.658754, 0.6533185, 0.6561683, 0.6517018, 0.6530478, 
    0.6539826, 0.6535724, 0.6557012, 0.6562027, 0.6582396, 0.6571867, 
    0.6634479, 0.6606798, 0.6683527, 0.6662109, 0.6517163, 0.6523986, 
    0.6547723, 0.6536432, 0.6568706, 0.6576645, 0.6583095, 0.659134, 
    0.659223, 0.6597113, 0.658911, 0.6596797, 0.6567708, 0.6580711, 0.654501, 
    0.6553704, 0.6549705, 0.6545317, 0.6558856, 0.6573274, 0.6573579, 
    0.6578201, 0.6591223, 0.6568837, 0.6638052, 0.6595333, 0.6531426, 
    0.6544563, 0.6546437, 0.6541349, 0.6575849, 0.6563354, 0.6596994, 
    0.6587906, 0.6602794, 0.6595398, 0.6594309, 0.6584805, 0.6578887, 
    0.6563928, 0.6551749, 0.6542087, 0.6544334, 0.6554946, 0.6574154, 
    0.6592311, 0.6588335, 0.6601663, 0.6566368, 0.6581175, 0.6575453, 
    0.6590368, 0.6557674, 0.6585523, 0.6550551, 0.6553619, 0.6563106, 
    0.658218, 0.6586395, 0.6590899, 0.6588119, 0.6574641, 0.6572432, 
    0.6562875, 0.6560237, 0.6552951, 0.6546918, 0.655243, 0.6558219, 
    0.6574647, 0.6589443, 0.6605564, 0.6609507, 0.6628332, 0.6613012, 
    0.6638291, 0.6616805, 0.6653984, 0.6587133, 0.6616169, 0.6563537, 
    0.6569212, 0.6579475, 0.6602995, 0.6590298, 0.6605145, 0.6572345, 
    0.6555313, 0.6550902, 0.6542674, 0.655109, 0.6550406, 0.6558457, 
    0.655587, 0.6575192, 0.6564814, 0.6594282, 0.6605027, 0.6635345, 
    0.6653913, 0.6672795, 0.6681129, 0.6683664, 0.6684724,
  0.65618, 0.6580042, 0.6576495, 0.659121, 0.6583046, 0.6592683, 0.6565498, 
    0.6580766, 0.6571018, 0.6563441, 0.6619779, 0.6591867, 0.6648777, 
    0.6630968, 0.667571, 0.6646006, 0.6681701, 0.6674851, 0.6695464, 
    0.6689558, 0.6715935, 0.6698191, 0.6729609, 0.6711696, 0.6714498, 
    0.6697605, 0.6597481, 0.6616304, 0.6596367, 0.659905, 0.6597846, 
    0.6583216, 0.6575845, 0.6560405, 0.6563208, 0.6574547, 0.6600257, 
    0.6591527, 0.6613526, 0.661303, 0.663753, 0.6626482, 0.6667672, 
    0.6655962, 0.6689805, 0.6681293, 0.6689405, 0.6686945, 0.6689437, 
    0.6676953, 0.6682302, 0.6671317, 0.6628551, 0.6641118, 0.6603646, 
    0.6581126, 0.6566167, 0.6555555, 0.6557056, 0.6559916, 0.6574613, 
    0.6588433, 0.6598967, 0.6606014, 0.6612958, 0.6633987, 0.6645115, 
    0.6670042, 0.6665541, 0.6673164, 0.6680446, 0.6692675, 0.6690661, 
    0.669605, 0.6672962, 0.6688306, 0.6662977, 0.6669905, 0.6614853, 
    0.6593882, 0.6584976, 0.6577176, 0.6558209, 0.6571308, 0.6566144, 
    0.6578428, 0.6586235, 0.6582373, 0.6606207, 0.659694, 0.6645774, 
    0.6624736, 0.6679596, 0.6666464, 0.6682744, 0.6674436, 0.6688672, 
    0.667586, 0.6698055, 0.670289, 0.6699586, 0.6712276, 0.667515, 0.6689406, 
    0.6582265, 0.6582895, 0.6585829, 0.6572934, 0.6572145, 0.6560329, 
    0.6570842, 0.657532, 0.6586687, 0.6593412, 0.6599805, 0.6613863, 
    0.6629568, 0.6651533, 0.6667315, 0.6677898, 0.6671408, 0.6677138, 
    0.6670733, 0.6667731, 0.6701078, 0.6682352, 0.6710451, 0.6708895, 
    0.6696178, 0.670907, 0.6583337, 0.6579713, 0.6567134, 0.6576978, 
    0.6559042, 0.6569082, 0.6574856, 0.6597135, 0.660203, 0.660657, 
    0.6615537, 0.6627048, 0.6647244, 0.6664821, 0.6680869, 0.6679693, 
    0.6680107, 0.6683694, 0.6674811, 0.6685151, 0.6686888, 0.6682349, 
    0.6708687, 0.6701161, 0.6708862, 0.6703962, 0.6580891, 0.6586989, 
    0.6583694, 0.6589891, 0.6585525, 0.6604939, 0.6610761, 0.6638005, 
    0.6626821, 0.664462, 0.6628628, 0.6631463, 0.6645204, 0.6629492, 
    0.6663853, 0.6640558, 0.6683832, 0.6660566, 0.6685291, 0.66808, 
    0.6688235, 0.6694897, 0.6703276, 0.6718743, 0.6715161, 0.6728097, 
    0.659608, 0.6603992, 0.6603294, 0.6611574, 0.6617697, 0.6630971, 
    0.6652268, 0.6644258, 0.6658961, 0.6661914, 0.6639575, 0.6653292, 
    0.6609286, 0.6616395, 0.6612161, 0.6596705, 0.6646106, 0.6620749, 
    0.6667577, 0.6653835, 0.6693947, 0.6673997, 0.6713189, 0.6729954, 
    0.6745731, 0.6764179, 0.6608309, 0.6602933, 0.6612558, 0.6625879, 
    0.6638238, 0.6654673, 0.6656355, 0.6659434, 0.6667411, 0.667412, 
    0.666041, 0.6675801, 0.6618047, 0.6648306, 0.6600901, 0.6615174, 
    0.6625093, 0.6620741, 0.6643342, 0.6648671, 0.6670328, 0.6659131, 
    0.6725817, 0.6696305, 0.6778226, 0.6755323, 0.6601055, 0.6608289, 
    0.6633477, 0.6621491, 0.665577, 0.6664211, 0.6671072, 0.6679846, 
    0.6680793, 0.6685991, 0.6677473, 0.6685655, 0.6654708, 0.6668535, 
    0.6630596, 0.6639829, 0.6635581, 0.6630923, 0.6645302, 0.6660626, 
    0.6660951, 0.6665866, 0.6679721, 0.6655909, 0.6729631, 0.6684096, 
    0.661618, 0.6630122, 0.6632111, 0.662671, 0.6663365, 0.6650081, 
    0.6685864, 0.6676191, 0.6692041, 0.6684164, 0.6683006, 0.6672891, 
    0.6666595, 0.6650691, 0.6637753, 0.6627493, 0.6629878, 0.6641148, 
    0.6661563, 0.6680879, 0.6676648, 0.6690836, 0.6653284, 0.6669029, 
    0.6662944, 0.6678811, 0.6644046, 0.6673656, 0.663648, 0.6639738, 
    0.6649818, 0.6670098, 0.6674583, 0.6679375, 0.6676418, 0.6662081, 
    0.6659731, 0.6649572, 0.6646768, 0.6639029, 0.6632622, 0.6638476, 
    0.6644624, 0.6662086, 0.6677827, 0.6694992, 0.6699192, 0.671926, 
    0.6702926, 0.6729885, 0.6706969, 0.6746641, 0.6675369, 0.6706291, 
    0.6650276, 0.6656308, 0.6667221, 0.6692255, 0.6678737, 0.6694545, 
    0.6659639, 0.6641538, 0.6636853, 0.6628117, 0.6637053, 0.6636326, 
    0.6644878, 0.6642129, 0.6662666, 0.6651634, 0.6682978, 0.6694419, 
    0.6726741, 0.6746565, 0.6766747, 0.6775661, 0.6778374, 0.6779508,
  0.6732581, 0.6752667, 0.6748759, 0.6764982, 0.6755978, 0.6766607, 
    0.6736649, 0.6753466, 0.6742727, 0.6734386, 0.6796541, 0.6765706, 
    0.6828659, 0.6808923, 0.6858573, 0.6825587, 0.6865237, 0.6857617, 
    0.6880563, 0.6873984, 0.6903397, 0.6883601, 0.6918676, 0.6898665, 
    0.6901793, 0.6882949, 0.6771902, 0.6792697, 0.6770672, 0.6773634, 
    0.6772304, 0.6756166, 0.6748043, 0.6731046, 0.6734129, 0.6746613, 
    0.6774967, 0.6765332, 0.6789626, 0.6789077, 0.6816191, 0.6803957, 
    0.6849638, 0.6836632, 0.6874259, 0.6864783, 0.6873813, 0.6871074, 
    0.6873849, 0.6859956, 0.6865906, 0.6853688, 0.6806248, 0.6820168, 
    0.6778709, 0.6753863, 0.6737387, 0.6725712, 0.6727362, 0.6730508, 
    0.6746687, 0.6761919, 0.6773542, 0.6781324, 0.6788998, 0.6812266, 
    0.6824598, 0.685227, 0.6847269, 0.6855742, 0.686384, 0.6877455, 
    0.6875212, 0.6881216, 0.6855517, 0.687259, 0.6844422, 0.6852118, 
    0.6791092, 0.676793, 0.6758106, 0.674951, 0.672863, 0.6743045, 0.6737361, 
    0.6750888, 0.6759494, 0.6755237, 0.6781538, 0.6771305, 0.682533, 
    0.6802024, 0.6862895, 0.6848295, 0.6866398, 0.6857156, 0.6872997, 
    0.6858739, 0.688345, 0.688884, 0.6885157, 0.6899312, 0.6857949, 
    0.6873814, 0.6755118, 0.6755812, 0.6759046, 0.6744837, 0.6743968, 
    0.6730962, 0.6742533, 0.6747465, 0.6759993, 0.6767411, 0.6774467, 
    0.6789998, 0.6807373, 0.6831717, 0.6849241, 0.6861006, 0.685379, 
    0.686016, 0.6853039, 0.6849703, 0.6886821, 0.6865962, 0.6897275, 
    0.6895539, 0.6881359, 0.6895735, 0.67563, 0.6752305, 0.673845, 0.6749291, 
    0.6729546, 0.6740595, 0.6746954, 0.677152, 0.6776924, 0.6781939, 
    0.6791849, 0.6804583, 0.682696, 0.6846469, 0.6864312, 0.6863003, 
    0.6863464, 0.6867454, 0.6857573, 0.6869078, 0.687101, 0.6865959, 
    0.6895307, 0.6886913, 0.6895502, 0.6890036, 0.6753603, 0.6760326, 
    0.6756693, 0.6763526, 0.6758712, 0.6780137, 0.6786569, 0.6816719, 
    0.6804333, 0.682405, 0.6806333, 0.6809471, 0.6824697, 0.6807289, 
    0.6845394, 0.6819547, 0.686761, 0.6841744, 0.6869233, 0.6864234, 
    0.6872511, 0.687993, 0.6889271, 0.6906533, 0.6902533, 0.6916985, 
    0.6770356, 0.6779091, 0.677832, 0.6787468, 0.6794238, 0.6808927, 
    0.6832532, 0.6823649, 0.6839962, 0.684324, 0.6818458, 0.6833668, 
    0.678494, 0.6792798, 0.6788117, 0.6771045, 0.6825697, 0.6797614, 
    0.6849531, 0.6834272, 0.6878873, 0.6856667, 0.6900331, 0.6919062, 
    0.6936718, 0.6957403, 0.678386, 0.6777921, 0.6788555, 0.680329, 
    0.6816976, 0.6835202, 0.6837068, 0.6840487, 0.6849347, 0.6856804, 
    0.684157, 0.6858674, 0.6794624, 0.6828138, 0.6775678, 0.6791448, 
    0.680242, 0.6797604, 0.6822634, 0.6828542, 0.6852589, 0.684015, 
    0.6914437, 0.68815, 0.6973178, 0.6947468, 0.6775847, 0.6783838, 
    0.6811702, 0.6798435, 0.6836419, 0.6845791, 0.6853416, 0.6863173, 
    0.6864226, 0.6870012, 0.6860533, 0.6869637, 0.6835241, 0.6850597, 
    0.6808512, 0.6818739, 0.6814032, 0.6808873, 0.6824806, 0.684181, 
    0.6842171, 0.684763, 0.6863034, 0.6836573, 0.6918701, 0.6867902, 
    0.679256, 0.6807986, 0.6810189, 0.6804209, 0.6844851, 0.6830107, 
    0.6869871, 0.6859108, 0.6876749, 0.6867979, 0.6866689, 0.6855438, 
    0.6848441, 0.6830783, 0.6816438, 0.6805076, 0.6807717, 0.6820201, 
    0.684285, 0.6864322, 0.6859615, 0.6875407, 0.683366, 0.6851145, 
    0.6844384, 0.6862022, 0.6823413, 0.6856288, 0.6815028, 0.6818638, 
    0.6829814, 0.6852334, 0.6857319, 0.686265, 0.685936, 0.6843426, 
    0.6840817, 0.6829542, 0.6826432, 0.6817852, 0.6810755, 0.681724, 
    0.6824055, 0.6843432, 0.6860927, 0.6880037, 0.6884718, 0.690711, 
    0.6888881, 0.6918985, 0.689339, 0.6937739, 0.6858193, 0.6892633, 
    0.6830322, 0.6837016, 0.6849136, 0.6876987, 0.6861939, 0.6879539, 
    0.6840714, 0.6820633, 0.6815442, 0.6805767, 0.6815663, 0.6814858, 
    0.6824335, 0.6821289, 0.6844075, 0.6831829, 0.6866658, 0.6879399, 
    0.691547, 0.6937653, 0.6960285, 0.6970295, 0.6973344, 0.6974619,
  0.6968738, 0.6993591, 0.6988748, 0.7008876, 0.6997698, 0.7010895, 
    0.6973764, 0.6994581, 0.698128, 0.6970968, 0.7048212, 0.7009776, 0.70885, 
    0.7063712, 0.7126261, 0.7084634, 0.7134706, 0.7125052, 0.7154173, 
    0.7145808, 0.7183295, 0.7158039, 0.7202864, 0.7177247, 0.7181244, 
    0.7157209, 0.701748, 0.7043408, 0.7015949, 0.7019636, 0.7017981, 
    0.6997929, 0.6987861, 0.6966842, 0.6970651, 0.6986091, 0.7021294, 
    0.7009311, 0.7039573, 0.7038887, 0.707283, 0.7057492, 0.7114957, 
    0.7098542, 0.7146157, 0.713413, 0.7145591, 0.7142112, 0.7145637, 
    0.7128012, 0.7135554, 0.7120079, 0.706036, 0.7077823, 0.7025955, 
    0.6995073, 0.6974676, 0.696026, 0.6962295, 0.6966178, 0.6986181, 
    0.700507, 0.7019521, 0.7029215, 0.7038788, 0.7067904, 0.7083392, 
    0.7118286, 0.7111964, 0.7122678, 0.7132935, 0.7150219, 0.7147369, 
    0.7155003, 0.7122393, 0.7144037, 0.7108368, 0.7118093, 0.7041403, 
    0.701254, 0.7000338, 0.6989679, 0.6963861, 0.6981674, 0.6974643, 
    0.6991386, 0.700206, 0.6996778, 0.702948, 0.7016737, 0.7084311, 
    0.7055072, 0.7131737, 0.7113261, 0.7136178, 0.7124467, 0.7144555, 
    0.7126472, 0.7157847, 0.7164713, 0.716002, 0.7178074, 0.7125472, 
    0.7145593, 0.699663, 0.6997491, 0.7001504, 0.6983892, 0.6982816, 
    0.6966739, 0.698104, 0.6987146, 0.7002679, 0.7011895, 0.7020673, 
    0.7040038, 0.7061771, 0.7092348, 0.7114456, 0.7129343, 0.7120208, 
    0.7128271, 0.7119258, 0.711504, 0.7162139, 0.7135625, 0.7175472, 
    0.7173256, 0.7155185, 0.7173506, 0.6998096, 0.6993142, 0.697599, 
    0.6989408, 0.6964991, 0.6978643, 0.6986512, 0.7017005, 0.7023731, 
    0.7029981, 0.7042349, 0.7058275, 0.7086362, 0.7110954, 0.7133532, 
    0.7131873, 0.7132457, 0.7137519, 0.7124996, 0.7139578, 0.7142031, 
    0.7135621, 0.7172959, 0.7162256, 0.7173209, 0.7166236, 0.6994752, 
    0.7003093, 0.6998584, 0.7007067, 0.7001089, 0.7027735, 0.7035757, 
    0.7073491, 0.7057962, 0.7082702, 0.7060468, 0.7064399, 0.7083516, 
    0.7061665, 0.7109596, 0.7077044, 0.7137715, 0.7104988, 0.7139775, 
    0.7133434, 0.7143937, 0.7153367, 0.7165262, 0.7187305, 0.7182189, 
    0.7200694, 0.7015556, 0.7026431, 0.7025471, 0.7036877, 0.7045333, 
    0.7063718, 0.7093375, 0.7082198, 0.710274, 0.7106877, 0.7075676, 
    0.7094806, 0.7033724, 0.7043534, 0.7037689, 0.7016414, 0.7084773, 
    0.7049553, 0.7114823, 0.7095567, 0.7152022, 0.7123849, 0.7179376, 
    0.7203358, 0.7226056, 0.7252764, 0.7032376, 0.7024974, 0.7038236, 
    0.7056656, 0.7073814, 0.7096739, 0.7099091, 0.7103403, 0.711459, 
    0.7124022, 0.7104769, 0.7126389, 0.7045816, 0.7087843, 0.702218, 
    0.7041848, 0.7055567, 0.7049541, 0.7080922, 0.7088352, 0.7118689, 
    0.7102978, 0.7197427, 0.7155365, 0.7273219, 0.723992, 0.7022391, 
    0.703235, 0.7067196, 0.705058, 0.7098273, 0.7110098, 0.7119735, 0.713209, 
    0.7133424, 0.7140765, 0.7128744, 0.7140288, 0.7096788, 0.711617, 
    0.7063197, 0.7076029, 0.707012, 0.706365, 0.7083652, 0.7105072, 
    0.7105528, 0.7112421, 0.7131913, 0.7098467, 0.7202895, 0.7138087, 
    0.7043236, 0.7062538, 0.70653, 0.7057807, 0.7108911, 0.7090322, 
    0.7140585, 0.7126939, 0.7149321, 0.7138184, 0.7136548, 0.7122293, 
    0.7113444, 0.7091173, 0.7073139, 0.7058893, 0.7062201, 0.7077865, 
    0.7106385, 0.7133546, 0.7127581, 0.7147616, 0.7094796, 0.7116863, 
    0.7108321, 0.7130631, 0.7081901, 0.7123369, 0.707137, 0.7075902, 
    0.7089953, 0.7118366, 0.7124674, 0.7131426, 0.7127258, 0.7107111, 
    0.7103818, 0.7089611, 0.7085698, 0.7074915, 0.7066009, 0.7074146, 
    0.7082708, 0.7107118, 0.7129242, 0.7153502, 0.7159461, 0.7188044, 
    0.7164764, 0.7203259, 0.7170513, 0.7227371, 0.7125781, 0.7169549, 
    0.7090593, 0.7099025, 0.7114323, 0.7149624, 0.7130525, 0.7152869, 
    0.7103689, 0.7078408, 0.7071888, 0.7059758, 0.7072166, 0.7071156, 
    0.7083061, 0.7079232, 0.7107931, 0.709249, 0.7136508, 0.7152691, 
    0.7198752, 0.722726, 0.7256494, 0.7269474, 0.7273434, 0.727509,
  0.7536336, 0.7576361, 0.7568524, 0.7601215, 0.7583021, 0.7604513, 
    0.7544393, 0.7577966, 0.7556476, 0.7539909, 0.7666051, 0.7602684, 
    0.7733833, 0.769196, 0.7798715, 0.7727266, 0.7813413, 0.7796615, 
    0.7847567, 0.7832844, 0.7899396, 0.7854396, 0.7934738, 0.7888559, 
    0.7895718, 0.7852929, 0.7615289, 0.7658064, 0.7612781, 0.7618824, 
    0.7616109, 0.7583396, 0.7567092, 0.7533303, 0.75394, 0.7564232, 
    0.7621546, 0.7601925, 0.7651701, 0.7650564, 0.7707297, 0.7681537, 
    0.7779149, 0.7750956, 0.7833456, 0.7812408, 0.7832464, 0.7826362, 
    0.7832544, 0.7801757, 0.7814893, 0.7788, 0.7686339, 0.7715728, 0.7629209, 
    0.7578763, 0.7545856, 0.752279, 0.7526037, 0.753224, 0.7564378, 
    0.7595009, 0.7618635, 0.763458, 0.7650401, 0.7699003, 0.7725158, 
    0.7784898, 0.7773989, 0.7792498, 0.7810325, 0.78406, 0.7835586, 
    0.7849032, 0.7792005, 0.7829736, 0.7767802, 0.7784564, 0.7654737, 
    0.7607201, 0.7587309, 0.7570029, 0.7528537, 0.7557111, 0.7545804, 
    0.7572792, 0.759011, 0.7581527, 0.7635017, 0.7614071, 0.7726718, 
    0.7677492, 0.7808238, 0.7776224, 0.7815983, 0.7795601, 0.7830645, 
    0.779908, 0.7854057, 0.7866222, 0.7857901, 0.7890038, 0.7797344, 
    0.7832466, 0.7581288, 0.7582685, 0.7589206, 0.7560684, 0.755895, 
    0.7533137, 0.755609, 0.7565935, 0.7591116, 0.7606146, 0.7620526, 
    0.7652472, 0.7688702, 0.7740384, 0.7778285, 0.780407, 0.7788221, 
    0.7802207, 0.7786579, 0.7779292, 0.7861657, 0.7815017, 0.7885385, 
    0.7881429, 0.7849354, 0.7881874, 0.7583667, 0.7575634, 0.7547967, 
    0.756959, 0.7530343, 0.7552231, 0.7564912, 0.761451, 0.7625551, 
    0.7635843, 0.7656305, 0.7682848, 0.7730199, 0.777225, 0.7811366, 
    0.7808475, 0.7809492, 0.7818323, 0.7796518, 0.7821925, 0.782622, 
    0.7815009, 0.78809, 0.7861864, 0.7881345, 0.7868928, 0.7578242, 
    0.7591789, 0.7584459, 0.7598264, 0.7588531, 0.7632141, 0.7645382, 
    0.7708414, 0.7682323, 0.7723989, 0.7686518, 0.7693112, 0.7725368, 
    0.7688527, 0.7769913, 0.7714411, 0.7818667, 0.7761997, 0.782227, 
    0.7811195, 0.7829561, 0.7846147, 0.7867197, 0.7906605, 0.7897412, 
    0.7930799, 0.7612137, 0.7629993, 0.7628412, 0.7647237, 0.7661263, 
    0.7691969, 0.7742134, 0.7723134, 0.7758142, 0.7765239, 0.77121, 
    0.7744575, 0.7642021, 0.7658274, 0.7648581, 0.7613541, 0.7727501, 
    0.7668286, 0.7778918, 0.7745873, 0.7843775, 0.7794529, 0.789237, 
    0.7935637, 0.7977186, 0.8026853, 0.7639796, 0.7627594, 0.7649486, 
    0.7680139, 0.7708958, 0.7747874, 0.7751894, 0.7759277, 0.7778517, 
    0.7794829, 0.776162, 0.7798938, 0.7662066, 0.7732716, 0.7623001, 
    0.7655474, 0.7678319, 0.7668266, 0.7720972, 0.7733582, 0.7785594, 
    0.7758549, 0.7924877, 0.7849671, 0.8065489, 0.8002861, 0.7623348, 
    0.7639752, 0.7697812, 0.7669997, 0.7750496, 0.7770777, 0.7787403, 
    0.7808852, 0.7811177, 0.7824002, 0.7803028, 0.7823168, 0.7747958, 
    0.7781242, 0.7691095, 0.7712697, 0.7702731, 0.7691855, 0.7725599, 
    0.7762139, 0.7762922, 0.7774776, 0.7808545, 0.7750828, 0.7934795, 
    0.7819318, 0.7657779, 0.768999, 0.7694625, 0.7682065, 0.7768735, 
    0.7736932, 0.7823688, 0.7799891, 0.783902, 0.7819487, 0.7816628, 
    0.7791833, 0.7776541, 0.7738381, 0.7707819, 0.7683882, 0.7689424, 
    0.77158, 0.7764394, 0.7811391, 0.7801008, 0.7836021, 0.7744558, 
    0.7782439, 0.776772, 0.7806311, 0.7722632, 0.7793697, 0.7704836, 
    0.7712482, 0.7736306, 0.7785036, 0.779596, 0.7807695, 0.7800446, 
    0.7765641, 0.775999, 0.7735722, 0.7729072, 0.7710815, 0.7695817, 
    0.7709517, 0.7723999, 0.7765653, 0.7803896, 0.7846385, 0.7856911, 
    0.7907935, 0.7866313, 0.7935457, 0.7876538, 0.797961, 0.779788, 0.787482, 
    0.7737394, 0.7751782, 0.7778056, 0.7839553, 0.7806128, 0.7845268, 
    0.7759768, 0.7716718, 0.7705711, 0.7685331, 0.7706179, 0.7704476, 
    0.7724597, 0.7718111, 0.776705, 0.7740625, 0.7816558, 0.7844955, 
    0.7927276, 0.7979407, 0.8033861, 0.8058377, 0.8065898, 0.806905,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 XSMRPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 XSMRPOOL_RECOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZBOT =
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5 ;

 ZWT =
  8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882 ;

 ZWT_CH4_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZWT_PERCH =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 o2_decomp_depth_unsat =
  3.698585e-11, 3.714113e-11, 3.711087e-11, 3.723616e-11, 3.716662e-11, 
    3.72486e-11, 3.701715e-11, 3.714701e-11, 3.706406e-11, 3.699952e-11, 
    3.747913e-11, 3.724145e-11, 3.77266e-11, 3.757467e-11, 3.795644e-11, 
    3.770282e-11, 3.800759e-11, 3.794908e-11, 3.81252e-11, 3.807466e-11, 
    3.829991e-11, 3.814839e-11, 3.841682e-11, 3.826368e-11, 3.828755e-11, 
    3.814319e-11, 3.72896e-11, 3.74498e-11, 3.728002e-11, 3.730286e-11, 
    3.729258e-11, 3.716787e-11, 3.710503e-11, 3.697367e-11, 3.699746e-11, 
    3.709393e-11, 3.731285e-11, 3.723847e-11, 3.74259e-11, 3.742168e-11, 
    3.763049e-11, 3.753628e-11, 3.788773e-11, 3.778772e-11, 3.807673e-11, 
    3.800393e-11, 3.807322e-11, 3.805215e-11, 3.807338e-11, 3.796673e-11, 
    3.801233e-11, 3.791853e-11, 3.755438e-11, 3.76615e-11, 3.734196e-11, 
    3.714994e-11, 3.702266e-11, 3.69324e-11, 3.694508e-11, 3.69694e-11, 
    3.709441e-11, 3.721208e-11, 3.730181e-11, 3.73618e-11, 3.742095e-11, 
    3.760009e-11, 3.769507e-11, 3.790783e-11, 3.786944e-11, 3.793443e-11, 
    3.799665e-11, 3.810106e-11, 3.808385e-11, 3.812981e-11, 3.793254e-11, 
    3.806358e-11, 3.784723e-11, 3.790636e-11, 3.743722e-11, 3.72587e-11, 
    3.71827e-11, 3.711632e-11, 3.695485e-11, 3.70663e-11, 3.702231e-11, 
    3.712685e-11, 3.719331e-11, 3.716038e-11, 3.73634e-11, 3.728437e-11, 
    3.770063e-11, 3.752121e-11, 3.798944e-11, 3.787723e-11, 3.801623e-11, 
    3.794528e-11, 3.806677e-11, 3.795736e-11, 3.814688e-11, 3.818817e-11, 
    3.815987e-11, 3.826837e-11, 3.795104e-11, 3.80728e-11, 3.715968e-11, 
    3.716505e-11, 3.718999e-11, 3.708008e-11, 3.707336e-11, 3.697276e-11, 
    3.706218e-11, 3.710029e-11, 3.719708e-11, 3.725428e-11, 3.730869e-11, 
    3.742852e-11, 3.756232e-11, 3.774968e-11, 3.788445e-11, 3.797478e-11, 
    3.791935e-11, 3.796821e-11, 3.79135e-11, 3.788781e-11, 3.817257e-11, 
    3.801259e-11, 3.825264e-11, 3.823936e-11, 3.813059e-11, 3.824075e-11, 
    3.716873e-11, 3.713783e-11, 3.703069e-11, 3.711446e-11, 3.696174e-11, 
    3.704716e-11, 3.709622e-11, 3.728591e-11, 3.732763e-11, 3.736631e-11, 
    3.744272e-11, 3.754079e-11, 3.771305e-11, 3.786303e-11, 3.800012e-11, 
    3.799001e-11, 3.799353e-11, 3.802409e-11, 3.794821e-11, 3.803647e-11, 
    3.805122e-11, 3.801249e-11, 3.823747e-11, 3.817316e-11, 3.823892e-11, 
    3.819698e-11, 3.714782e-11, 3.719967e-11, 3.717156e-11, 3.722432e-11, 
    3.718705e-11, 3.735241e-11, 3.740195e-11, 3.763424e-11, 3.753885e-11, 
    3.769067e-11, 3.75542e-11, 3.757836e-11, 3.76954e-11, 3.756149e-11, 
    3.785459e-11, 3.765567e-11, 3.802523e-11, 3.782633e-11, 3.803761e-11, 
    3.79992e-11, 3.806267e-11, 3.811957e-11, 3.819111e-11, 3.832328e-11, 
    3.829259e-11, 3.840321e-11, 3.727707e-11, 3.734438e-11, 3.733847e-11, 
    3.740897e-11, 3.74611e-11, 3.757434e-11, 3.775597e-11, 3.768758e-11, 
    3.781303e-11, 3.783822e-11, 3.76475e-11, 3.77645e-11, 3.738911e-11, 
    3.744959e-11, 3.741355e-11, 3.728175e-11, 3.770293e-11, 3.748657e-11, 
    3.788619e-11, 3.776883e-11, 3.811133e-11, 3.794086e-11, 3.827571e-11, 
    3.841895e-11, 3.855398e-11, 3.871166e-11, 3.738116e-11, 3.73353e-11, 
    3.741729e-11, 3.753079e-11, 3.763619e-11, 3.777645e-11, 3.779078e-11, 
    3.781699e-11, 3.788507e-11, 3.794236e-11, 3.782516e-11, 3.795661e-11, 
    3.74635e-11, 3.772173e-11, 3.731744e-11, 3.743902e-11, 3.752356e-11, 
    3.748648e-11, 3.767927e-11, 3.772466e-11, 3.790944e-11, 3.78139e-11, 
    3.838343e-11, 3.813123e-11, 3.883189e-11, 3.863582e-11, 3.731926e-11, 
    3.738086e-11, 3.759551e-11, 3.749333e-11, 3.778572e-11, 3.785777e-11, 
    3.79163e-11, 3.79912e-11, 3.799923e-11, 3.804363e-11, 3.79708e-11, 
    3.80407e-11, 3.777632e-11, 3.78944e-11, 3.757057e-11, 3.764924e-11, 
    3.761302e-11, 3.757322e-11, 3.769583e-11, 3.782655e-11, 3.782936e-11, 
    3.787121e-11, 3.798924e-11, 3.778618e-11, 3.841573e-11, 3.802651e-11, 
    3.744807e-11, 3.756679e-11, 3.758379e-11, 3.753776e-11, 3.785043e-11, 
    3.773705e-11, 3.804256e-11, 3.795988e-11, 3.809522e-11, 3.802794e-11, 
    3.801795e-11, 3.793157e-11, 3.78777e-11, 3.774192e-11, 3.763143e-11, 
    3.754397e-11, 3.756423e-11, 3.766033e-11, 3.783444e-11, 3.799944e-11, 
    3.796323e-11, 3.808443e-11, 3.776368e-11, 3.789807e-11, 3.784601e-11, 
    3.798157e-11, 3.768558e-11, 3.793811e-11, 3.762102e-11, 3.764875e-11, 
    3.773468e-11, 3.790774e-11, 3.794606e-11, 3.798697e-11, 3.796166e-11, 
    3.783918e-11, 3.78191e-11, 3.773235e-11, 3.770834e-11, 3.764235e-11, 
    3.758761e-11, 3.763753e-11, 3.768987e-11, 3.783894e-11, 3.797328e-11, 
    3.811988e-11, 3.815579e-11, 3.832706e-11, 3.818746e-11, 3.841768e-11, 
    3.822172e-11, 3.856103e-11, 3.795274e-11, 3.821692e-11, 3.773863e-11, 
    3.779005e-11, 3.788312e-11, 3.809685e-11, 3.798142e-11, 3.81164e-11, 
    3.781829e-11, 3.766368e-11, 3.762374e-11, 3.754922e-11, 3.762537e-11, 
    3.761918e-11, 3.76921e-11, 3.766859e-11, 3.784378e-11, 3.774964e-11, 
    3.801715e-11, 3.811488e-11, 3.839113e-11, 3.856058e-11, 3.873336e-11, 
    3.880958e-11, 3.88328e-11, 3.884246e-11,
  2.482071e-11, 2.495144e-11, 2.492602e-11, 2.503156e-11, 2.497302e-11, 
    2.504213e-11, 2.484722e-11, 2.495662e-11, 2.488678e-11, 2.48325e-11, 
    2.523665e-11, 2.503628e-11, 2.544547e-11, 2.53173e-11, 2.563967e-11, 
    2.542549e-11, 2.568292e-11, 2.563353e-11, 2.578238e-11, 2.573972e-11, 
    2.593025e-11, 2.580208e-11, 2.602924e-11, 2.589966e-11, 2.59199e-11, 
    2.579785e-11, 2.507661e-11, 2.521167e-11, 2.50686e-11, 2.508785e-11, 
    2.507922e-11, 2.497421e-11, 2.492131e-11, 2.481076e-11, 2.483082e-11, 
    2.491204e-11, 2.509651e-11, 2.503388e-11, 2.51919e-11, 2.518833e-11, 
    2.536454e-11, 2.528504e-11, 2.558174e-11, 2.549733e-11, 2.57415e-11, 
    2.568003e-11, 2.57386e-11, 2.572085e-11, 2.573884e-11, 2.56487e-11, 
    2.56873e-11, 2.560805e-11, 2.529991e-11, 2.539035e-11, 2.512087e-11, 
    2.495914e-11, 2.485201e-11, 2.477602e-11, 2.478676e-11, 2.480723e-11, 
    2.491252e-11, 2.501167e-11, 2.508729e-11, 2.513791e-11, 2.518781e-11, 
    2.533891e-11, 2.54191e-11, 2.55988e-11, 2.556638e-11, 2.562133e-11, 
    2.567392e-11, 2.576221e-11, 2.574768e-11, 2.578659e-11, 2.561991e-11, 
    2.573064e-11, 2.554792e-11, 2.559785e-11, 2.520122e-11, 2.505078e-11, 
    2.498677e-11, 2.49309e-11, 2.479502e-11, 2.488883e-11, 2.485183e-11, 
    2.493991e-11, 2.49959e-11, 2.496821e-11, 2.513929e-11, 2.507273e-11, 
    2.542385e-11, 2.527245e-11, 2.566778e-11, 2.557304e-11, 2.569051e-11, 
    2.563056e-11, 2.57333e-11, 2.564083e-11, 2.580109e-11, 2.5836e-11, 
    2.581214e-11, 2.590389e-11, 2.56357e-11, 2.573859e-11, 2.496742e-11, 
    2.497194e-11, 2.499299e-11, 2.490048e-11, 2.489483e-11, 2.48102e-11, 
    2.488552e-11, 2.49176e-11, 2.499916e-11, 2.50474e-11, 2.50933e-11, 
    2.51943e-11, 2.53072e-11, 2.546536e-11, 2.557918e-11, 2.565554e-11, 
    2.560872e-11, 2.565005e-11, 2.560384e-11, 2.55822e-11, 2.58229e-11, 
    2.568766e-11, 2.589069e-11, 2.587945e-11, 2.578751e-11, 2.588071e-11, 
    2.497511e-11, 2.494913e-11, 2.485893e-11, 2.492951e-11, 2.480099e-11, 
    2.487289e-11, 2.491424e-11, 2.507409e-11, 2.510929e-11, 2.514189e-11, 
    2.520634e-11, 2.528911e-11, 2.543448e-11, 2.556116e-11, 2.567698e-11, 
    2.56685e-11, 2.567148e-11, 2.569736e-11, 2.563326e-11, 2.570789e-11, 
    2.57204e-11, 2.568766e-11, 2.587794e-11, 2.582354e-11, 2.587921e-11, 
    2.584379e-11, 2.495758e-11, 2.500131e-11, 2.497767e-11, 2.502212e-11, 
    2.499079e-11, 2.513012e-11, 2.517194e-11, 2.536791e-11, 2.528747e-11, 
    2.541556e-11, 2.530049e-11, 2.532086e-11, 2.541968e-11, 2.530672e-11, 
    2.555414e-11, 2.538626e-11, 2.569836e-11, 2.55304e-11, 2.57089e-11, 
    2.567648e-11, 2.573017e-11, 2.577826e-11, 2.583883e-11, 2.595062e-11, 
    2.592473e-11, 2.601833e-11, 2.506656e-11, 2.512334e-11, 2.511837e-11, 
    2.517785e-11, 2.522186e-11, 2.531735e-11, 2.547068e-11, 2.541301e-11, 
    2.551895e-11, 2.554022e-11, 2.537929e-11, 2.547804e-11, 2.516139e-11, 
    2.521244e-11, 2.518206e-11, 2.507102e-11, 2.542625e-11, 2.524375e-11, 
    2.558105e-11, 2.548199e-11, 2.57714e-11, 2.562733e-11, 2.591047e-11, 
    2.603168e-11, 2.614604e-11, 2.627966e-11, 2.515438e-11, 2.511578e-11, 
    2.518494e-11, 2.528065e-11, 2.536964e-11, 2.548802e-11, 2.550016e-11, 
    2.552235e-11, 2.557989e-11, 2.562827e-11, 2.552934e-11, 2.564041e-11, 
    2.522422e-11, 2.544212e-11, 2.510116e-11, 2.520365e-11, 2.527502e-11, 
    2.524374e-11, 2.540642e-11, 2.54448e-11, 2.560088e-11, 2.552018e-11, 
    2.600172e-11, 2.578838e-11, 2.638163e-11, 2.621548e-11, 2.510229e-11, 
    2.515426e-11, 2.533534e-11, 2.524914e-11, 2.549595e-11, 2.555678e-11, 
    2.560629e-11, 2.566957e-11, 2.567643e-11, 2.571394e-11, 2.565247e-11, 
    2.571152e-11, 2.548827e-11, 2.558798e-11, 2.531467e-11, 2.53811e-11, 
    2.535054e-11, 2.531701e-11, 2.542053e-11, 2.553088e-11, 2.553329e-11, 
    2.55687e-11, 2.566845e-11, 2.549695e-11, 2.60292e-11, 2.570007e-11, 
    2.521097e-11, 2.531116e-11, 2.532554e-11, 2.52867e-11, 2.555068e-11, 
    2.545494e-11, 2.571304e-11, 2.564322e-11, 2.575765e-11, 2.570077e-11, 
    2.56924e-11, 2.561941e-11, 2.557398e-11, 2.545932e-11, 2.536614e-11, 
    2.529234e-11, 2.53095e-11, 2.539058e-11, 2.553765e-11, 2.567702e-11, 
    2.564647e-11, 2.574895e-11, 2.547803e-11, 2.559151e-11, 2.554762e-11, 
    2.566212e-11, 2.541146e-11, 2.562472e-11, 2.535701e-11, 2.538046e-11, 
    2.545304e-11, 2.559918e-11, 2.563162e-11, 2.566617e-11, 2.564486e-11, 
    2.55414e-11, 2.552448e-11, 2.545129e-11, 2.543106e-11, 2.537536e-11, 
    2.532924e-11, 2.537136e-11, 2.541561e-11, 2.554146e-11, 2.565499e-11, 
    2.577894e-11, 2.580931e-11, 2.595425e-11, 2.583618e-11, 2.603102e-11, 
    2.586524e-11, 2.615245e-11, 2.563716e-11, 2.586047e-11, 2.545636e-11, 
    2.549983e-11, 2.557844e-11, 2.57591e-11, 2.566158e-11, 2.577567e-11, 
    2.552382e-11, 2.539336e-11, 2.535969e-11, 2.529681e-11, 2.536113e-11, 
    2.53559e-11, 2.541748e-11, 2.539769e-11, 2.554564e-11, 2.546614e-11, 
    2.569218e-11, 2.577478e-11, 2.600849e-11, 2.615201e-11, 2.629838e-11, 
    2.636304e-11, 2.638273e-11, 2.639096e-11,
  2.659881e-11, 2.674073e-11, 2.671313e-11, 2.682772e-11, 2.676415e-11, 
    2.68392e-11, 2.662758e-11, 2.674635e-11, 2.667052e-11, 2.66116e-11, 
    2.70505e-11, 2.683284e-11, 2.727736e-11, 2.713808e-11, 2.748846e-11, 
    2.725565e-11, 2.753549e-11, 2.748178e-11, 2.764364e-11, 2.759724e-11, 
    2.780451e-11, 2.766506e-11, 2.791221e-11, 2.777121e-11, 2.779323e-11, 
    2.766046e-11, 2.687663e-11, 2.702335e-11, 2.686794e-11, 2.688884e-11, 
    2.687947e-11, 2.676545e-11, 2.670802e-11, 2.6588e-11, 2.660979e-11, 
    2.669795e-11, 2.689825e-11, 2.683023e-11, 2.700184e-11, 2.699796e-11, 
    2.71894e-11, 2.710303e-11, 2.742548e-11, 2.733372e-11, 2.759917e-11, 
    2.753233e-11, 2.759603e-11, 2.757671e-11, 2.759628e-11, 2.749827e-11, 
    2.754024e-11, 2.745407e-11, 2.711919e-11, 2.721746e-11, 2.69247e-11, 
    2.67491e-11, 2.663278e-11, 2.655031e-11, 2.656196e-11, 2.658417e-11, 
    2.669847e-11, 2.680611e-11, 2.688823e-11, 2.69432e-11, 2.69974e-11, 
    2.716159e-11, 2.72487e-11, 2.744402e-11, 2.740877e-11, 2.746852e-11, 
    2.752569e-11, 2.76217e-11, 2.76059e-11, 2.764822e-11, 2.746697e-11, 
    2.758737e-11, 2.73887e-11, 2.744298e-11, 2.701201e-11, 2.684858e-11, 
    2.67791e-11, 2.671843e-11, 2.657092e-11, 2.667275e-11, 2.663259e-11, 
    2.672819e-11, 2.678899e-11, 2.675892e-11, 2.69447e-11, 2.687242e-11, 
    2.725387e-11, 2.708935e-11, 2.751902e-11, 2.741601e-11, 2.754373e-11, 
    2.747854e-11, 2.759026e-11, 2.748971e-11, 2.766398e-11, 2.770196e-11, 
    2.7676e-11, 2.77758e-11, 2.748413e-11, 2.759601e-11, 2.675807e-11, 
    2.676297e-11, 2.678583e-11, 2.668541e-11, 2.667927e-11, 2.65874e-11, 
    2.666915e-11, 2.670398e-11, 2.679252e-11, 2.684491e-11, 2.689475e-11, 
    2.700445e-11, 2.712711e-11, 2.729897e-11, 2.742268e-11, 2.75057e-11, 
    2.745479e-11, 2.749973e-11, 2.744949e-11, 2.742596e-11, 2.768772e-11, 
    2.754063e-11, 2.776144e-11, 2.774921e-11, 2.764922e-11, 2.775059e-11, 
    2.676642e-11, 2.673821e-11, 2.66403e-11, 2.671691e-11, 2.65774e-11, 
    2.665545e-11, 2.670035e-11, 2.68739e-11, 2.691211e-11, 2.694752e-11, 
    2.701753e-11, 2.710744e-11, 2.726541e-11, 2.74031e-11, 2.752902e-11, 
    2.751979e-11, 2.752304e-11, 2.755117e-11, 2.748148e-11, 2.756262e-11, 
    2.757624e-11, 2.754063e-11, 2.774758e-11, 2.768841e-11, 2.774895e-11, 
    2.771043e-11, 2.674738e-11, 2.679486e-11, 2.67692e-11, 2.681746e-11, 
    2.678345e-11, 2.693475e-11, 2.698018e-11, 2.719307e-11, 2.710567e-11, 
    2.724486e-11, 2.711981e-11, 2.714194e-11, 2.724934e-11, 2.712657e-11, 
    2.739548e-11, 2.721303e-11, 2.755227e-11, 2.736968e-11, 2.756372e-11, 
    2.752847e-11, 2.758685e-11, 2.763916e-11, 2.770503e-11, 2.782666e-11, 
    2.779848e-11, 2.790032e-11, 2.686572e-11, 2.692739e-11, 2.692198e-11, 
    2.698658e-11, 2.703439e-11, 2.713813e-11, 2.730475e-11, 2.724207e-11, 
    2.735721e-11, 2.738034e-11, 2.720543e-11, 2.731275e-11, 2.696871e-11, 
    2.702417e-11, 2.699116e-11, 2.687057e-11, 2.725647e-11, 2.705819e-11, 
    2.742472e-11, 2.731704e-11, 2.763169e-11, 2.747504e-11, 2.778297e-11, 
    2.791487e-11, 2.803931e-11, 2.81848e-11, 2.696109e-11, 2.691916e-11, 
    2.699428e-11, 2.709827e-11, 2.719494e-11, 2.73236e-11, 2.733679e-11, 
    2.736091e-11, 2.742345e-11, 2.747605e-11, 2.736851e-11, 2.748925e-11, 
    2.703699e-11, 2.727371e-11, 2.69033e-11, 2.701463e-11, 2.709214e-11, 
    2.705816e-11, 2.723491e-11, 2.727661e-11, 2.744628e-11, 2.735855e-11, 
    2.788227e-11, 2.765017e-11, 2.829582e-11, 2.811491e-11, 2.690451e-11, 
    2.696096e-11, 2.715769e-11, 2.706403e-11, 2.733221e-11, 2.739834e-11, 
    2.745216e-11, 2.752096e-11, 2.752841e-11, 2.756921e-11, 2.750236e-11, 
    2.756658e-11, 2.732387e-11, 2.743225e-11, 2.713521e-11, 2.720739e-11, 
    2.717419e-11, 2.713776e-11, 2.725024e-11, 2.737019e-11, 2.73728e-11, 
    2.74113e-11, 2.751979e-11, 2.73333e-11, 2.79122e-11, 2.755416e-11, 
    2.702256e-11, 2.713142e-11, 2.714703e-11, 2.710482e-11, 2.73917e-11, 
    2.728764e-11, 2.756822e-11, 2.749231e-11, 2.761674e-11, 2.755488e-11, 
    2.754578e-11, 2.746642e-11, 2.741703e-11, 2.72924e-11, 2.719114e-11, 
    2.711095e-11, 2.71296e-11, 2.721771e-11, 2.737755e-11, 2.752907e-11, 
    2.749585e-11, 2.760727e-11, 2.731274e-11, 2.74361e-11, 2.738838e-11, 
    2.751286e-11, 2.724039e-11, 2.747223e-11, 2.718122e-11, 2.72067e-11, 
    2.728558e-11, 2.744444e-11, 2.747969e-11, 2.751727e-11, 2.749409e-11, 
    2.738162e-11, 2.736322e-11, 2.728367e-11, 2.72617e-11, 2.720116e-11, 
    2.715105e-11, 2.719682e-11, 2.724491e-11, 2.738168e-11, 2.750511e-11, 
    2.763989e-11, 2.767293e-11, 2.783063e-11, 2.770218e-11, 2.791419e-11, 
    2.773382e-11, 2.804632e-11, 2.748575e-11, 2.77286e-11, 2.728918e-11, 
    2.733642e-11, 2.74219e-11, 2.761833e-11, 2.751227e-11, 2.763635e-11, 
    2.736251e-11, 2.722073e-11, 2.718413e-11, 2.711581e-11, 2.718569e-11, 
    2.718001e-11, 2.724693e-11, 2.722542e-11, 2.738623e-11, 2.729981e-11, 
    2.754554e-11, 2.763538e-11, 2.788963e-11, 2.804582e-11, 2.820516e-11, 
    2.827557e-11, 2.829702e-11, 2.830598e-11,
  2.832771e-11, 2.848203e-11, 2.845201e-11, 2.857668e-11, 2.850751e-11, 
    2.858917e-11, 2.835898e-11, 2.848816e-11, 2.840567e-11, 2.83416e-11, 
    2.881922e-11, 2.858225e-11, 2.906635e-11, 2.891457e-11, 2.929652e-11, 
    2.90427e-11, 2.934782e-11, 2.928921e-11, 2.946581e-11, 2.941517e-11, 
    2.964147e-11, 2.948919e-11, 2.97591e-11, 2.960509e-11, 2.962915e-11, 
    2.948417e-11, 2.86299e-11, 2.878967e-11, 2.862044e-11, 2.86432e-11, 
    2.863298e-11, 2.850892e-11, 2.844647e-11, 2.831594e-11, 2.833962e-11, 
    2.843551e-11, 2.865343e-11, 2.85794e-11, 2.876618e-11, 2.876196e-11, 
    2.897048e-11, 2.887639e-11, 2.92278e-11, 2.912775e-11, 2.941728e-11, 
    2.934436e-11, 2.941385e-11, 2.939278e-11, 2.941413e-11, 2.93072e-11, 
    2.935299e-11, 2.925898e-11, 2.889399e-11, 2.900105e-11, 2.868221e-11, 
    2.849117e-11, 2.836463e-11, 2.827497e-11, 2.828763e-11, 2.831179e-11, 
    2.843608e-11, 2.855316e-11, 2.864251e-11, 2.870234e-11, 2.876136e-11, 
    2.894021e-11, 2.903512e-11, 2.924804e-11, 2.920959e-11, 2.927476e-11, 
    2.933711e-11, 2.944187e-11, 2.942462e-11, 2.947081e-11, 2.927306e-11, 
    2.940442e-11, 2.918769e-11, 2.92469e-11, 2.877732e-11, 2.859937e-11, 
    2.852379e-11, 2.845778e-11, 2.829738e-11, 2.84081e-11, 2.836443e-11, 
    2.846839e-11, 2.853452e-11, 2.850181e-11, 2.870398e-11, 2.862531e-11, 
    2.904074e-11, 2.88615e-11, 2.932983e-11, 2.921748e-11, 2.935679e-11, 
    2.928567e-11, 2.940756e-11, 2.929786e-11, 2.948802e-11, 2.952949e-11, 
    2.950114e-11, 2.96101e-11, 2.929178e-11, 2.941385e-11, 2.850089e-11, 
    2.850623e-11, 2.853109e-11, 2.842187e-11, 2.841519e-11, 2.831529e-11, 
    2.840418e-11, 2.844207e-11, 2.853837e-11, 2.859537e-11, 2.864962e-11, 
    2.876903e-11, 2.890263e-11, 2.90899e-11, 2.922476e-11, 2.93153e-11, 
    2.925977e-11, 2.930879e-11, 2.9254e-11, 2.922833e-11, 2.951394e-11, 
    2.935342e-11, 2.959442e-11, 2.958107e-11, 2.947191e-11, 2.958257e-11, 
    2.850997e-11, 2.847928e-11, 2.837281e-11, 2.845612e-11, 2.830442e-11, 
    2.838928e-11, 2.843812e-11, 2.862693e-11, 2.866851e-11, 2.870706e-11, 
    2.878327e-11, 2.888119e-11, 2.905331e-11, 2.920341e-11, 2.934074e-11, 
    2.933067e-11, 2.933422e-11, 2.936492e-11, 2.928888e-11, 2.937741e-11, 
    2.939227e-11, 2.935341e-11, 2.957928e-11, 2.951468e-11, 2.958078e-11, 
    2.953872e-11, 2.848926e-11, 2.854092e-11, 2.8513e-11, 2.856551e-11, 
    2.85285e-11, 2.869317e-11, 2.874262e-11, 2.89745e-11, 2.887926e-11, 
    2.903091e-11, 2.889466e-11, 2.891878e-11, 2.903583e-11, 2.890202e-11, 
    2.919511e-11, 2.899624e-11, 2.936611e-11, 2.9167e-11, 2.93786e-11, 
    2.934014e-11, 2.940384e-11, 2.946092e-11, 2.953282e-11, 2.966565e-11, 
    2.963487e-11, 2.974611e-11, 2.861801e-11, 2.868514e-11, 2.867925e-11, 
    2.874958e-11, 2.880163e-11, 2.891462e-11, 2.909619e-11, 2.902786e-11, 
    2.915337e-11, 2.917859e-11, 2.898794e-11, 2.910492e-11, 2.873012e-11, 
    2.879052e-11, 2.875457e-11, 2.86233e-11, 2.904357e-11, 2.882756e-11, 
    2.922699e-11, 2.910958e-11, 2.945278e-11, 2.928188e-11, 2.961793e-11, 
    2.976203e-11, 2.9898e-11, 3.005712e-11, 2.872183e-11, 2.867618e-11, 
    2.875795e-11, 2.887121e-11, 2.897652e-11, 2.911673e-11, 2.91311e-11, 
    2.91574e-11, 2.922559e-11, 2.928296e-11, 2.91657e-11, 2.929735e-11, 
    2.880451e-11, 2.906236e-11, 2.865892e-11, 2.878013e-11, 2.886454e-11, 
    2.882752e-11, 2.902006e-11, 2.906551e-11, 2.92505e-11, 2.915482e-11, 
    2.972643e-11, 2.947297e-11, 3.017855e-11, 2.998068e-11, 2.866024e-11, 
    2.872168e-11, 2.893593e-11, 2.883391e-11, 2.912611e-11, 2.919821e-11, 
    2.92569e-11, 2.933196e-11, 2.934008e-11, 2.93846e-11, 2.931166e-11, 
    2.938172e-11, 2.911703e-11, 2.923519e-11, 2.891143e-11, 2.899008e-11, 
    2.895389e-11, 2.891421e-11, 2.903676e-11, 2.916754e-11, 2.917037e-11, 
    2.921235e-11, 2.933075e-11, 2.91273e-11, 2.975916e-11, 2.936824e-11, 
    2.878874e-11, 2.890733e-11, 2.892431e-11, 2.887834e-11, 2.919098e-11, 
    2.907754e-11, 2.938351e-11, 2.930069e-11, 2.943645e-11, 2.936896e-11, 
    2.935903e-11, 2.927246e-11, 2.92186e-11, 2.908273e-11, 2.897237e-11, 
    2.888501e-11, 2.890532e-11, 2.900132e-11, 2.917556e-11, 2.93408e-11, 
    2.930457e-11, 2.942612e-11, 2.910489e-11, 2.92394e-11, 2.918737e-11, 
    2.932311e-11, 2.902604e-11, 2.927885e-11, 2.896155e-11, 2.898932e-11, 
    2.907529e-11, 2.924851e-11, 2.928693e-11, 2.932793e-11, 2.930263e-11, 
    2.917999e-11, 2.915993e-11, 2.90732e-11, 2.904926e-11, 2.898328e-11, 
    2.892868e-11, 2.897856e-11, 2.903097e-11, 2.918005e-11, 2.931467e-11, 
    2.946173e-11, 2.949778e-11, 2.967002e-11, 2.952975e-11, 2.976134e-11, 
    2.956435e-11, 2.990572e-11, 2.929358e-11, 2.95586e-11, 2.907921e-11, 
    2.91307e-11, 2.922392e-11, 2.943822e-11, 2.932248e-11, 2.945787e-11, 
    2.915914e-11, 2.900463e-11, 2.896473e-11, 2.889031e-11, 2.896643e-11, 
    2.896024e-11, 2.903315e-11, 2.900971e-11, 2.918501e-11, 2.90908e-11, 
    2.935878e-11, 2.945681e-11, 2.973443e-11, 2.990514e-11, 3.007936e-11, 
    3.015639e-11, 3.017985e-11, 3.018966e-11,
  2.872595e-11, 2.888845e-11, 2.885682e-11, 2.898819e-11, 2.891528e-11, 
    2.900135e-11, 2.875886e-11, 2.889491e-11, 2.880802e-11, 2.874056e-11, 
    2.924409e-11, 2.899406e-11, 2.950513e-11, 2.934471e-11, 2.974865e-11, 
    2.948013e-11, 2.980297e-11, 2.97409e-11, 2.992797e-11, 2.987431e-11, 
    3.011432e-11, 2.995276e-11, 3.023918e-11, 3.00757e-11, 3.010123e-11, 
    2.994744e-11, 2.904428e-11, 2.921289e-11, 2.903431e-11, 2.905831e-11, 
    2.904754e-11, 2.891678e-11, 2.885101e-11, 2.871356e-11, 2.873848e-11, 
    2.883945e-11, 2.906911e-11, 2.899104e-11, 2.918803e-11, 2.918358e-11, 
    2.940377e-11, 2.930437e-11, 2.967589e-11, 2.957003e-11, 2.987655e-11, 
    2.979929e-11, 2.987291e-11, 2.985058e-11, 2.98732e-11, 2.975994e-11, 
    2.980844e-11, 2.970889e-11, 2.932297e-11, 2.943609e-11, 2.909946e-11, 
    2.889811e-11, 2.876482e-11, 2.867044e-11, 2.868377e-11, 2.870919e-11, 
    2.884005e-11, 2.896338e-11, 2.905758e-11, 2.912068e-11, 2.918294e-11, 
    2.937183e-11, 2.947211e-11, 2.969732e-11, 2.965661e-11, 2.97256e-11, 
    2.979161e-11, 2.990261e-11, 2.988432e-11, 2.993329e-11, 2.972379e-11, 
    2.986292e-11, 2.963343e-11, 2.96961e-11, 2.919986e-11, 2.901209e-11, 
    2.893247e-11, 2.88629e-11, 2.869402e-11, 2.881058e-11, 2.87646e-11, 
    2.887407e-11, 2.894375e-11, 2.890927e-11, 2.912241e-11, 2.903944e-11, 
    2.947805e-11, 2.928867e-11, 2.97839e-11, 2.966496e-11, 2.981245e-11, 
    2.973714e-11, 2.986625e-11, 2.975004e-11, 2.995152e-11, 2.99955e-11, 
    2.996544e-11, 3.008099e-11, 2.974361e-11, 2.987291e-11, 2.890831e-11, 
    2.891393e-11, 2.894012e-11, 2.882508e-11, 2.881805e-11, 2.871287e-11, 
    2.880645e-11, 2.884635e-11, 2.894779e-11, 2.900788e-11, 2.906508e-11, 
    2.919105e-11, 2.933211e-11, 2.953001e-11, 2.967267e-11, 2.976851e-11, 
    2.970972e-11, 2.976162e-11, 2.97036e-11, 2.967643e-11, 2.997901e-11, 
    2.980889e-11, 3.006436e-11, 3.005019e-11, 2.993445e-11, 3.005178e-11, 
    2.891788e-11, 2.888554e-11, 2.877342e-11, 2.886114e-11, 2.870143e-11, 
    2.879076e-11, 2.88422e-11, 2.904117e-11, 2.908499e-11, 2.912566e-11, 
    2.920607e-11, 2.930945e-11, 2.949132e-11, 2.965008e-11, 2.979545e-11, 
    2.978479e-11, 2.978854e-11, 2.982107e-11, 2.974054e-11, 2.983429e-11, 
    2.985005e-11, 2.980887e-11, 3.004829e-11, 2.997978e-11, 3.004989e-11, 
    3.000527e-11, 2.889605e-11, 2.895048e-11, 2.892106e-11, 2.89764e-11, 
    2.893741e-11, 2.911103e-11, 2.916321e-11, 2.940804e-11, 2.930742e-11, 
    2.946765e-11, 2.932367e-11, 2.934916e-11, 2.947288e-11, 2.933145e-11, 
    2.964131e-11, 2.943103e-11, 2.982233e-11, 2.961159e-11, 2.983556e-11, 
    2.979482e-11, 2.98623e-11, 2.99228e-11, 2.999903e-11, 3.013996e-11, 
    3.010729e-11, 3.022537e-11, 2.903175e-11, 2.910255e-11, 2.909632e-11, 
    2.917051e-11, 2.922546e-11, 2.934475e-11, 2.953665e-11, 2.946441e-11, 
    2.959712e-11, 2.962381e-11, 2.942221e-11, 2.954589e-11, 2.915e-11, 
    2.921375e-11, 2.917578e-11, 2.903733e-11, 2.948104e-11, 2.925285e-11, 
    2.967503e-11, 2.955081e-11, 2.991417e-11, 2.973315e-11, 3.008932e-11, 
    3.024232e-11, 3.038675e-11, 3.055602e-11, 2.914124e-11, 2.909308e-11, 
    2.917935e-11, 2.929893e-11, 2.941015e-11, 2.955838e-11, 2.957357e-11, 
    2.960139e-11, 2.967354e-11, 2.973427e-11, 2.961019e-11, 2.974951e-11, 
    2.922855e-11, 2.950089e-11, 2.907489e-11, 2.920279e-11, 2.929188e-11, 
    2.925278e-11, 2.945616e-11, 2.95042e-11, 2.969992e-11, 2.959866e-11, 
    3.020451e-11, 2.993559e-11, 3.068529e-11, 3.047469e-11, 2.907627e-11, 
    2.914107e-11, 2.936728e-11, 2.925953e-11, 2.956829e-11, 2.964457e-11, 
    2.970667e-11, 2.978616e-11, 2.979476e-11, 2.984192e-11, 2.976466e-11, 
    2.983886e-11, 2.95587e-11, 2.968371e-11, 2.934138e-11, 2.942448e-11, 
    2.938624e-11, 2.934431e-11, 2.947382e-11, 2.961214e-11, 2.961511e-11, 
    2.965954e-11, 2.978496e-11, 2.956955e-11, 3.023931e-11, 2.982466e-11, 
    2.921184e-11, 2.933708e-11, 2.9355e-11, 2.930643e-11, 2.963692e-11, 
    2.951693e-11, 2.984077e-11, 2.975304e-11, 2.989686e-11, 2.982534e-11, 
    2.981483e-11, 2.972315e-11, 2.966614e-11, 2.952242e-11, 2.940578e-11, 
    2.931347e-11, 2.933492e-11, 2.943637e-11, 2.962062e-11, 2.979553e-11, 
    2.975717e-11, 2.988591e-11, 2.954584e-11, 2.968817e-11, 2.963311e-11, 
    2.977679e-11, 2.946249e-11, 2.973e-11, 2.939433e-11, 2.942367e-11, 
    2.951455e-11, 2.969783e-11, 2.973847e-11, 2.97819e-11, 2.975509e-11, 
    2.962531e-11, 2.960407e-11, 2.951234e-11, 2.948703e-11, 2.941728e-11, 
    2.935961e-11, 2.94123e-11, 2.94677e-11, 2.962536e-11, 2.976785e-11, 
    2.992366e-11, 2.996187e-11, 3.014463e-11, 2.99958e-11, 3.024163e-11, 
    3.003256e-11, 3.039503e-11, 2.974555e-11, 3.002642e-11, 2.951869e-11, 
    2.957315e-11, 2.96718e-11, 2.989876e-11, 2.977611e-11, 2.991959e-11, 
    2.960324e-11, 2.943987e-11, 2.939769e-11, 2.931908e-11, 2.939949e-11, 
    2.939294e-11, 2.947e-11, 2.944522e-11, 2.96306e-11, 2.953094e-11, 
    2.981457e-11, 2.991846e-11, 3.021298e-11, 3.039436e-11, 3.057966e-11, 
    3.066167e-11, 3.068665e-11, 3.069711e-11,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
