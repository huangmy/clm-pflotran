netcdf ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-4.clm2.h0.0001-12-02-00000 {
dimensions:
	lndgrid = 338 ;
	gridcell = 338 ;
	landunit = 1352 ;
	column = 5408 ;
	pft = 10816 ;
	levgrnd = 15 ;
	levurb = 5 ;
	levlak = 10 ;
	numrad = 2 ;
	levsno = 5 ;
	ltype = 9 ;
	natpft = 17 ;
	string_length = 8 ;
	levdcmp = 15 ;
	hist_interval = 2 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float levgrnd(levgrnd) ;
		levgrnd:long_name = "coordinate soil levels" ;
		levgrnd:units = "m" ;
	float levlak(levlak) ;
		levlak:long_name = "coordinate lake levels" ;
		levlak:units = "m" ;
	float levdcmp(levdcmp) ;
		levdcmp:long_name = "coordinate soil levels" ;
		levdcmp:units = "m" ;
	float time(time) ;
		time:long_name = "time" ;
		time:units = "days since 0001-12-01 00:00:00" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bounds" ;
	int mcdate(time) ;
		mcdate:long_name = "current date (YYYYMMDD)" ;
	int mcsec(time) ;
		mcsec:long_name = "current seconds of current date" ;
		mcsec:units = "s" ;
	int mdcur(time) ;
		mdcur:long_name = "current day (from base day)" ;
	int mscur(time) ;
		mscur:long_name = "current seconds of current day" ;
	int nstep(time) ;
		nstep:long_name = "time step" ;
	double time_bounds(time, hist_interval) ;
		time_bounds:long_name = "history time interval endpoints" ;
	char date_written(time, string_length) ;
	char time_written(time, string_length) ;
	float lon(lndgrid) ;
		lon:long_name = "coordinate longitude" ;
		lon:units = "degrees_east" ;
		lon:_FillValue = 1.e+36f ;
		lon:missing_value = 1.e+36f ;
	float lat(lndgrid) ;
		lat:long_name = "coordinate latitude" ;
		lat:units = "degrees_north" ;
		lat:_FillValue = 1.e+36f ;
		lat:missing_value = 1.e+36f ;
	float area(lndgrid) ;
		area:long_name = "grid cell areas" ;
		area:units = "km^2" ;
		area:_FillValue = 1.e+36f ;
		area:missing_value = 1.e+36f ;
	float topo(lndgrid) ;
		topo:long_name = "grid cell topography" ;
		topo:units = "m" ;
		topo:_FillValue = 1.e+36f ;
		topo:missing_value = 1.e+36f ;
	float landfrac(lndgrid) ;
		landfrac:long_name = "land fraction" ;
		landfrac:_FillValue = 1.e+36f ;
		landfrac:missing_value = 1.e+36f ;
	int landmask(lndgrid) ;
		landmask:long_name = "land/ocean mask (0.=ocean and 1.=land)" ;
		landmask:_FillValue = -9999 ;
		landmask:missing_value = -9999 ;
	int pftmask(lndgrid) ;
		pftmask:long_name = "pft real/fake mask (0.=fake and 1.=real)" ;
		pftmask:_FillValue = -9999 ;
		pftmask:missing_value = -9999 ;
	float ACTUAL_IMMOB(time, lndgrid) ;
		ACTUAL_IMMOB:long_name = "actual N immobilization" ;
		ACTUAL_IMMOB:units = "gN/m^2/s" ;
		ACTUAL_IMMOB:cell_methods = "time: mean" ;
		ACTUAL_IMMOB:_FillValue = 1.e+36f ;
		ACTUAL_IMMOB:missing_value = 1.e+36f ;
	float AGNPP(time, lndgrid) ;
		AGNPP:long_name = "aboveground NPP" ;
		AGNPP:units = "gC/m^2/s" ;
		AGNPP:cell_methods = "time: mean" ;
		AGNPP:_FillValue = 1.e+36f ;
		AGNPP:missing_value = 1.e+36f ;
	float ALT(time, lndgrid) ;
		ALT:long_name = "current active layer thickness" ;
		ALT:units = "m" ;
		ALT:cell_methods = "time: mean" ;
		ALT:_FillValue = 1.e+36f ;
		ALT:missing_value = 1.e+36f ;
	float ALTMAX(time, lndgrid) ;
		ALTMAX:long_name = "maximum annual active layer thickness" ;
		ALTMAX:units = "m" ;
		ALTMAX:cell_methods = "time: mean" ;
		ALTMAX:_FillValue = 1.e+36f ;
		ALTMAX:missing_value = 1.e+36f ;
	float ALTMAX_LASTYEAR(time, lndgrid) ;
		ALTMAX_LASTYEAR:long_name = "maximum prior year active layer thickness" ;
		ALTMAX_LASTYEAR:units = "m" ;
		ALTMAX_LASTYEAR:cell_methods = "time: mean" ;
		ALTMAX_LASTYEAR:_FillValue = 1.e+36f ;
		ALTMAX_LASTYEAR:missing_value = 1.e+36f ;
	float AR(time, lndgrid) ;
		AR:long_name = "autotrophic respiration (MR + GR)" ;
		AR:units = "gC/m^2/s" ;
		AR:cell_methods = "time: mean" ;
		AR:_FillValue = 1.e+36f ;
		AR:missing_value = 1.e+36f ;
	float BAF_CROP(time, lndgrid) ;
		BAF_CROP:long_name = "fractional area burned for crop" ;
		BAF_CROP:units = "proportion/sec" ;
		BAF_CROP:cell_methods = "time: mean" ;
		BAF_CROP:_FillValue = 1.e+36f ;
		BAF_CROP:missing_value = 1.e+36f ;
	float BAF_PEATF(time, lndgrid) ;
		BAF_PEATF:long_name = "fractional area burned in peatland" ;
		BAF_PEATF:units = "proportion/sec" ;
		BAF_PEATF:cell_methods = "time: mean" ;
		BAF_PEATF:_FillValue = 1.e+36f ;
		BAF_PEATF:missing_value = 1.e+36f ;
	float BCDEP(time, lndgrid) ;
		BCDEP:long_name = "total BC deposition (dry+wet) from atmosphere" ;
		BCDEP:units = "kg/m^2/s" ;
		BCDEP:cell_methods = "time: mean" ;
		BCDEP:_FillValue = 1.e+36f ;
		BCDEP:missing_value = 1.e+36f ;
	float BGNPP(time, lndgrid) ;
		BGNPP:long_name = "belowground NPP" ;
		BGNPP:units = "gC/m^2/s" ;
		BGNPP:cell_methods = "time: mean" ;
		BGNPP:_FillValue = 1.e+36f ;
		BGNPP:missing_value = 1.e+36f ;
	float BTRAN(time, lndgrid) ;
		BTRAN:long_name = "transpiration beta factor" ;
		BTRAN:units = "unitless" ;
		BTRAN:cell_methods = "time: mean" ;
		BTRAN:_FillValue = 1.e+36f ;
		BTRAN:missing_value = 1.e+36f ;
	float BUILDHEAT(time, lndgrid) ;
		BUILDHEAT:long_name = "heat flux from urban building interior to walls and roof" ;
		BUILDHEAT:units = "W/m^2" ;
		BUILDHEAT:cell_methods = "time: mean" ;
		BUILDHEAT:_FillValue = 1.e+36f ;
		BUILDHEAT:missing_value = 1.e+36f ;
	float CH4PROD(time, lndgrid) ;
		CH4PROD:long_name = "Gridcell total production of CH4" ;
		CH4PROD:units = "gC/m2/s" ;
		CH4PROD:cell_methods = "time: mean" ;
		CH4PROD:_FillValue = 1.e+36f ;
		CH4PROD:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_SAT(time, lndgrid) ;
		CH4_SURF_AERE_SAT:long_name = "aerenchyma surface CH4 flux for inundated area; (+ to atm)" ;
		CH4_SURF_AERE_SAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_SAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_AERE_UNSAT(time, lndgrid) ;
		CH4_SURF_AERE_UNSAT:long_name = "aerenchyma surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_AERE_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_AERE_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_AERE_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_AERE_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_SAT(time, lndgrid) ;
		CH4_SURF_DIFF_SAT:long_name = "diffusive surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_DIFF_SAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_SAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_DIFF_UNSAT(time, lndgrid) ;
		CH4_SURF_DIFF_UNSAT:long_name = "diffusive surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_DIFF_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_DIFF_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_DIFF_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_DIFF_UNSAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_SAT(time, lndgrid) ;
		CH4_SURF_EBUL_SAT:long_name = "ebullition surface CH4 flux for inundated / lake area; (+ to atm)" ;
		CH4_SURF_EBUL_SAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_SAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_SAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_SAT:missing_value = 1.e+36f ;
	float CH4_SURF_EBUL_UNSAT(time, lndgrid) ;
		CH4_SURF_EBUL_UNSAT:long_name = "ebullition surface CH4 flux for non-inundated area; (+ to atm)" ;
		CH4_SURF_EBUL_UNSAT:units = "mol/m2/s" ;
		CH4_SURF_EBUL_UNSAT:cell_methods = "time: mean" ;
		CH4_SURF_EBUL_UNSAT:_FillValue = 1.e+36f ;
		CH4_SURF_EBUL_UNSAT:missing_value = 1.e+36f ;
	float COL_CTRUNC(time, lndgrid) ;
		COL_CTRUNC:long_name = "column-level sink for C truncation" ;
		COL_CTRUNC:units = "gC/m^2" ;
		COL_CTRUNC:cell_methods = "time: mean" ;
		COL_CTRUNC:_FillValue = 1.e+36f ;
		COL_CTRUNC:missing_value = 1.e+36f ;
	float COL_FIRE_CLOSS(time, lndgrid) ;
		COL_FIRE_CLOSS:long_name = "total column-level fire C loss for non-peat fires outside land-type converted region" ;
		COL_FIRE_CLOSS:units = "gC/m^2/s" ;
		COL_FIRE_CLOSS:cell_methods = "time: mean" ;
		COL_FIRE_CLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_CLOSS:missing_value = 1.e+36f ;
	float COL_FIRE_NLOSS(time, lndgrid) ;
		COL_FIRE_NLOSS:long_name = "total column-level fire N loss" ;
		COL_FIRE_NLOSS:units = "gN/m^2/s" ;
		COL_FIRE_NLOSS:cell_methods = "time: mean" ;
		COL_FIRE_NLOSS:_FillValue = 1.e+36f ;
		COL_FIRE_NLOSS:missing_value = 1.e+36f ;
	float COL_NTRUNC(time, lndgrid) ;
		COL_NTRUNC:long_name = "column-level sink for N truncation" ;
		COL_NTRUNC:units = "gN/m^2" ;
		COL_NTRUNC:cell_methods = "time: mean" ;
		COL_NTRUNC:_FillValue = 1.e+36f ;
		COL_NTRUNC:missing_value = 1.e+36f ;
	float CONC_CH4_SAT(time, levgrnd, lndgrid) ;
		CONC_CH4_SAT:long_name = "CH4 soil Concentration for inundated / lake area" ;
		CONC_CH4_SAT:units = "mol/m3" ;
		CONC_CH4_SAT:cell_methods = "time: mean" ;
		CONC_CH4_SAT:_FillValue = 1.e+36f ;
		CONC_CH4_SAT:missing_value = 1.e+36f ;
	float CONC_CH4_UNSAT(time, levgrnd, lndgrid) ;
		CONC_CH4_UNSAT:long_name = "CH4 soil Concentration for non-inundated area" ;
		CONC_CH4_UNSAT:units = "mol/m3" ;
		CONC_CH4_UNSAT:cell_methods = "time: mean" ;
		CONC_CH4_UNSAT:_FillValue = 1.e+36f ;
		CONC_CH4_UNSAT:missing_value = 1.e+36f ;
	float CONC_O2_SAT(time, levgrnd, lndgrid) ;
		CONC_O2_SAT:long_name = "O2 soil Concentration for inundated / lake area" ;
		CONC_O2_SAT:units = "mol/m3" ;
		CONC_O2_SAT:cell_methods = "time: mean" ;
		CONC_O2_SAT:_FillValue = 1.e+36f ;
		CONC_O2_SAT:missing_value = 1.e+36f ;
	float CONC_O2_UNSAT(time, levgrnd, lndgrid) ;
		CONC_O2_UNSAT:long_name = "O2 soil Concentration for non-inundated area" ;
		CONC_O2_UNSAT:units = "mol/m3" ;
		CONC_O2_UNSAT:cell_methods = "time: mean" ;
		CONC_O2_UNSAT:_FillValue = 1.e+36f ;
		CONC_O2_UNSAT:missing_value = 1.e+36f ;
	float CPOOL(time, lndgrid) ;
		CPOOL:long_name = "temporary photosynthate C pool" ;
		CPOOL:units = "gC/m^2" ;
		CPOOL:cell_methods = "time: mean" ;
		CPOOL:_FillValue = 1.e+36f ;
		CPOOL:missing_value = 1.e+36f ;
	float CWDC(time, lndgrid) ;
		CWDC:long_name = "CWD C" ;
		CWDC:units = "gC/m^2" ;
		CWDC:cell_methods = "time: mean" ;
		CWDC:_FillValue = 1.e+36f ;
		CWDC:missing_value = 1.e+36f ;
	float CWDC_HR(time, lndgrid) ;
		CWDC_HR:long_name = "coarse woody debris C heterotrophic respiration" ;
		CWDC_HR:units = "gC/m^2/s" ;
		CWDC_HR:cell_methods = "time: mean" ;
		CWDC_HR:_FillValue = 1.e+36f ;
		CWDC_HR:missing_value = 1.e+36f ;
	float CWDC_LOSS(time, lndgrid) ;
		CWDC_LOSS:long_name = "coarse woody debris C loss" ;
		CWDC_LOSS:units = "gC/m^2/s" ;
		CWDC_LOSS:cell_methods = "time: mean" ;
		CWDC_LOSS:_FillValue = 1.e+36f ;
		CWDC_LOSS:missing_value = 1.e+36f ;
	float CWDC_TO_LITR2C(time, lndgrid) ;
		CWDC_TO_LITR2C:long_name = "decomp. of coarse woody debris C to litter 2 C" ;
		CWDC_TO_LITR2C:units = "gC/m^2/s" ;
		CWDC_TO_LITR2C:cell_methods = "time: mean" ;
		CWDC_TO_LITR2C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR2C:missing_value = 1.e+36f ;
	float CWDC_TO_LITR3C(time, lndgrid) ;
		CWDC_TO_LITR3C:long_name = "decomp. of coarse woody debris C to litter 3 C" ;
		CWDC_TO_LITR3C:units = "gC/m^2/s" ;
		CWDC_TO_LITR3C:cell_methods = "time: mean" ;
		CWDC_TO_LITR3C:_FillValue = 1.e+36f ;
		CWDC_TO_LITR3C:missing_value = 1.e+36f ;
	float CWDC_vr(time, levdcmp, lndgrid) ;
		CWDC_vr:long_name = "CWD C (vertically resolved)" ;
		CWDC_vr:units = "gC/m^3" ;
		CWDC_vr:cell_methods = "time: mean" ;
		CWDC_vr:_FillValue = 1.e+36f ;
		CWDC_vr:missing_value = 1.e+36f ;
	float CWDN(time, lndgrid) ;
		CWDN:long_name = "CWD N" ;
		CWDN:units = "gN/m^2" ;
		CWDN:cell_methods = "time: mean" ;
		CWDN:_FillValue = 1.e+36f ;
		CWDN:missing_value = 1.e+36f ;
	float CWDN_TO_LITR2N(time, lndgrid) ;
		CWDN_TO_LITR2N:long_name = "decomp. of coarse woody debris N to litter 2 N" ;
		CWDN_TO_LITR2N:units = "gN/m^2" ;
		CWDN_TO_LITR2N:cell_methods = "time: mean" ;
		CWDN_TO_LITR2N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR2N:missing_value = 1.e+36f ;
	float CWDN_TO_LITR3N(time, lndgrid) ;
		CWDN_TO_LITR3N:long_name = "decomp. of coarse woody debris N to litter 3 N" ;
		CWDN_TO_LITR3N:units = "gN/m^2" ;
		CWDN_TO_LITR3N:cell_methods = "time: mean" ;
		CWDN_TO_LITR3N:_FillValue = 1.e+36f ;
		CWDN_TO_LITR3N:missing_value = 1.e+36f ;
	float CWDN_vr(time, levdcmp, lndgrid) ;
		CWDN_vr:long_name = "CWD N (vertically resolved)" ;
		CWDN_vr:units = "gN/m^3" ;
		CWDN_vr:cell_methods = "time: mean" ;
		CWDN_vr:_FillValue = 1.e+36f ;
		CWDN_vr:missing_value = 1.e+36f ;
	float DEADCROOTC(time, lndgrid) ;
		DEADCROOTC:long_name = "dead coarse root C" ;
		DEADCROOTC:units = "gC/m^2" ;
		DEADCROOTC:cell_methods = "time: mean" ;
		DEADCROOTC:_FillValue = 1.e+36f ;
		DEADCROOTC:missing_value = 1.e+36f ;
	float DEADCROOTN(time, lndgrid) ;
		DEADCROOTN:long_name = "dead coarse root N" ;
		DEADCROOTN:units = "gN/m^2" ;
		DEADCROOTN:cell_methods = "time: mean" ;
		DEADCROOTN:_FillValue = 1.e+36f ;
		DEADCROOTN:missing_value = 1.e+36f ;
	float DEADSTEMC(time, lndgrid) ;
		DEADSTEMC:long_name = "dead stem C" ;
		DEADSTEMC:units = "gC/m^2" ;
		DEADSTEMC:cell_methods = "time: mean" ;
		DEADSTEMC:_FillValue = 1.e+36f ;
		DEADSTEMC:missing_value = 1.e+36f ;
	float DEADSTEMN(time, lndgrid) ;
		DEADSTEMN:long_name = "dead stem N" ;
		DEADSTEMN:units = "gN/m^2" ;
		DEADSTEMN:cell_methods = "time: mean" ;
		DEADSTEMN:_FillValue = 1.e+36f ;
		DEADSTEMN:missing_value = 1.e+36f ;
	float DENIT(time, lndgrid) ;
		DENIT:long_name = "total rate of denitrification" ;
		DENIT:units = "gN/m^2/s" ;
		DENIT:cell_methods = "time: mean" ;
		DENIT:_FillValue = 1.e+36f ;
		DENIT:missing_value = 1.e+36f ;
	float DISPVEGC(time, lndgrid) ;
		DISPVEGC:long_name = "displayed veg carbon, excluding storage and cpool" ;
		DISPVEGC:units = "gC/m^2" ;
		DISPVEGC:cell_methods = "time: mean" ;
		DISPVEGC:_FillValue = 1.e+36f ;
		DISPVEGC:missing_value = 1.e+36f ;
	float DISPVEGN(time, lndgrid) ;
		DISPVEGN:long_name = "displayed vegetation nitrogen" ;
		DISPVEGN:units = "gN/m^2" ;
		DISPVEGN:cell_methods = "time: mean" ;
		DISPVEGN:_FillValue = 1.e+36f ;
		DISPVEGN:missing_value = 1.e+36f ;
	float DSTDEP(time, lndgrid) ;
		DSTDEP:long_name = "total dust deposition (dry+wet) from atmosphere" ;
		DSTDEP:units = "kg/m^2/s" ;
		DSTDEP:cell_methods = "time: mean" ;
		DSTDEP:_FillValue = 1.e+36f ;
		DSTDEP:missing_value = 1.e+36f ;
	float DSTFLXT(time, lndgrid) ;
		DSTFLXT:long_name = "total surface dust emission" ;
		DSTFLXT:units = "kg/m2/s" ;
		DSTFLXT:cell_methods = "time: mean" ;
		DSTFLXT:_FillValue = 1.e+36f ;
		DSTFLXT:missing_value = 1.e+36f ;
	float DWT_CLOSS(time, lndgrid) ;
		DWT_CLOSS:long_name = "total carbon loss from land cover conversion" ;
		DWT_CLOSS:units = "gC/m^2/s" ;
		DWT_CLOSS:cell_methods = "time: mean" ;
		DWT_CLOSS:_FillValue = 1.e+36f ;
		DWT_CLOSS:missing_value = 1.e+36f ;
	float DWT_CONV_CFLUX(time, lndgrid) ;
		DWT_CONV_CFLUX:long_name = "conversion C flux (immediate loss to atm)" ;
		DWT_CONV_CFLUX:units = "gC/m^2/s" ;
		DWT_CONV_CFLUX:cell_methods = "time: mean" ;
		DWT_CONV_CFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_CFLUX:missing_value = 1.e+36f ;
	float DWT_CONV_NFLUX(time, lndgrid) ;
		DWT_CONV_NFLUX:long_name = "conversion N flux (immediate loss to atm)" ;
		DWT_CONV_NFLUX:units = "gN/m^2/s" ;
		DWT_CONV_NFLUX:cell_methods = "time: mean" ;
		DWT_CONV_NFLUX:_FillValue = 1.e+36f ;
		DWT_CONV_NFLUX:missing_value = 1.e+36f ;
	float DWT_NLOSS(time, lndgrid) ;
		DWT_NLOSS:long_name = "total nitrogen loss from landcover conversion" ;
		DWT_NLOSS:units = "gN/m^2/s" ;
		DWT_NLOSS:cell_methods = "time: mean" ;
		DWT_NLOSS:_FillValue = 1.e+36f ;
		DWT_NLOSS:missing_value = 1.e+36f ;
	float DWT_PROD100C_GAIN(time, lndgrid) ;
		DWT_PROD100C_GAIN:long_name = "landcover change-driven addition to 100-yr wood product pool" ;
		DWT_PROD100C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD100C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD100N_GAIN(time, lndgrid) ;
		DWT_PROD100N_GAIN:long_name = "addition to 100-yr wood product pool" ;
		DWT_PROD100N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD100N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD100N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD100N_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10C_GAIN(time, lndgrid) ;
		DWT_PROD10C_GAIN:long_name = "landcover change-driven addition to 10-yr wood product pool" ;
		DWT_PROD10C_GAIN:units = "gC/m^2/s" ;
		DWT_PROD10C_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10C_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10C_GAIN:missing_value = 1.e+36f ;
	float DWT_PROD10N_GAIN(time, lndgrid) ;
		DWT_PROD10N_GAIN:long_name = "addition to 10-yr wood product pool" ;
		DWT_PROD10N_GAIN:units = "gN/m^2/s" ;
		DWT_PROD10N_GAIN:cell_methods = "time: mean" ;
		DWT_PROD10N_GAIN:_FillValue = 1.e+36f ;
		DWT_PROD10N_GAIN:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDC_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDC_TO_DEADSTEM:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDC_TO_LEAF(time, lndgrid) ;
		DWT_SEEDC_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDC_TO_LEAF:units = "gC/m^2/s" ;
		DWT_SEEDC_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDC_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDC_TO_LEAF:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_DEADSTEM(time, lndgrid) ;
		DWT_SEEDN_TO_DEADSTEM:long_name = "seed source to PFT-level deadstem" ;
		DWT_SEEDN_TO_DEADSTEM:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_DEADSTEM:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_DEADSTEM:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_DEADSTEM:missing_value = 1.e+36f ;
	float DWT_SEEDN_TO_LEAF(time, lndgrid) ;
		DWT_SEEDN_TO_LEAF:long_name = "seed source to PFT-level leaf" ;
		DWT_SEEDN_TO_LEAF:units = "gN/m^2/s" ;
		DWT_SEEDN_TO_LEAF:cell_methods = "time: mean" ;
		DWT_SEEDN_TO_LEAF:_FillValue = 1.e+36f ;
		DWT_SEEDN_TO_LEAF:missing_value = 1.e+36f ;
	float EFLX_DYNBAL(time, lndgrid) ;
		EFLX_DYNBAL:long_name = "dynamic land cover change conversion energy flux" ;
		EFLX_DYNBAL:units = "W/m^2" ;
		EFLX_DYNBAL:cell_methods = "time: mean" ;
		EFLX_DYNBAL:_FillValue = 1.e+36f ;
		EFLX_DYNBAL:missing_value = 1.e+36f ;
	float EFLX_GRND_LAKE(time, lndgrid) ;
		EFLX_GRND_LAKE:long_name = "net heat flux into lake/snow surface, excluding light transmission" ;
		EFLX_GRND_LAKE:units = "W/m^2" ;
		EFLX_GRND_LAKE:cell_methods = "time: mean" ;
		EFLX_GRND_LAKE:_FillValue = 1.e+36f ;
		EFLX_GRND_LAKE:missing_value = 1.e+36f ;
	float EFLX_LH_TOT(time, lndgrid) ;
		EFLX_LH_TOT:long_name = "total latent heat flux [+ to atm]" ;
		EFLX_LH_TOT:units = "W/m^2" ;
		EFLX_LH_TOT:cell_methods = "time: mean" ;
		EFLX_LH_TOT:_FillValue = 1.e+36f ;
		EFLX_LH_TOT:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_R(time, lndgrid) ;
		EFLX_LH_TOT_R:long_name = "Rural total evaporation" ;
		EFLX_LH_TOT_R:units = "W/m^2" ;
		EFLX_LH_TOT_R:cell_methods = "time: mean" ;
		EFLX_LH_TOT_R:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_R:missing_value = 1.e+36f ;
	float EFLX_LH_TOT_U(time, lndgrid) ;
		EFLX_LH_TOT_U:long_name = "Urban total evaporation" ;
		EFLX_LH_TOT_U:units = "W/m^2" ;
		EFLX_LH_TOT_U:cell_methods = "time: mean" ;
		EFLX_LH_TOT_U:_FillValue = 1.e+36f ;
		EFLX_LH_TOT_U:missing_value = 1.e+36f ;
	float ELAI(time, lndgrid) ;
		ELAI:long_name = "exposed one-sided leaf area index" ;
		ELAI:units = "m^2/m^2" ;
		ELAI:cell_methods = "time: mean" ;
		ELAI:_FillValue = 1.e+36f ;
		ELAI:missing_value = 1.e+36f ;
	float ER(time, lndgrid) ;
		ER:long_name = "total ecosystem respiration, autotrophic + heterotrophic" ;
		ER:units = "gC/m^2/s" ;
		ER:cell_methods = "time: mean" ;
		ER:_FillValue = 1.e+36f ;
		ER:missing_value = 1.e+36f ;
	float ERRH2O(time, lndgrid) ;
		ERRH2O:long_name = "total water conservation error" ;
		ERRH2O:units = "mm" ;
		ERRH2O:cell_methods = "time: mean" ;
		ERRH2O:_FillValue = 1.e+36f ;
		ERRH2O:missing_value = 1.e+36f ;
	float ERRH2OSNO(time, lndgrid) ;
		ERRH2OSNO:long_name = "imbalance in snow depth (liquid water)" ;
		ERRH2OSNO:units = "mm" ;
		ERRH2OSNO:cell_methods = "time: mean" ;
		ERRH2OSNO:_FillValue = 1.e+36f ;
		ERRH2OSNO:missing_value = 1.e+36f ;
	float ERRSEB(time, lndgrid) ;
		ERRSEB:long_name = "surface energy conservation error" ;
		ERRSEB:units = "W/m^2" ;
		ERRSEB:cell_methods = "time: mean" ;
		ERRSEB:_FillValue = 1.e+36f ;
		ERRSEB:missing_value = 1.e+36f ;
	float ERRSOI(time, lndgrid) ;
		ERRSOI:long_name = "soil/lake energy conservation error" ;
		ERRSOI:units = "W/m^2" ;
		ERRSOI:cell_methods = "time: mean" ;
		ERRSOI:_FillValue = 1.e+36f ;
		ERRSOI:missing_value = 1.e+36f ;
	float ERRSOL(time, lndgrid) ;
		ERRSOL:long_name = "solar radiation conservation error" ;
		ERRSOL:units = "W/m^2" ;
		ERRSOL:cell_methods = "time: mean" ;
		ERRSOL:_FillValue = 1.e+36f ;
		ERRSOL:missing_value = 1.e+36f ;
	float ESAI(time, lndgrid) ;
		ESAI:long_name = "exposed one-sided stem area index" ;
		ESAI:units = "m^2/m^2" ;
		ESAI:cell_methods = "time: mean" ;
		ESAI:_FillValue = 1.e+36f ;
		ESAI:missing_value = 1.e+36f ;
	float FAREA_BURNED(time, lndgrid) ;
		FAREA_BURNED:long_name = "fractional area burned" ;
		FAREA_BURNED:units = "proportion/sec" ;
		FAREA_BURNED:cell_methods = "time: mean" ;
		FAREA_BURNED:_FillValue = 1.e+36f ;
		FAREA_BURNED:missing_value = 1.e+36f ;
	float FCEV(time, lndgrid) ;
		FCEV:long_name = "canopy evaporation" ;
		FCEV:units = "W/m^2" ;
		FCEV:cell_methods = "time: mean" ;
		FCEV:_FillValue = 1.e+36f ;
		FCEV:missing_value = 1.e+36f ;
	float FCH4(time, lndgrid) ;
		FCH4:long_name = "Gridcell surface CH4 flux to atmosphere (+ to atm)" ;
		FCH4:units = "kgC/m2/s" ;
		FCH4:cell_methods = "time: mean" ;
		FCH4:_FillValue = 1.e+36f ;
		FCH4:missing_value = 1.e+36f ;
	float FCH4TOCO2(time, lndgrid) ;
		FCH4TOCO2:long_name = "Gridcell oxidation of CH4 to CO2" ;
		FCH4TOCO2:units = "gC/m2/s" ;
		FCH4TOCO2:cell_methods = "time: mean" ;
		FCH4TOCO2:_FillValue = 1.e+36f ;
		FCH4TOCO2:missing_value = 1.e+36f ;
	float FCH4_DFSAT(time, lndgrid) ;
		FCH4_DFSAT:long_name = "CH4 additional flux due to changing fsat, vegetated landunits only" ;
		FCH4_DFSAT:units = "kgC/m2/s" ;
		FCH4_DFSAT:cell_methods = "time: mean" ;
		FCH4_DFSAT:_FillValue = 1.e+36f ;
		FCH4_DFSAT:missing_value = 1.e+36f ;
	float FCOV(time, lndgrid) ;
		FCOV:long_name = "fractional impermeable area" ;
		FCOV:units = "unitless" ;
		FCOV:cell_methods = "time: mean" ;
		FCOV:_FillValue = 1.e+36f ;
		FCOV:missing_value = 1.e+36f ;
	float FCTR(time, lndgrid) ;
		FCTR:long_name = "canopy transpiration" ;
		FCTR:units = "W/m^2" ;
		FCTR:cell_methods = "time: mean" ;
		FCTR:_FillValue = 1.e+36f ;
		FCTR:missing_value = 1.e+36f ;
	float FGEV(time, lndgrid) ;
		FGEV:long_name = "ground evaporation" ;
		FGEV:units = "W/m^2" ;
		FGEV:cell_methods = "time: mean" ;
		FGEV:_FillValue = 1.e+36f ;
		FGEV:missing_value = 1.e+36f ;
	float FGR(time, lndgrid) ;
		FGR:long_name = "heat flux into soil/snow including snow melt and lake / snow light transmission" ;
		FGR:units = "W/m^2" ;
		FGR:cell_methods = "time: mean" ;
		FGR:_FillValue = 1.e+36f ;
		FGR:missing_value = 1.e+36f ;
	float FGR12(time, lndgrid) ;
		FGR12:long_name = "heat flux between soil layers 1 and 2" ;
		FGR12:units = "W/m^2" ;
		FGR12:cell_methods = "time: mean" ;
		FGR12:_FillValue = 1.e+36f ;
		FGR12:missing_value = 1.e+36f ;
	float FGR_R(time, lndgrid) ;
		FGR_R:long_name = "Rural heat flux into soil/snow including snow melt and snow light transmission" ;
		FGR_R:units = "W/m^2" ;
		FGR_R:cell_methods = "time: mean" ;
		FGR_R:_FillValue = 1.e+36f ;
		FGR_R:missing_value = 1.e+36f ;
	float FGR_U(time, lndgrid) ;
		FGR_U:long_name = "Urban heat flux into soil/snow including snow melt" ;
		FGR_U:units = "W/m^2" ;
		FGR_U:cell_methods = "time: mean" ;
		FGR_U:_FillValue = 1.e+36f ;
		FGR_U:missing_value = 1.e+36f ;
	float FH2OSFC(time, lndgrid) ;
		FH2OSFC:long_name = "fraction of ground covered by surface water" ;
		FH2OSFC:units = "unitless" ;
		FH2OSFC:cell_methods = "time: mean" ;
		FH2OSFC:_FillValue = 1.e+36f ;
		FH2OSFC:missing_value = 1.e+36f ;
	float FINUNDATED(time, lndgrid) ;
		FINUNDATED:long_name = "fractional inundated area of vegetated columns" ;
		FINUNDATED:units = "unitless" ;
		FINUNDATED:cell_methods = "time: mean" ;
		FINUNDATED:_FillValue = 1.e+36f ;
		FINUNDATED:missing_value = 1.e+36f ;
	float FINUNDATED_LAG(time, lndgrid) ;
		FINUNDATED_LAG:long_name = "time-lagged inundated fraction of vegetated columns" ;
		FINUNDATED_LAG:units = "unitless" ;
		FINUNDATED_LAG:cell_methods = "time: mean" ;
		FINUNDATED_LAG:_FillValue = 1.e+36f ;
		FINUNDATED_LAG:missing_value = 1.e+36f ;
	float FIRA(time, lndgrid) ;
		FIRA:long_name = "net infrared (longwave) radiation" ;
		FIRA:units = "W/m^2" ;
		FIRA:cell_methods = "time: mean" ;
		FIRA:_FillValue = 1.e+36f ;
		FIRA:missing_value = 1.e+36f ;
	float FIRA_R(time, lndgrid) ;
		FIRA_R:long_name = "Rural net infrared (longwave) radiation" ;
		FIRA_R:units = "W/m^2" ;
		FIRA_R:cell_methods = "time: mean" ;
		FIRA_R:_FillValue = 1.e+36f ;
		FIRA_R:missing_value = 1.e+36f ;
	float FIRA_U(time, lndgrid) ;
		FIRA_U:long_name = "Urban net infrared (longwave) radiation" ;
		FIRA_U:units = "W/m^2" ;
		FIRA_U:cell_methods = "time: mean" ;
		FIRA_U:_FillValue = 1.e+36f ;
		FIRA_U:missing_value = 1.e+36f ;
	float FIRE(time, lndgrid) ;
		FIRE:long_name = "emitted infrared (longwave) radiation" ;
		FIRE:units = "W/m^2" ;
		FIRE:cell_methods = "time: mean" ;
		FIRE:_FillValue = 1.e+36f ;
		FIRE:missing_value = 1.e+36f ;
	float FIRE_R(time, lndgrid) ;
		FIRE_R:long_name = "Rural emitted infrared (longwave) radiation" ;
		FIRE_R:units = "W/m^2" ;
		FIRE_R:cell_methods = "time: mean" ;
		FIRE_R:_FillValue = 1.e+36f ;
		FIRE_R:missing_value = 1.e+36f ;
	float FIRE_U(time, lndgrid) ;
		FIRE_U:long_name = "Urban emitted infrared (longwave) radiation" ;
		FIRE_U:units = "W/m^2" ;
		FIRE_U:cell_methods = "time: mean" ;
		FIRE_U:_FillValue = 1.e+36f ;
		FIRE_U:missing_value = 1.e+36f ;
	float FLDS(time, lndgrid) ;
		FLDS:long_name = "atmospheric longwave radiation" ;
		FLDS:units = "W/m^2" ;
		FLDS:cell_methods = "time: mean" ;
		FLDS:_FillValue = 1.e+36f ;
		FLDS:missing_value = 1.e+36f ;
	float FPG(time, lndgrid) ;
		FPG:long_name = "fraction of potential gpp" ;
		FPG:units = "proportion" ;
		FPG:cell_methods = "time: mean" ;
		FPG:_FillValue = 1.e+36f ;
		FPG:missing_value = 1.e+36f ;
	float FPI(time, lndgrid) ;
		FPI:long_name = "fraction of potential immobilization" ;
		FPI:units = "proportion" ;
		FPI:cell_methods = "time: mean" ;
		FPI:_FillValue = 1.e+36f ;
		FPI:missing_value = 1.e+36f ;
	float FPI_vr(time, levdcmp, lndgrid) ;
		FPI_vr:long_name = "fraction of potential immobilization" ;
		FPI_vr:units = "proportion" ;
		FPI_vr:cell_methods = "time: mean" ;
		FPI_vr:_FillValue = 1.e+36f ;
		FPI_vr:missing_value = 1.e+36f ;
	float FPSN(time, lndgrid) ;
		FPSN:long_name = "photosynthesis" ;
		FPSN:units = "umol/m2s" ;
		FPSN:cell_methods = "time: mean" ;
		FPSN:_FillValue = 1.e+36f ;
		FPSN:missing_value = 1.e+36f ;
	float FPSN_WC(time, lndgrid) ;
		FPSN_WC:long_name = "Rubisco-limited photosynthesis" ;
		FPSN_WC:units = "umol/m2s" ;
		FPSN_WC:cell_methods = "time: mean" ;
		FPSN_WC:_FillValue = 1.e+36f ;
		FPSN_WC:missing_value = 1.e+36f ;
	float FPSN_WJ(time, lndgrid) ;
		FPSN_WJ:long_name = "RuBP-limited photosynthesis" ;
		FPSN_WJ:units = "umol/m2s" ;
		FPSN_WJ:cell_methods = "time: mean" ;
		FPSN_WJ:_FillValue = 1.e+36f ;
		FPSN_WJ:missing_value = 1.e+36f ;
	float FPSN_WP(time, lndgrid) ;
		FPSN_WP:long_name = "Product-limited photosynthesis" ;
		FPSN_WP:units = "umol/m2s" ;
		FPSN_WP:cell_methods = "time: mean" ;
		FPSN_WP:_FillValue = 1.e+36f ;
		FPSN_WP:missing_value = 1.e+36f ;
	float FROOTC(time, lndgrid) ;
		FROOTC:long_name = "fine root C" ;
		FROOTC:units = "gC/m^2" ;
		FROOTC:cell_methods = "time: mean" ;
		FROOTC:_FillValue = 1.e+36f ;
		FROOTC:missing_value = 1.e+36f ;
	float FROOTC_ALLOC(time, lndgrid) ;
		FROOTC_ALLOC:long_name = "fine root C allocation" ;
		FROOTC_ALLOC:units = "gC/m^2/s" ;
		FROOTC_ALLOC:cell_methods = "time: mean" ;
		FROOTC_ALLOC:_FillValue = 1.e+36f ;
		FROOTC_ALLOC:missing_value = 1.e+36f ;
	float FROOTC_LOSS(time, lndgrid) ;
		FROOTC_LOSS:long_name = "fine root C loss" ;
		FROOTC_LOSS:units = "gC/m^2/s" ;
		FROOTC_LOSS:cell_methods = "time: mean" ;
		FROOTC_LOSS:_FillValue = 1.e+36f ;
		FROOTC_LOSS:missing_value = 1.e+36f ;
	float FROOTN(time, lndgrid) ;
		FROOTN:long_name = "fine root N" ;
		FROOTN:units = "gN/m^2" ;
		FROOTN:cell_methods = "time: mean" ;
		FROOTN:_FillValue = 1.e+36f ;
		FROOTN:missing_value = 1.e+36f ;
	float FROST_TABLE(time, lndgrid) ;
		FROST_TABLE:long_name = "frost table depth (vegetated landunits only)" ;
		FROST_TABLE:units = "m" ;
		FROST_TABLE:cell_methods = "time: mean" ;
		FROST_TABLE:_FillValue = 1.e+36f ;
		FROST_TABLE:missing_value = 1.e+36f ;
	float FSA(time, lndgrid) ;
		FSA:long_name = "absorbed solar radiation" ;
		FSA:units = "W/m^2" ;
		FSA:cell_methods = "time: mean" ;
		FSA:_FillValue = 1.e+36f ;
		FSA:missing_value = 1.e+36f ;
	float FSAT(time, lndgrid) ;
		FSAT:long_name = "fractional area with water table at surface" ;
		FSAT:units = "unitless" ;
		FSAT:cell_methods = "time: mean" ;
		FSAT:_FillValue = 1.e+36f ;
		FSAT:missing_value = 1.e+36f ;
	float FSA_R(time, lndgrid) ;
		FSA_R:long_name = "Rural absorbed solar radiation" ;
		FSA_R:units = "W/m^2" ;
		FSA_R:cell_methods = "time: mean" ;
		FSA_R:_FillValue = 1.e+36f ;
		FSA_R:missing_value = 1.e+36f ;
	float FSA_U(time, lndgrid) ;
		FSA_U:long_name = "Urban absorbed solar radiation" ;
		FSA_U:units = "W/m^2" ;
		FSA_U:cell_methods = "time: mean" ;
		FSA_U:_FillValue = 1.e+36f ;
		FSA_U:missing_value = 1.e+36f ;
	float FSDS(time, lndgrid) ;
		FSDS:long_name = "atmospheric incident solar radiation" ;
		FSDS:units = "W/m^2" ;
		FSDS:cell_methods = "time: mean" ;
		FSDS:_FillValue = 1.e+36f ;
		FSDS:missing_value = 1.e+36f ;
	float FSDSND(time, lndgrid) ;
		FSDSND:long_name = "direct nir incident solar radiation" ;
		FSDSND:units = "W/m^2" ;
		FSDSND:cell_methods = "time: mean" ;
		FSDSND:_FillValue = 1.e+36f ;
		FSDSND:missing_value = 1.e+36f ;
	float FSDSNDLN(time, lndgrid) ;
		FSDSNDLN:long_name = "direct nir incident solar radiation at local noon" ;
		FSDSNDLN:units = "W/m^2" ;
		FSDSNDLN:cell_methods = "time: mean" ;
		FSDSNDLN:_FillValue = 1.e+36f ;
		FSDSNDLN:missing_value = 1.e+36f ;
	float FSDSNI(time, lndgrid) ;
		FSDSNI:long_name = "diffuse nir incident solar radiation" ;
		FSDSNI:units = "W/m^2" ;
		FSDSNI:cell_methods = "time: mean" ;
		FSDSNI:_FillValue = 1.e+36f ;
		FSDSNI:missing_value = 1.e+36f ;
	float FSDSVD(time, lndgrid) ;
		FSDSVD:long_name = "direct vis incident solar radiation" ;
		FSDSVD:units = "W/m^2" ;
		FSDSVD:cell_methods = "time: mean" ;
		FSDSVD:_FillValue = 1.e+36f ;
		FSDSVD:missing_value = 1.e+36f ;
	float FSDSVDLN(time, lndgrid) ;
		FSDSVDLN:long_name = "direct vis incident solar radiation at local noon" ;
		FSDSVDLN:units = "W/m^2" ;
		FSDSVDLN:cell_methods = "time: mean" ;
		FSDSVDLN:_FillValue = 1.e+36f ;
		FSDSVDLN:missing_value = 1.e+36f ;
	float FSDSVI(time, lndgrid) ;
		FSDSVI:long_name = "diffuse vis incident solar radiation" ;
		FSDSVI:units = "W/m^2" ;
		FSDSVI:cell_methods = "time: mean" ;
		FSDSVI:_FillValue = 1.e+36f ;
		FSDSVI:missing_value = 1.e+36f ;
	float FSDSVILN(time, lndgrid) ;
		FSDSVILN:long_name = "diffuse vis incident solar radiation at local noon" ;
		FSDSVILN:units = "W/m^2" ;
		FSDSVILN:cell_methods = "time: mean" ;
		FSDSVILN:_FillValue = 1.e+36f ;
		FSDSVILN:missing_value = 1.e+36f ;
	float FSH(time, lndgrid) ;
		FSH:long_name = "sensible heat" ;
		FSH:units = "W/m^2" ;
		FSH:cell_methods = "time: mean" ;
		FSH:_FillValue = 1.e+36f ;
		FSH:missing_value = 1.e+36f ;
	float FSH_G(time, lndgrid) ;
		FSH_G:long_name = "sensible heat from ground" ;
		FSH_G:units = "W/m^2" ;
		FSH_G:cell_methods = "time: mean" ;
		FSH_G:_FillValue = 1.e+36f ;
		FSH_G:missing_value = 1.e+36f ;
	float FSH_NODYNLNDUSE(time, lndgrid) ;
		FSH_NODYNLNDUSE:long_name = "sensible heat not including correction for land use change" ;
		FSH_NODYNLNDUSE:units = "W/m^2" ;
		FSH_NODYNLNDUSE:cell_methods = "time: mean" ;
		FSH_NODYNLNDUSE:_FillValue = 1.e+36f ;
		FSH_NODYNLNDUSE:missing_value = 1.e+36f ;
	float FSH_R(time, lndgrid) ;
		FSH_R:long_name = "Rural sensible heat" ;
		FSH_R:units = "W/m^2" ;
		FSH_R:cell_methods = "time: mean" ;
		FSH_R:_FillValue = 1.e+36f ;
		FSH_R:missing_value = 1.e+36f ;
	float FSH_U(time, lndgrid) ;
		FSH_U:long_name = "Urban sensible heat" ;
		FSH_U:units = "W/m^2" ;
		FSH_U:cell_methods = "time: mean" ;
		FSH_U:_FillValue = 1.e+36f ;
		FSH_U:missing_value = 1.e+36f ;
	float FSH_V(time, lndgrid) ;
		FSH_V:long_name = "sensible heat from veg" ;
		FSH_V:units = "W/m^2" ;
		FSH_V:cell_methods = "time: mean" ;
		FSH_V:_FillValue = 1.e+36f ;
		FSH_V:missing_value = 1.e+36f ;
	float FSM(time, lndgrid) ;
		FSM:long_name = "snow melt heat flux" ;
		FSM:units = "W/m^2" ;
		FSM:cell_methods = "time: mean" ;
		FSM:_FillValue = 1.e+36f ;
		FSM:missing_value = 1.e+36f ;
	float FSM_R(time, lndgrid) ;
		FSM_R:long_name = "Rural snow melt heat flux" ;
		FSM_R:units = "W/m^2" ;
		FSM_R:cell_methods = "time: mean" ;
		FSM_R:_FillValue = 1.e+36f ;
		FSM_R:missing_value = 1.e+36f ;
	float FSM_U(time, lndgrid) ;
		FSM_U:long_name = "Urban snow melt heat flux" ;
		FSM_U:units = "W/m^2" ;
		FSM_U:cell_methods = "time: mean" ;
		FSM_U:_FillValue = 1.e+36f ;
		FSM_U:missing_value = 1.e+36f ;
	float FSNO(time, lndgrid) ;
		FSNO:long_name = "fraction of ground covered by snow" ;
		FSNO:units = "unitless" ;
		FSNO:cell_methods = "time: mean" ;
		FSNO:_FillValue = 1.e+36f ;
		FSNO:missing_value = 1.e+36f ;
	float FSNO_EFF(time, lndgrid) ;
		FSNO_EFF:long_name = "effective fraction of ground covered by snow" ;
		FSNO_EFF:units = "unitless" ;
		FSNO_EFF:cell_methods = "time: mean" ;
		FSNO_EFF:_FillValue = 1.e+36f ;
		FSNO_EFF:missing_value = 1.e+36f ;
	float FSR(time, lndgrid) ;
		FSR:long_name = "reflected solar radiation" ;
		FSR:units = "W/m^2" ;
		FSR:cell_methods = "time: mean" ;
		FSR:_FillValue = 1.e+36f ;
		FSR:missing_value = 1.e+36f ;
	float FSRND(time, lndgrid) ;
		FSRND:long_name = "direct nir reflected solar radiation" ;
		FSRND:units = "W/m^2" ;
		FSRND:cell_methods = "time: mean" ;
		FSRND:_FillValue = 1.e+36f ;
		FSRND:missing_value = 1.e+36f ;
	float FSRNDLN(time, lndgrid) ;
		FSRNDLN:long_name = "direct nir reflected solar radiation at local noon" ;
		FSRNDLN:units = "W/m^2" ;
		FSRNDLN:cell_methods = "time: mean" ;
		FSRNDLN:_FillValue = 1.e+36f ;
		FSRNDLN:missing_value = 1.e+36f ;
	float FSRNI(time, lndgrid) ;
		FSRNI:long_name = "diffuse nir reflected solar radiation" ;
		FSRNI:units = "W/m^2" ;
		FSRNI:cell_methods = "time: mean" ;
		FSRNI:_FillValue = 1.e+36f ;
		FSRNI:missing_value = 1.e+36f ;
	float FSRVD(time, lndgrid) ;
		FSRVD:long_name = "direct vis reflected solar radiation" ;
		FSRVD:units = "W/m^2" ;
		FSRVD:cell_methods = "time: mean" ;
		FSRVD:_FillValue = 1.e+36f ;
		FSRVD:missing_value = 1.e+36f ;
	float FSRVDLN(time, lndgrid) ;
		FSRVDLN:long_name = "direct vis reflected solar radiation at local noon" ;
		FSRVDLN:units = "W/m^2" ;
		FSRVDLN:cell_methods = "time: mean" ;
		FSRVDLN:_FillValue = 1.e+36f ;
		FSRVDLN:missing_value = 1.e+36f ;
	float FSRVI(time, lndgrid) ;
		FSRVI:long_name = "diffuse vis reflected solar radiation" ;
		FSRVI:units = "W/m^2" ;
		FSRVI:cell_methods = "time: mean" ;
		FSRVI:_FillValue = 1.e+36f ;
		FSRVI:missing_value = 1.e+36f ;
	float FUELC(time, lndgrid) ;
		FUELC:long_name = "fuel load" ;
		FUELC:units = "gC/m^2" ;
		FUELC:cell_methods = "time: mean" ;
		FUELC:_FillValue = 1.e+36f ;
		FUELC:missing_value = 1.e+36f ;
	float F_DENIT(time, lndgrid) ;
		F_DENIT:long_name = "denitrification flux" ;
		F_DENIT:units = "gN/m^2/s" ;
		F_DENIT:cell_methods = "time: mean" ;
		F_DENIT:_FillValue = 1.e+36f ;
		F_DENIT:missing_value = 1.e+36f ;
	float F_DENIT_vr(time, levdcmp, lndgrid) ;
		F_DENIT_vr:long_name = "denitrification flux" ;
		F_DENIT_vr:units = "gN/m^3/s" ;
		F_DENIT_vr:cell_methods = "time: mean" ;
		F_DENIT_vr:_FillValue = 1.e+36f ;
		F_DENIT_vr:missing_value = 1.e+36f ;
	float F_N2O_DENIT(time, lndgrid) ;
		F_N2O_DENIT:long_name = "denitrification N2O flux" ;
		F_N2O_DENIT:units = "gN/m^2/s" ;
		F_N2O_DENIT:cell_methods = "time: mean" ;
		F_N2O_DENIT:_FillValue = 1.e+36f ;
		F_N2O_DENIT:missing_value = 1.e+36f ;
	float F_N2O_NIT(time, lndgrid) ;
		F_N2O_NIT:long_name = "nitrification N2O flux" ;
		F_N2O_NIT:units = "gN/m^2/s" ;
		F_N2O_NIT:cell_methods = "time: mean" ;
		F_N2O_NIT:_FillValue = 1.e+36f ;
		F_N2O_NIT:missing_value = 1.e+36f ;
	float F_NIT(time, lndgrid) ;
		F_NIT:long_name = "nitrification flux" ;
		F_NIT:units = "gN/m^2/s" ;
		F_NIT:cell_methods = "time: mean" ;
		F_NIT:_FillValue = 1.e+36f ;
		F_NIT:missing_value = 1.e+36f ;
	float F_NIT_vr(time, levdcmp, lndgrid) ;
		F_NIT_vr:long_name = "nitrification flux" ;
		F_NIT_vr:units = "gN/m^3/s" ;
		F_NIT_vr:cell_methods = "time: mean" ;
		F_NIT_vr:_FillValue = 1.e+36f ;
		F_NIT_vr:missing_value = 1.e+36f ;
	float GC_HEAT1(time, lndgrid) ;
		GC_HEAT1:long_name = "initial gridcell total heat content" ;
		GC_HEAT1:units = "J/m^2" ;
		GC_HEAT1:cell_methods = "time: mean" ;
		GC_HEAT1:_FillValue = 1.e+36f ;
		GC_HEAT1:missing_value = 1.e+36f ;
	float GC_ICE1(time, lndgrid) ;
		GC_ICE1:long_name = "initial gridcell total ice content" ;
		GC_ICE1:units = "mm" ;
		GC_ICE1:cell_methods = "time: mean" ;
		GC_ICE1:_FillValue = 1.e+36f ;
		GC_ICE1:missing_value = 1.e+36f ;
	float GC_LIQ1(time, lndgrid) ;
		GC_LIQ1:long_name = "initial gridcell total liq content" ;
		GC_LIQ1:units = "mm" ;
		GC_LIQ1:cell_methods = "time: mean" ;
		GC_LIQ1:_FillValue = 1.e+36f ;
		GC_LIQ1:missing_value = 1.e+36f ;
	float GPP(time, lndgrid) ;
		GPP:long_name = "gross primary production" ;
		GPP:units = "gC/m^2/s" ;
		GPP:cell_methods = "time: mean" ;
		GPP:_FillValue = 1.e+36f ;
		GPP:missing_value = 1.e+36f ;
	float GR(time, lndgrid) ;
		GR:long_name = "total growth respiration" ;
		GR:units = "gC/m^2/s" ;
		GR:cell_methods = "time: mean" ;
		GR:_FillValue = 1.e+36f ;
		GR:missing_value = 1.e+36f ;
	float GROSS_NMIN(time, lndgrid) ;
		GROSS_NMIN:long_name = "gross rate of N mineralization" ;
		GROSS_NMIN:units = "gN/m^2/s" ;
		GROSS_NMIN:cell_methods = "time: mean" ;
		GROSS_NMIN:_FillValue = 1.e+36f ;
		GROSS_NMIN:missing_value = 1.e+36f ;
	float H2OCAN(time, lndgrid) ;
		H2OCAN:long_name = "intercepted water" ;
		H2OCAN:units = "mm" ;
		H2OCAN:cell_methods = "time: mean" ;
		H2OCAN:_FillValue = 1.e+36f ;
		H2OCAN:missing_value = 1.e+36f ;
	float H2OSFC(time, lndgrid) ;
		H2OSFC:long_name = "surface water depth" ;
		H2OSFC:units = "mm" ;
		H2OSFC:cell_methods = "time: mean" ;
		H2OSFC:_FillValue = 1.e+36f ;
		H2OSFC:missing_value = 1.e+36f ;
	float H2OSNO(time, lndgrid) ;
		H2OSNO:long_name = "snow depth (liquid water)" ;
		H2OSNO:units = "mm" ;
		H2OSNO:cell_methods = "time: mean" ;
		H2OSNO:_FillValue = 1.e+36f ;
		H2OSNO:missing_value = 1.e+36f ;
	float H2OSNO_TOP(time, lndgrid) ;
		H2OSNO_TOP:long_name = "mass of snow in top snow layer" ;
		H2OSNO_TOP:units = "kg/m2" ;
		H2OSNO_TOP:cell_methods = "time: mean" ;
		H2OSNO_TOP:_FillValue = 1.e+36f ;
		H2OSNO_TOP:missing_value = 1.e+36f ;
	float H2OSOI(time, levgrnd, lndgrid) ;
		H2OSOI:long_name = "volumetric soil water (vegetated landunits only)" ;
		H2OSOI:units = "mm3/mm3" ;
		H2OSOI:cell_methods = "time: mean" ;
		H2OSOI:_FillValue = 1.e+36f ;
		H2OSOI:missing_value = 1.e+36f ;
	float HC(time, lndgrid) ;
		HC:long_name = "heat content of soil/snow/lake" ;
		HC:units = "MJ/m2" ;
		HC:cell_methods = "time: mean" ;
		HC:_FillValue = 1.e+36f ;
		HC:missing_value = 1.e+36f ;
	float HCSOI(time, lndgrid) ;
		HCSOI:long_name = "soil heat content" ;
		HCSOI:units = "MJ/m2" ;
		HCSOI:cell_methods = "time: mean" ;
		HCSOI:_FillValue = 1.e+36f ;
		HCSOI:missing_value = 1.e+36f ;
	float HEAT_FROM_AC(time, lndgrid) ;
		HEAT_FROM_AC:long_name = "sensible heat flux put into canyon due to heat removed from air conditioning" ;
		HEAT_FROM_AC:units = "W/m^2" ;
		HEAT_FROM_AC:cell_methods = "time: mean" ;
		HEAT_FROM_AC:_FillValue = 1.e+36f ;
		HEAT_FROM_AC:missing_value = 1.e+36f ;
	float HR(time, lndgrid) ;
		HR:long_name = "total heterotrophic respiration" ;
		HR:units = "gC/m^2/s" ;
		HR:cell_methods = "time: mean" ;
		HR:_FillValue = 1.e+36f ;
		HR:missing_value = 1.e+36f ;
	float HR_vr(time, levdcmp, lndgrid) ;
		HR_vr:long_name = "total vertically resolved heterotrophic respiration" ;
		HR_vr:units = "gC/m^3/s" ;
		HR_vr:cell_methods = "time: mean" ;
		HR_vr:_FillValue = 1.e+36f ;
		HR_vr:missing_value = 1.e+36f ;
	float HTOP(time, lndgrid) ;
		HTOP:long_name = "canopy top" ;
		HTOP:units = "m" ;
		HTOP:cell_methods = "time: mean" ;
		HTOP:_FillValue = 1.e+36f ;
		HTOP:missing_value = 1.e+36f ;
	float INT_SNOW(time, lndgrid) ;
		INT_SNOW:long_name = "accumulated swe (vegetated landunits only)" ;
		INT_SNOW:units = "mm" ;
		INT_SNOW:cell_methods = "time: mean" ;
		INT_SNOW:_FillValue = 1.e+36f ;
		INT_SNOW:missing_value = 1.e+36f ;
	float LAISHA(time, lndgrid) ;
		LAISHA:long_name = "shaded projected leaf area index" ;
		LAISHA:units = "none" ;
		LAISHA:cell_methods = "time: mean" ;
		LAISHA:_FillValue = 1.e+36f ;
		LAISHA:missing_value = 1.e+36f ;
	float LAISUN(time, lndgrid) ;
		LAISUN:long_name = "sunlit projected leaf area index" ;
		LAISUN:units = "none" ;
		LAISUN:cell_methods = "time: mean" ;
		LAISUN:_FillValue = 1.e+36f ;
		LAISUN:missing_value = 1.e+36f ;
	float LAKEICEFRAC(time, levlak, lndgrid) ;
		LAKEICEFRAC:long_name = "lake layer ice mass fraction" ;
		LAKEICEFRAC:units = "unitless" ;
		LAKEICEFRAC:cell_methods = "time: mean" ;
		LAKEICEFRAC:_FillValue = 1.e+36f ;
		LAKEICEFRAC:missing_value = 1.e+36f ;
	float LAKEICETHICK(time, lndgrid) ;
		LAKEICETHICK:long_name = "thickness of lake ice (including physical expansion on freezing)" ;
		LAKEICETHICK:units = "m" ;
		LAKEICETHICK:cell_methods = "time: mean" ;
		LAKEICETHICK:_FillValue = 1.e+36f ;
		LAKEICETHICK:missing_value = 1.e+36f ;
	float LAND_UPTAKE(time, lndgrid) ;
		LAND_UPTAKE:long_name = "NEE minus LAND_USE_FLUX, negative for update" ;
		LAND_UPTAKE:units = "gC/m^2/s" ;
		LAND_UPTAKE:cell_methods = "time: mean" ;
		LAND_UPTAKE:_FillValue = 1.e+36f ;
		LAND_UPTAKE:missing_value = 1.e+36f ;
	float LAND_USE_FLUX(time, lndgrid) ;
		LAND_USE_FLUX:long_name = "total C emitted from land cover conversion and wood product pools" ;
		LAND_USE_FLUX:units = "gC/m^2/s" ;
		LAND_USE_FLUX:cell_methods = "time: mean" ;
		LAND_USE_FLUX:_FillValue = 1.e+36f ;
		LAND_USE_FLUX:missing_value = 1.e+36f ;
	float LEAFC(time, lndgrid) ;
		LEAFC:long_name = "leaf C" ;
		LEAFC:units = "gC/m^2" ;
		LEAFC:cell_methods = "time: mean" ;
		LEAFC:_FillValue = 1.e+36f ;
		LEAFC:missing_value = 1.e+36f ;
	float LEAFC_ALLOC(time, lndgrid) ;
		LEAFC_ALLOC:long_name = "leaf C allocation" ;
		LEAFC_ALLOC:units = "gC/m^2/s" ;
		LEAFC_ALLOC:cell_methods = "time: mean" ;
		LEAFC_ALLOC:_FillValue = 1.e+36f ;
		LEAFC_ALLOC:missing_value = 1.e+36f ;
	float LEAFC_LOSS(time, lndgrid) ;
		LEAFC_LOSS:long_name = "leaf C loss" ;
		LEAFC_LOSS:units = "gC/m^2/s" ;
		LEAFC_LOSS:cell_methods = "time: mean" ;
		LEAFC_LOSS:_FillValue = 1.e+36f ;
		LEAFC_LOSS:missing_value = 1.e+36f ;
	float LEAFN(time, lndgrid) ;
		LEAFN:long_name = "leaf N" ;
		LEAFN:units = "gN/m^2" ;
		LEAFN:cell_methods = "time: mean" ;
		LEAFN:_FillValue = 1.e+36f ;
		LEAFN:missing_value = 1.e+36f ;
	float LEAF_MR(time, lndgrid) ;
		LEAF_MR:long_name = "leaf maintenance respiration" ;
		LEAF_MR:units = "gC/m^2/s" ;
		LEAF_MR:cell_methods = "time: mean" ;
		LEAF_MR:_FillValue = 1.e+36f ;
		LEAF_MR:missing_value = 1.e+36f ;
	float LFC2(time, lndgrid) ;
		LFC2:long_name = "conversion area fraction of BET and BDT that burned" ;
		LFC2:units = "per sec" ;
		LFC2:cell_methods = "time: mean" ;
		LFC2:_FillValue = 1.e+36f ;
		LFC2:missing_value = 1.e+36f ;
	float LF_CONV_CFLUX(time, lndgrid) ;
		LF_CONV_CFLUX:long_name = "conversion carbon due to BET and BDT area decreasing" ;
		LF_CONV_CFLUX:units = "gC/m^2/s" ;
		LF_CONV_CFLUX:cell_methods = "time: mean" ;
		LF_CONV_CFLUX:_FillValue = 1.e+36f ;
		LF_CONV_CFLUX:missing_value = 1.e+36f ;
	float LITFALL(time, lndgrid) ;
		LITFALL:long_name = "litterfall (leaves and fine roots)" ;
		LITFALL:units = "gC/m^2/s" ;
		LITFALL:cell_methods = "time: mean" ;
		LITFALL:_FillValue = 1.e+36f ;
		LITFALL:missing_value = 1.e+36f ;
	float LITHR(time, lndgrid) ;
		LITHR:long_name = "litter heterotrophic respiration" ;
		LITHR:units = "gC/m^2/s" ;
		LITHR:cell_methods = "time: mean" ;
		LITHR:_FillValue = 1.e+36f ;
		LITHR:missing_value = 1.e+36f ;
	float LITR1C(time, lndgrid) ;
		LITR1C:long_name = "LITR1 C" ;
		LITR1C:units = "gC/m^2" ;
		LITR1C:cell_methods = "time: mean" ;
		LITR1C:_FillValue = 1.e+36f ;
		LITR1C:missing_value = 1.e+36f ;
	float LITR1C_TO_SOIL1C(time, lndgrid) ;
		LITR1C_TO_SOIL1C:long_name = "decomp. of litter 1 C to soil 1 C" ;
		LITR1C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR1C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR1C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR1C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR1C_vr(time, levdcmp, lndgrid) ;
		LITR1C_vr:long_name = "LITR1 C (vertically resolved)" ;
		LITR1C_vr:units = "gC/m^3" ;
		LITR1C_vr:cell_methods = "time: mean" ;
		LITR1C_vr:_FillValue = 1.e+36f ;
		LITR1C_vr:missing_value = 1.e+36f ;
	float LITR1N(time, lndgrid) ;
		LITR1N:long_name = "LITR1 N" ;
		LITR1N:units = "gN/m^2" ;
		LITR1N:cell_methods = "time: mean" ;
		LITR1N:_FillValue = 1.e+36f ;
		LITR1N:missing_value = 1.e+36f ;
	float LITR1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR1N_TNDNCY_VERT_TRANS:long_name = "litter 1 N tendency due to vertical transport" ;
		LITR1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR1N_TO_SOIL1N(time, lndgrid) ;
		LITR1N_TO_SOIL1N:long_name = "decomp. of litter 1 N to soil 1 N" ;
		LITR1N_TO_SOIL1N:units = "gN/m^2" ;
		LITR1N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR1N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR1N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR1N_vr(time, levdcmp, lndgrid) ;
		LITR1N_vr:long_name = "LITR1 N (vertically resolved)" ;
		LITR1N_vr:units = "gN/m^3" ;
		LITR1N_vr:cell_methods = "time: mean" ;
		LITR1N_vr:_FillValue = 1.e+36f ;
		LITR1N_vr:missing_value = 1.e+36f ;
	float LITR1_HR(time, lndgrid) ;
		LITR1_HR:long_name = "Het. Resp. from litter 1" ;
		LITR1_HR:units = "gC/m^2/s" ;
		LITR1_HR:cell_methods = "time: mean" ;
		LITR1_HR:_FillValue = 1.e+36f ;
		LITR1_HR:missing_value = 1.e+36f ;
	float LITR2C(time, lndgrid) ;
		LITR2C:long_name = "LITR2 C" ;
		LITR2C:units = "gC/m^2" ;
		LITR2C:cell_methods = "time: mean" ;
		LITR2C:_FillValue = 1.e+36f ;
		LITR2C:missing_value = 1.e+36f ;
	float LITR2C_TO_SOIL1C(time, lndgrid) ;
		LITR2C_TO_SOIL1C:long_name = "decomp. of litter 2 C to soil 1 C" ;
		LITR2C_TO_SOIL1C:units = "gC/m^2/s" ;
		LITR2C_TO_SOIL1C:cell_methods = "time: mean" ;
		LITR2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		LITR2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float LITR2C_vr(time, levdcmp, lndgrid) ;
		LITR2C_vr:long_name = "LITR2 C (vertically resolved)" ;
		LITR2C_vr:units = "gC/m^3" ;
		LITR2C_vr:cell_methods = "time: mean" ;
		LITR2C_vr:_FillValue = 1.e+36f ;
		LITR2C_vr:missing_value = 1.e+36f ;
	float LITR2N(time, lndgrid) ;
		LITR2N:long_name = "LITR2 N" ;
		LITR2N:units = "gN/m^2" ;
		LITR2N:cell_methods = "time: mean" ;
		LITR2N:_FillValue = 1.e+36f ;
		LITR2N:missing_value = 1.e+36f ;
	float LITR2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR2N_TNDNCY_VERT_TRANS:long_name = "litter 2 N tendency due to vertical transport" ;
		LITR2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR2N_TO_SOIL1N(time, lndgrid) ;
		LITR2N_TO_SOIL1N:long_name = "decomp. of litter 2 N to soil 1 N" ;
		LITR2N_TO_SOIL1N:units = "gN/m^2" ;
		LITR2N_TO_SOIL1N:cell_methods = "time: mean" ;
		LITR2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		LITR2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float LITR2N_vr(time, levdcmp, lndgrid) ;
		LITR2N_vr:long_name = "LITR2 N (vertically resolved)" ;
		LITR2N_vr:units = "gN/m^3" ;
		LITR2N_vr:cell_methods = "time: mean" ;
		LITR2N_vr:_FillValue = 1.e+36f ;
		LITR2N_vr:missing_value = 1.e+36f ;
	float LITR2_HR(time, lndgrid) ;
		LITR2_HR:long_name = "Het. Resp. from litter 2" ;
		LITR2_HR:units = "gC/m^2/s" ;
		LITR2_HR:cell_methods = "time: mean" ;
		LITR2_HR:_FillValue = 1.e+36f ;
		LITR2_HR:missing_value = 1.e+36f ;
	float LITR3C(time, lndgrid) ;
		LITR3C:long_name = "LITR3 C" ;
		LITR3C:units = "gC/m^2" ;
		LITR3C:cell_methods = "time: mean" ;
		LITR3C:_FillValue = 1.e+36f ;
		LITR3C:missing_value = 1.e+36f ;
	float LITR3C_TO_SOIL2C(time, lndgrid) ;
		LITR3C_TO_SOIL2C:long_name = "decomp. of litter 3 C to soil 2 C" ;
		LITR3C_TO_SOIL2C:units = "gC/m^2/s" ;
		LITR3C_TO_SOIL2C:cell_methods = "time: mean" ;
		LITR3C_TO_SOIL2C:_FillValue = 1.e+36f ;
		LITR3C_TO_SOIL2C:missing_value = 1.e+36f ;
	float LITR3C_vr(time, levdcmp, lndgrid) ;
		LITR3C_vr:long_name = "LITR3 C (vertically resolved)" ;
		LITR3C_vr:units = "gC/m^3" ;
		LITR3C_vr:cell_methods = "time: mean" ;
		LITR3C_vr:_FillValue = 1.e+36f ;
		LITR3C_vr:missing_value = 1.e+36f ;
	float LITR3N(time, lndgrid) ;
		LITR3N:long_name = "LITR3 N" ;
		LITR3N:units = "gN/m^2" ;
		LITR3N:cell_methods = "time: mean" ;
		LITR3N:_FillValue = 1.e+36f ;
		LITR3N:missing_value = 1.e+36f ;
	float LITR3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		LITR3N_TNDNCY_VERT_TRANS:long_name = "litter 3 N tendency due to vertical transport" ;
		LITR3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		LITR3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		LITR3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		LITR3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float LITR3N_TO_SOIL2N(time, lndgrid) ;
		LITR3N_TO_SOIL2N:long_name = "decomp. of litter 3 N to soil 2 N" ;
		LITR3N_TO_SOIL2N:units = "gN/m^2" ;
		LITR3N_TO_SOIL2N:cell_methods = "time: mean" ;
		LITR3N_TO_SOIL2N:_FillValue = 1.e+36f ;
		LITR3N_TO_SOIL2N:missing_value = 1.e+36f ;
	float LITR3N_vr(time, levdcmp, lndgrid) ;
		LITR3N_vr:long_name = "LITR3 N (vertically resolved)" ;
		LITR3N_vr:units = "gN/m^3" ;
		LITR3N_vr:cell_methods = "time: mean" ;
		LITR3N_vr:_FillValue = 1.e+36f ;
		LITR3N_vr:missing_value = 1.e+36f ;
	float LITR3_HR(time, lndgrid) ;
		LITR3_HR:long_name = "Het. Resp. from litter 3" ;
		LITR3_HR:units = "gC/m^2/s" ;
		LITR3_HR:cell_methods = "time: mean" ;
		LITR3_HR:_FillValue = 1.e+36f ;
		LITR3_HR:missing_value = 1.e+36f ;
	float LITTERC(time, lndgrid) ;
		LITTERC:long_name = "litter C" ;
		LITTERC:units = "gC/m^2" ;
		LITTERC:cell_methods = "time: mean" ;
		LITTERC:_FillValue = 1.e+36f ;
		LITTERC:missing_value = 1.e+36f ;
	float LITTERC_HR(time, lndgrid) ;
		LITTERC_HR:long_name = "litter C heterotrophic respiration" ;
		LITTERC_HR:units = "gC/m^2/s" ;
		LITTERC_HR:cell_methods = "time: mean" ;
		LITTERC_HR:_FillValue = 1.e+36f ;
		LITTERC_HR:missing_value = 1.e+36f ;
	float LITTERC_LOSS(time, lndgrid) ;
		LITTERC_LOSS:long_name = "litter C loss" ;
		LITTERC_LOSS:units = "gC/m^2/s" ;
		LITTERC_LOSS:cell_methods = "time: mean" ;
		LITTERC_LOSS:_FillValue = 1.e+36f ;
		LITTERC_LOSS:missing_value = 1.e+36f ;
	float LIVECROOTC(time, lndgrid) ;
		LIVECROOTC:long_name = "live coarse root C" ;
		LIVECROOTC:units = "gC/m^2" ;
		LIVECROOTC:cell_methods = "time: mean" ;
		LIVECROOTC:_FillValue = 1.e+36f ;
		LIVECROOTC:missing_value = 1.e+36f ;
	float LIVECROOTN(time, lndgrid) ;
		LIVECROOTN:long_name = "live coarse root N" ;
		LIVECROOTN:units = "gN/m^2" ;
		LIVECROOTN:cell_methods = "time: mean" ;
		LIVECROOTN:_FillValue = 1.e+36f ;
		LIVECROOTN:missing_value = 1.e+36f ;
	float LIVESTEMC(time, lndgrid) ;
		LIVESTEMC:long_name = "live stem C" ;
		LIVESTEMC:units = "gC/m^2" ;
		LIVESTEMC:cell_methods = "time: mean" ;
		LIVESTEMC:_FillValue = 1.e+36f ;
		LIVESTEMC:missing_value = 1.e+36f ;
	float LIVESTEMN(time, lndgrid) ;
		LIVESTEMN:long_name = "live stem N" ;
		LIVESTEMN:units = "gN/m^2" ;
		LIVESTEMN:cell_methods = "time: mean" ;
		LIVESTEMN:_FillValue = 1.e+36f ;
		LIVESTEMN:missing_value = 1.e+36f ;
	float MEG_acetaldehyde(time, lndgrid) ;
		MEG_acetaldehyde:long_name = "MEGAN flux" ;
		MEG_acetaldehyde:units = "kg/m2/sec" ;
		MEG_acetaldehyde:cell_methods = "time: mean" ;
		MEG_acetaldehyde:_FillValue = 1.e+36f ;
		MEG_acetaldehyde:missing_value = 1.e+36f ;
	float MEG_acetic_acid(time, lndgrid) ;
		MEG_acetic_acid:long_name = "MEGAN flux" ;
		MEG_acetic_acid:units = "kg/m2/sec" ;
		MEG_acetic_acid:cell_methods = "time: mean" ;
		MEG_acetic_acid:_FillValue = 1.e+36f ;
		MEG_acetic_acid:missing_value = 1.e+36f ;
	float MEG_acetone(time, lndgrid) ;
		MEG_acetone:long_name = "MEGAN flux" ;
		MEG_acetone:units = "kg/m2/sec" ;
		MEG_acetone:cell_methods = "time: mean" ;
		MEG_acetone:_FillValue = 1.e+36f ;
		MEG_acetone:missing_value = 1.e+36f ;
	float MEG_carene_3(time, lndgrid) ;
		MEG_carene_3:long_name = "MEGAN flux" ;
		MEG_carene_3:units = "kg/m2/sec" ;
		MEG_carene_3:cell_methods = "time: mean" ;
		MEG_carene_3:_FillValue = 1.e+36f ;
		MEG_carene_3:missing_value = 1.e+36f ;
	float MEG_ethanol(time, lndgrid) ;
		MEG_ethanol:long_name = "MEGAN flux" ;
		MEG_ethanol:units = "kg/m2/sec" ;
		MEG_ethanol:cell_methods = "time: mean" ;
		MEG_ethanol:_FillValue = 1.e+36f ;
		MEG_ethanol:missing_value = 1.e+36f ;
	float MEG_formaldehyde(time, lndgrid) ;
		MEG_formaldehyde:long_name = "MEGAN flux" ;
		MEG_formaldehyde:units = "kg/m2/sec" ;
		MEG_formaldehyde:cell_methods = "time: mean" ;
		MEG_formaldehyde:_FillValue = 1.e+36f ;
		MEG_formaldehyde:missing_value = 1.e+36f ;
	float MEG_isoprene(time, lndgrid) ;
		MEG_isoprene:long_name = "MEGAN flux" ;
		MEG_isoprene:units = "kg/m2/sec" ;
		MEG_isoprene:cell_methods = "time: mean" ;
		MEG_isoprene:_FillValue = 1.e+36f ;
		MEG_isoprene:missing_value = 1.e+36f ;
	float MEG_methanol(time, lndgrid) ;
		MEG_methanol:long_name = "MEGAN flux" ;
		MEG_methanol:units = "kg/m2/sec" ;
		MEG_methanol:cell_methods = "time: mean" ;
		MEG_methanol:_FillValue = 1.e+36f ;
		MEG_methanol:missing_value = 1.e+36f ;
	float MEG_pinene_a(time, lndgrid) ;
		MEG_pinene_a:long_name = "MEGAN flux" ;
		MEG_pinene_a:units = "kg/m2/sec" ;
		MEG_pinene_a:cell_methods = "time: mean" ;
		MEG_pinene_a:_FillValue = 1.e+36f ;
		MEG_pinene_a:missing_value = 1.e+36f ;
	float MEG_thujene_a(time, lndgrid) ;
		MEG_thujene_a:long_name = "MEGAN flux" ;
		MEG_thujene_a:units = "kg/m2/sec" ;
		MEG_thujene_a:cell_methods = "time: mean" ;
		MEG_thujene_a:_FillValue = 1.e+36f ;
		MEG_thujene_a:missing_value = 1.e+36f ;
	float MR(time, lndgrid) ;
		MR:long_name = "maintenance respiration" ;
		MR:units = "gC/m^2/s" ;
		MR:cell_methods = "time: mean" ;
		MR:_FillValue = 1.e+36f ;
		MR:missing_value = 1.e+36f ;
	float M_LITR1C_TO_LEACHING(time, lndgrid) ;
		M_LITR1C_TO_LEACHING:long_name = "litter 1 C leaching loss" ;
		M_LITR1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR2C_TO_LEACHING(time, lndgrid) ;
		M_LITR2C_TO_LEACHING:long_name = "litter 2 C leaching loss" ;
		M_LITR2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_LITR3C_TO_LEACHING(time, lndgrid) ;
		M_LITR3C_TO_LEACHING:long_name = "litter 3 C leaching loss" ;
		M_LITR3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_LITR3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_LITR3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_LITR3C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL1C_TO_LEACHING(time, lndgrid) ;
		M_SOIL1C_TO_LEACHING:long_name = "soil 1 C leaching loss" ;
		M_SOIL1C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL1C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL1C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL1C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL2C_TO_LEACHING(time, lndgrid) ;
		M_SOIL2C_TO_LEACHING:long_name = "soil 2 C leaching loss" ;
		M_SOIL2C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL2C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL2C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL2C_TO_LEACHING:missing_value = 1.e+36f ;
	float M_SOIL3C_TO_LEACHING(time, lndgrid) ;
		M_SOIL3C_TO_LEACHING:long_name = "soil 3 C leaching loss" ;
		M_SOIL3C_TO_LEACHING:units = "gC/m^2/s" ;
		M_SOIL3C_TO_LEACHING:cell_methods = "time: mean" ;
		M_SOIL3C_TO_LEACHING:_FillValue = 1.e+36f ;
		M_SOIL3C_TO_LEACHING:missing_value = 1.e+36f ;
	float NBP(time, lndgrid) ;
		NBP:long_name = "net biome production, includes fire, landuse, and harvest flux, positive for sink" ;
		NBP:units = "gC/m^2/s" ;
		NBP:cell_methods = "time: mean" ;
		NBP:_FillValue = 1.e+36f ;
		NBP:missing_value = 1.e+36f ;
	float NDEPLOY(time, lndgrid) ;
		NDEPLOY:long_name = "total N deployed in new growth" ;
		NDEPLOY:units = "gN/m^2/s" ;
		NDEPLOY:cell_methods = "time: mean" ;
		NDEPLOY:_FillValue = 1.e+36f ;
		NDEPLOY:missing_value = 1.e+36f ;
	float NDEP_TO_SMINN(time, lndgrid) ;
		NDEP_TO_SMINN:long_name = "atmospheric N deposition to soil mineral N" ;
		NDEP_TO_SMINN:units = "gN/m^2/s" ;
		NDEP_TO_SMINN:cell_methods = "time: mean" ;
		NDEP_TO_SMINN:_FillValue = 1.e+36f ;
		NDEP_TO_SMINN:missing_value = 1.e+36f ;
	float NEE(time, lndgrid) ;
		NEE:long_name = "net ecosystem exchange of carbon, includes fire, landuse, harvest, and hrv_xsmrpool flux, positive for source" ;
		NEE:units = "gC/m^2/s" ;
		NEE:cell_methods = "time: mean" ;
		NEE:_FillValue = 1.e+36f ;
		NEE:missing_value = 1.e+36f ;
	float NEM(time, lndgrid) ;
		NEM:long_name = "Gridcell net adjustment to NEE passed to atm. for methane production" ;
		NEM:units = "gC/m2/s" ;
		NEM:cell_methods = "time: mean" ;
		NEM:_FillValue = 1.e+36f ;
		NEM:missing_value = 1.e+36f ;
	float NEP(time, lndgrid) ;
		NEP:long_name = "net ecosystem production, excludes fire, landuse, and harvest flux, positive for sink" ;
		NEP:units = "gC/m^2/s" ;
		NEP:cell_methods = "time: mean" ;
		NEP:_FillValue = 1.e+36f ;
		NEP:missing_value = 1.e+36f ;
	float NET_NMIN(time, lndgrid) ;
		NET_NMIN:long_name = "net rate of N mineralization" ;
		NET_NMIN:units = "gN/m^2/s" ;
		NET_NMIN:cell_methods = "time: mean" ;
		NET_NMIN:_FillValue = 1.e+36f ;
		NET_NMIN:missing_value = 1.e+36f ;
	float NFIRE(time, lndgrid) ;
		NFIRE:long_name = "fire counts valid only in Reg.C" ;
		NFIRE:units = "counts/km2/sec" ;
		NFIRE:cell_methods = "time: mean" ;
		NFIRE:_FillValue = 1.e+36f ;
		NFIRE:missing_value = 1.e+36f ;
	float NFIX_TO_SMINN(time, lndgrid) ;
		NFIX_TO_SMINN:long_name = "symbiotic/asymbiotic N fixation to soil mineral N" ;
		NFIX_TO_SMINN:units = "gN/m^2/s" ;
		NFIX_TO_SMINN:cell_methods = "time: mean" ;
		NFIX_TO_SMINN:_FillValue = 1.e+36f ;
		NFIX_TO_SMINN:missing_value = 1.e+36f ;
	float NPP(time, lndgrid) ;
		NPP:long_name = "net primary production" ;
		NPP:units = "gC/m^2/s" ;
		NPP:cell_methods = "time: mean" ;
		NPP:_FillValue = 1.e+36f ;
		NPP:missing_value = 1.e+36f ;
	float OCDEP(time, lndgrid) ;
		OCDEP:long_name = "total OC deposition (dry+wet) from atmosphere" ;
		OCDEP:units = "kg/m^2/s" ;
		OCDEP:cell_methods = "time: mean" ;
		OCDEP:_FillValue = 1.e+36f ;
		OCDEP:missing_value = 1.e+36f ;
	float O_SCALAR(time, levdcmp, lndgrid) ;
		O_SCALAR:long_name = "fraction by which decomposition is reduced due to anoxia" ;
		O_SCALAR:units = "unitless" ;
		O_SCALAR:cell_methods = "time: mean" ;
		O_SCALAR:_FillValue = 1.e+36f ;
		O_SCALAR:missing_value = 1.e+36f ;
	float PARVEGLN(time, lndgrid) ;
		PARVEGLN:long_name = "absorbed par by vegetation at local noon" ;
		PARVEGLN:units = "W/m^2" ;
		PARVEGLN:cell_methods = "time: mean" ;
		PARVEGLN:_FillValue = 1.e+36f ;
		PARVEGLN:missing_value = 1.e+36f ;
	float PBOT(time, lndgrid) ;
		PBOT:long_name = "atmospheric pressure" ;
		PBOT:units = "Pa" ;
		PBOT:cell_methods = "time: mean" ;
		PBOT:_FillValue = 1.e+36f ;
		PBOT:missing_value = 1.e+36f ;
	float PCH4(time, lndgrid) ;
		PCH4:long_name = "atmospheric partial pressure of CH4" ;
		PCH4:units = "Pa" ;
		PCH4:cell_methods = "time: mean" ;
		PCH4:_FillValue = 1.e+36f ;
		PCH4:missing_value = 1.e+36f ;
	float PCO2(time, lndgrid) ;
		PCO2:long_name = "atmospheric partial pressure of CO2" ;
		PCO2:units = "Pa" ;
		PCO2:cell_methods = "time: mean" ;
		PCO2:_FillValue = 1.e+36f ;
		PCO2:missing_value = 1.e+36f ;
	float PCT_LANDUNIT(time, ltype, lndgrid) ;
		PCT_LANDUNIT:long_name = "% of each landunit on grid cell" ;
		PCT_LANDUNIT:units = "%" ;
		PCT_LANDUNIT:cell_methods = "time: mean" ;
		PCT_LANDUNIT:_FillValue = 1.e+36f ;
		PCT_LANDUNIT:missing_value = 1.e+36f ;
	float PCT_NAT_PFT(time, natpft, lndgrid) ;
		PCT_NAT_PFT:long_name = "% of each PFT on the natural vegetation (i.e., soil) landunit" ;
		PCT_NAT_PFT:units = "%" ;
		PCT_NAT_PFT:cell_methods = "time: mean" ;
		PCT_NAT_PFT:_FillValue = 1.e+36f ;
		PCT_NAT_PFT:missing_value = 1.e+36f ;
	float PFT_CTRUNC(time, lndgrid) ;
		PFT_CTRUNC:long_name = "pft-level sink for C truncation" ;
		PFT_CTRUNC:units = "gC/m^2" ;
		PFT_CTRUNC:cell_methods = "time: mean" ;
		PFT_CTRUNC:_FillValue = 1.e+36f ;
		PFT_CTRUNC:missing_value = 1.e+36f ;
	float PFT_FIRE_CLOSS(time, lndgrid) ;
		PFT_FIRE_CLOSS:long_name = "total pft-level fire C loss for non-peat fires outside land-type converted region" ;
		PFT_FIRE_CLOSS:units = "gC/m^2/s" ;
		PFT_FIRE_CLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_CLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_CLOSS:missing_value = 1.e+36f ;
	float PFT_FIRE_NLOSS(time, lndgrid) ;
		PFT_FIRE_NLOSS:long_name = "total pft-level fire N loss" ;
		PFT_FIRE_NLOSS:units = "gN/m^2/s" ;
		PFT_FIRE_NLOSS:cell_methods = "time: mean" ;
		PFT_FIRE_NLOSS:_FillValue = 1.e+36f ;
		PFT_FIRE_NLOSS:missing_value = 1.e+36f ;
	float PFT_NTRUNC(time, lndgrid) ;
		PFT_NTRUNC:long_name = "pft-level sink for N truncation" ;
		PFT_NTRUNC:units = "gN/m^2" ;
		PFT_NTRUNC:cell_methods = "time: mean" ;
		PFT_NTRUNC:_FillValue = 1.e+36f ;
		PFT_NTRUNC:missing_value = 1.e+36f ;
	float PLANT_NDEMAND(time, lndgrid) ;
		PLANT_NDEMAND:long_name = "N flux required to support initial GPP" ;
		PLANT_NDEMAND:units = "gN/m^2/s" ;
		PLANT_NDEMAND:cell_methods = "time: mean" ;
		PLANT_NDEMAND:_FillValue = 1.e+36f ;
		PLANT_NDEMAND:missing_value = 1.e+36f ;
	float POTENTIAL_IMMOB(time, lndgrid) ;
		POTENTIAL_IMMOB:long_name = "potential N immobilization" ;
		POTENTIAL_IMMOB:units = "gN/m^2/s" ;
		POTENTIAL_IMMOB:cell_methods = "time: mean" ;
		POTENTIAL_IMMOB:_FillValue = 1.e+36f ;
		POTENTIAL_IMMOB:missing_value = 1.e+36f ;
	float POT_F_DENIT(time, lndgrid) ;
		POT_F_DENIT:long_name = "potential denitrification flux" ;
		POT_F_DENIT:units = "gN/m^2/s" ;
		POT_F_DENIT:cell_methods = "time: mean" ;
		POT_F_DENIT:_FillValue = 1.e+36f ;
		POT_F_DENIT:missing_value = 1.e+36f ;
	float POT_F_NIT(time, lndgrid) ;
		POT_F_NIT:long_name = "potential nitrification flux" ;
		POT_F_NIT:units = "gN/m^2/s" ;
		POT_F_NIT:cell_methods = "time: mean" ;
		POT_F_NIT:_FillValue = 1.e+36f ;
		POT_F_NIT:missing_value = 1.e+36f ;
	float PROD100C(time, lndgrid) ;
		PROD100C:long_name = "100-yr wood product C" ;
		PROD100C:units = "gC/m^2" ;
		PROD100C:cell_methods = "time: mean" ;
		PROD100C:_FillValue = 1.e+36f ;
		PROD100C:missing_value = 1.e+36f ;
	float PROD100C_LOSS(time, lndgrid) ;
		PROD100C_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100C_LOSS:units = "gC/m^2/s" ;
		PROD100C_LOSS:cell_methods = "time: mean" ;
		PROD100C_LOSS:_FillValue = 1.e+36f ;
		PROD100C_LOSS:missing_value = 1.e+36f ;
	float PROD100N(time, lndgrid) ;
		PROD100N:long_name = "100-yr wood product N" ;
		PROD100N:units = "gN/m^2" ;
		PROD100N:cell_methods = "time: mean" ;
		PROD100N:_FillValue = 1.e+36f ;
		PROD100N:missing_value = 1.e+36f ;
	float PROD100N_LOSS(time, lndgrid) ;
		PROD100N_LOSS:long_name = "loss from 100-yr wood product pool" ;
		PROD100N_LOSS:units = "gN/m^2/s" ;
		PROD100N_LOSS:cell_methods = "time: mean" ;
		PROD100N_LOSS:_FillValue = 1.e+36f ;
		PROD100N_LOSS:missing_value = 1.e+36f ;
	float PROD10C(time, lndgrid) ;
		PROD10C:long_name = "10-yr wood product C" ;
		PROD10C:units = "gC/m^2" ;
		PROD10C:cell_methods = "time: mean" ;
		PROD10C:_FillValue = 1.e+36f ;
		PROD10C:missing_value = 1.e+36f ;
	float PROD10C_LOSS(time, lndgrid) ;
		PROD10C_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10C_LOSS:units = "gC/m^2/s" ;
		PROD10C_LOSS:cell_methods = "time: mean" ;
		PROD10C_LOSS:_FillValue = 1.e+36f ;
		PROD10C_LOSS:missing_value = 1.e+36f ;
	float PROD10N(time, lndgrid) ;
		PROD10N:long_name = "10-yr wood product N" ;
		PROD10N:units = "gN/m^2" ;
		PROD10N:cell_methods = "time: mean" ;
		PROD10N:_FillValue = 1.e+36f ;
		PROD10N:missing_value = 1.e+36f ;
	float PROD10N_LOSS(time, lndgrid) ;
		PROD10N_LOSS:long_name = "loss from 10-yr wood product pool" ;
		PROD10N_LOSS:units = "gN/m^2/s" ;
		PROD10N_LOSS:cell_methods = "time: mean" ;
		PROD10N_LOSS:_FillValue = 1.e+36f ;
		PROD10N_LOSS:missing_value = 1.e+36f ;
	float PRODUCT_CLOSS(time, lndgrid) ;
		PRODUCT_CLOSS:long_name = "total carbon loss from wood product pools" ;
		PRODUCT_CLOSS:units = "gC/m^2/s" ;
		PRODUCT_CLOSS:cell_methods = "time: mean" ;
		PRODUCT_CLOSS:_FillValue = 1.e+36f ;
		PRODUCT_CLOSS:missing_value = 1.e+36f ;
	float PRODUCT_NLOSS(time, lndgrid) ;
		PRODUCT_NLOSS:long_name = "total N loss from wood product pools" ;
		PRODUCT_NLOSS:units = "gN/m^2/s" ;
		PRODUCT_NLOSS:cell_methods = "time: mean" ;
		PRODUCT_NLOSS:_FillValue = 1.e+36f ;
		PRODUCT_NLOSS:missing_value = 1.e+36f ;
	float PSNSHA(time, lndgrid) ;
		PSNSHA:long_name = "shaded leaf photosynthesis" ;
		PSNSHA:units = "umolCO2/m^2/s" ;
		PSNSHA:cell_methods = "time: mean" ;
		PSNSHA:_FillValue = 1.e+36f ;
		PSNSHA:missing_value = 1.e+36f ;
	float PSNSHADE_TO_CPOOL(time, lndgrid) ;
		PSNSHADE_TO_CPOOL:long_name = "C fixation from shaded canopy" ;
		PSNSHADE_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSHADE_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSHADE_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSHADE_TO_CPOOL:missing_value = 1.e+36f ;
	float PSNSUN(time, lndgrid) ;
		PSNSUN:long_name = "sunlit leaf photosynthesis" ;
		PSNSUN:units = "umolCO2/m^2/s" ;
		PSNSUN:cell_methods = "time: mean" ;
		PSNSUN:_FillValue = 1.e+36f ;
		PSNSUN:missing_value = 1.e+36f ;
	float PSNSUN_TO_CPOOL(time, lndgrid) ;
		PSNSUN_TO_CPOOL:long_name = "C fixation from sunlit canopy" ;
		PSNSUN_TO_CPOOL:units = "gC/m^2/s" ;
		PSNSUN_TO_CPOOL:cell_methods = "time: mean" ;
		PSNSUN_TO_CPOOL:_FillValue = 1.e+36f ;
		PSNSUN_TO_CPOOL:missing_value = 1.e+36f ;
	float Q2M(time, lndgrid) ;
		Q2M:long_name = "2m specific humidity" ;
		Q2M:units = "kg/kg" ;
		Q2M:cell_methods = "time: mean" ;
		Q2M:_FillValue = 1.e+36f ;
		Q2M:missing_value = 1.e+36f ;
	float QBOT(time, lndgrid) ;
		QBOT:long_name = "atmospheric specific humidity" ;
		QBOT:units = "kg/kg" ;
		QBOT:cell_methods = "time: mean" ;
		QBOT:_FillValue = 1.e+36f ;
		QBOT:missing_value = 1.e+36f ;
	float QCHARGE(time, lndgrid) ;
		QCHARGE:long_name = "aquifer recharge rate (vegetated landunits only)" ;
		QCHARGE:units = "mm/s" ;
		QCHARGE:cell_methods = "time: mean" ;
		QCHARGE:_FillValue = 1.e+36f ;
		QCHARGE:missing_value = 1.e+36f ;
	float QDRAI(time, lndgrid) ;
		QDRAI:long_name = "sub-surface drainage" ;
		QDRAI:units = "mm/s" ;
		QDRAI:cell_methods = "time: mean" ;
		QDRAI:_FillValue = 1.e+36f ;
		QDRAI:missing_value = 1.e+36f ;
	float QDRAI_PERCH(time, lndgrid) ;
		QDRAI_PERCH:long_name = "perched wt drainage" ;
		QDRAI_PERCH:units = "mm/s" ;
		QDRAI_PERCH:cell_methods = "time: mean" ;
		QDRAI_PERCH:_FillValue = 1.e+36f ;
		QDRAI_PERCH:missing_value = 1.e+36f ;
	float QDRAI_XS(time, lndgrid) ;
		QDRAI_XS:long_name = "saturation excess drainage" ;
		QDRAI_XS:units = "mm/s" ;
		QDRAI_XS:cell_methods = "time: mean" ;
		QDRAI_XS:_FillValue = 1.e+36f ;
		QDRAI_XS:missing_value = 1.e+36f ;
	float QDRIP(time, lndgrid) ;
		QDRIP:long_name = "throughfall" ;
		QDRIP:units = "mm/s" ;
		QDRIP:cell_methods = "time: mean" ;
		QDRIP:_FillValue = 1.e+36f ;
		QDRIP:missing_value = 1.e+36f ;
	float QFLOOD(time, lndgrid) ;
		QFLOOD:long_name = "runoff from river flooding" ;
		QFLOOD:units = "mm/s" ;
		QFLOOD:cell_methods = "time: mean" ;
		QFLOOD:_FillValue = 1.e+36f ;
		QFLOOD:missing_value = 1.e+36f ;
	float QFLX_ICE_DYNBAL(time, lndgrid) ;
		QFLX_ICE_DYNBAL:long_name = "ice dynamic land cover change conversion runoff flux" ;
		QFLX_ICE_DYNBAL:units = "mm/s" ;
		QFLX_ICE_DYNBAL:cell_methods = "time: mean" ;
		QFLX_ICE_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_ICE_DYNBAL:missing_value = 1.e+36f ;
	float QFLX_LIQ_DYNBAL(time, lndgrid) ;
		QFLX_LIQ_DYNBAL:long_name = "liq dynamic land cover change conversion runoff flux" ;
		QFLX_LIQ_DYNBAL:units = "mm/s" ;
		QFLX_LIQ_DYNBAL:cell_methods = "time: mean" ;
		QFLX_LIQ_DYNBAL:_FillValue = 1.e+36f ;
		QFLX_LIQ_DYNBAL:missing_value = 1.e+36f ;
	float QH2OSFC(time, lndgrid) ;
		QH2OSFC:long_name = "surface water runoff" ;
		QH2OSFC:units = "mm/s" ;
		QH2OSFC:cell_methods = "time: mean" ;
		QH2OSFC:_FillValue = 1.e+36f ;
		QH2OSFC:missing_value = 1.e+36f ;
	float QINFL(time, lndgrid) ;
		QINFL:long_name = "infiltration" ;
		QINFL:units = "mm/s" ;
		QINFL:cell_methods = "time: mean" ;
		QINFL:_FillValue = 1.e+36f ;
		QINFL:missing_value = 1.e+36f ;
	float QINTR(time, lndgrid) ;
		QINTR:long_name = "interception" ;
		QINTR:units = "mm/s" ;
		QINTR:cell_methods = "time: mean" ;
		QINTR:_FillValue = 1.e+36f ;
		QINTR:missing_value = 1.e+36f ;
	float QIRRIG(time, lndgrid) ;
		QIRRIG:long_name = "water added through irrigation" ;
		QIRRIG:units = "mm/s" ;
		QIRRIG:cell_methods = "time: mean" ;
		QIRRIG:_FillValue = 1.e+36f ;
		QIRRIG:missing_value = 1.e+36f ;
	float QOVER(time, lndgrid) ;
		QOVER:long_name = "surface runoff" ;
		QOVER:units = "mm/s" ;
		QOVER:cell_methods = "time: mean" ;
		QOVER:_FillValue = 1.e+36f ;
		QOVER:missing_value = 1.e+36f ;
	float QOVER_LAG(time, lndgrid) ;
		QOVER_LAG:long_name = "time-lagged surface runoff for soil columns" ;
		QOVER_LAG:units = "mm/s" ;
		QOVER_LAG:cell_methods = "time: mean" ;
		QOVER_LAG:_FillValue = 1.e+36f ;
		QOVER_LAG:missing_value = 1.e+36f ;
	float QRGWL(time, lndgrid) ;
		QRGWL:long_name = "surface runoff at glaciers (liquid only), wetlands, lakes" ;
		QRGWL:units = "mm/s" ;
		QRGWL:cell_methods = "time: mean" ;
		QRGWL:_FillValue = 1.e+36f ;
		QRGWL:missing_value = 1.e+36f ;
	float QRUNOFF(time, lndgrid) ;
		QRUNOFF:long_name = "total liquid runoff (does not include QSNWCPICE)" ;
		QRUNOFF:units = "mm/s" ;
		QRUNOFF:cell_methods = "time: mean" ;
		QRUNOFF:_FillValue = 1.e+36f ;
		QRUNOFF:missing_value = 1.e+36f ;
	float QRUNOFF_NODYNLNDUSE(time, lndgrid) ;
		QRUNOFF_NODYNLNDUSE:long_name = "total liquid runoff (does not include QSNWCPICE) not including correction for land use change" ;
		QRUNOFF_NODYNLNDUSE:units = "mm/s" ;
		QRUNOFF_NODYNLNDUSE:cell_methods = "time: mean" ;
		QRUNOFF_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QRUNOFF_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QRUNOFF_R(time, lndgrid) ;
		QRUNOFF_R:long_name = "Rural total runoff" ;
		QRUNOFF_R:units = "mm/s" ;
		QRUNOFF_R:cell_methods = "time: mean" ;
		QRUNOFF_R:_FillValue = 1.e+36f ;
		QRUNOFF_R:missing_value = 1.e+36f ;
	float QRUNOFF_U(time, lndgrid) ;
		QRUNOFF_U:long_name = "Urban total runoff" ;
		QRUNOFF_U:units = "mm/s" ;
		QRUNOFF_U:cell_methods = "time: mean" ;
		QRUNOFF_U:_FillValue = 1.e+36f ;
		QRUNOFF_U:missing_value = 1.e+36f ;
	float QSNOMELT(time, lndgrid) ;
		QSNOMELT:long_name = "snow melt" ;
		QSNOMELT:units = "mm/s" ;
		QSNOMELT:cell_methods = "time: mean" ;
		QSNOMELT:_FillValue = 1.e+36f ;
		QSNOMELT:missing_value = 1.e+36f ;
	float QSNWCPICE(time, lndgrid) ;
		QSNWCPICE:long_name = "excess snowfall due to snow capping" ;
		QSNWCPICE:units = "mm/s" ;
		QSNWCPICE:cell_methods = "time: mean" ;
		QSNWCPICE:_FillValue = 1.e+36f ;
		QSNWCPICE:missing_value = 1.e+36f ;
	float QSNWCPICE_NODYNLNDUSE(time, lndgrid) ;
		QSNWCPICE_NODYNLNDUSE:long_name = "excess snowfall due to snow capping not including correction for land use change" ;
		QSNWCPICE_NODYNLNDUSE:units = "mm H2O/s" ;
		QSNWCPICE_NODYNLNDUSE:cell_methods = "time: mean" ;
		QSNWCPICE_NODYNLNDUSE:_FillValue = 1.e+36f ;
		QSNWCPICE_NODYNLNDUSE:missing_value = 1.e+36f ;
	float QSOIL(time, lndgrid) ;
		QSOIL:long_name = "Ground evaporation (soil/snow evaporation + soil/snow sublimation - dew)" ;
		QSOIL:units = "mm/s" ;
		QSOIL:cell_methods = "time: mean" ;
		QSOIL:_FillValue = 1.e+36f ;
		QSOIL:missing_value = 1.e+36f ;
	float QVEGE(time, lndgrid) ;
		QVEGE:long_name = "canopy evaporation" ;
		QVEGE:units = "mm/s" ;
		QVEGE:cell_methods = "time: mean" ;
		QVEGE:_FillValue = 1.e+36f ;
		QVEGE:missing_value = 1.e+36f ;
	float QVEGT(time, lndgrid) ;
		QVEGT:long_name = "canopy transpiration" ;
		QVEGT:units = "mm/s" ;
		QVEGT:cell_methods = "time: mean" ;
		QVEGT:_FillValue = 1.e+36f ;
		QVEGT:missing_value = 1.e+36f ;
	float RAIN(time, lndgrid) ;
		RAIN:long_name = "atmospheric rain" ;
		RAIN:units = "mm/s" ;
		RAIN:cell_methods = "time: mean" ;
		RAIN:_FillValue = 1.e+36f ;
		RAIN:missing_value = 1.e+36f ;
	float RETRANSN(time, lndgrid) ;
		RETRANSN:long_name = "plant pool of retranslocated N" ;
		RETRANSN:units = "gN/m^2" ;
		RETRANSN:cell_methods = "time: mean" ;
		RETRANSN:_FillValue = 1.e+36f ;
		RETRANSN:missing_value = 1.e+36f ;
	float RETRANSN_TO_NPOOL(time, lndgrid) ;
		RETRANSN_TO_NPOOL:long_name = "deployment of retranslocated N" ;
		RETRANSN_TO_NPOOL:units = "gN/m^2/s" ;
		RETRANSN_TO_NPOOL:cell_methods = "time: mean" ;
		RETRANSN_TO_NPOOL:_FillValue = 1.e+36f ;
		RETRANSN_TO_NPOOL:missing_value = 1.e+36f ;
	float RH2M(time, lndgrid) ;
		RH2M:long_name = "2m relative humidity" ;
		RH2M:units = "%" ;
		RH2M:cell_methods = "time: mean" ;
		RH2M:_FillValue = 1.e+36f ;
		RH2M:missing_value = 1.e+36f ;
	float RH2M_R(time, lndgrid) ;
		RH2M_R:long_name = "Rural 2m specific humidity" ;
		RH2M_R:units = "%" ;
		RH2M_R:cell_methods = "time: mean" ;
		RH2M_R:_FillValue = 1.e+36f ;
		RH2M_R:missing_value = 1.e+36f ;
	float RH2M_U(time, lndgrid) ;
		RH2M_U:long_name = "Urban 2m relative humidity" ;
		RH2M_U:units = "%" ;
		RH2M_U:cell_methods = "time: mean" ;
		RH2M_U:_FillValue = 1.e+36f ;
		RH2M_U:missing_value = 1.e+36f ;
	float RR(time, lndgrid) ;
		RR:long_name = "root respiration (fine root MR + total root GR)" ;
		RR:units = "gC/m^2/s" ;
		RR:cell_methods = "time: mean" ;
		RR:_FillValue = 1.e+36f ;
		RR:missing_value = 1.e+36f ;
	float SABG(time, lndgrid) ;
		SABG:long_name = "solar rad absorbed by ground" ;
		SABG:units = "W/m^2" ;
		SABG:cell_methods = "time: mean" ;
		SABG:_FillValue = 1.e+36f ;
		SABG:missing_value = 1.e+36f ;
	float SABG_PEN(time, lndgrid) ;
		SABG_PEN:long_name = "Rural solar rad penetrating top soil or snow layer" ;
		SABG_PEN:units = "watt/m^2" ;
		SABG_PEN:cell_methods = "time: mean" ;
		SABG_PEN:_FillValue = 1.e+36f ;
		SABG_PEN:missing_value = 1.e+36f ;
	float SABV(time, lndgrid) ;
		SABV:long_name = "solar rad absorbed by veg" ;
		SABV:units = "W/m^2" ;
		SABV:cell_methods = "time: mean" ;
		SABV:_FillValue = 1.e+36f ;
		SABV:missing_value = 1.e+36f ;
	float SEEDC(time, lndgrid) ;
		SEEDC:long_name = "pool for seeding new PFTs" ;
		SEEDC:units = "gC/m^2" ;
		SEEDC:cell_methods = "time: mean" ;
		SEEDC:_FillValue = 1.e+36f ;
		SEEDC:missing_value = 1.e+36f ;
	float SEEDN(time, lndgrid) ;
		SEEDN:long_name = "pool for seeding new PFTs" ;
		SEEDN:units = "gN/m^2" ;
		SEEDN:cell_methods = "time: mean" ;
		SEEDN:_FillValue = 1.e+36f ;
		SEEDN:missing_value = 1.e+36f ;
	float SMINN(time, lndgrid) ;
		SMINN:long_name = "soil mineral N" ;
		SMINN:units = "gN/m^2" ;
		SMINN:cell_methods = "time: mean" ;
		SMINN:_FillValue = 1.e+36f ;
		SMINN:missing_value = 1.e+36f ;
	float SMINN_TO_NPOOL(time, lndgrid) ;
		SMINN_TO_NPOOL:long_name = "deployment of soil mineral N uptake" ;
		SMINN_TO_NPOOL:units = "gN/m^2/s" ;
		SMINN_TO_NPOOL:cell_methods = "time: mean" ;
		SMINN_TO_NPOOL:_FillValue = 1.e+36f ;
		SMINN_TO_NPOOL:missing_value = 1.e+36f ;
	float SMINN_TO_PLANT(time, lndgrid) ;
		SMINN_TO_PLANT:long_name = "plant uptake of soil mineral N" ;
		SMINN_TO_PLANT:units = "gN/m^2/s" ;
		SMINN_TO_PLANT:cell_methods = "time: mean" ;
		SMINN_TO_PLANT:_FillValue = 1.e+36f ;
		SMINN_TO_PLANT:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L1(time, lndgrid) ;
		SMINN_TO_SOIL1N_L1:long_name = "mineral N flux for decomp. of LITR1to SOIL1" ;
		SMINN_TO_SOIL1N_L1:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_L2(time, lndgrid) ;
		SMINN_TO_SOIL1N_L2:long_name = "mineral N flux for decomp. of LITR2to SOIL1" ;
		SMINN_TO_SOIL1N_L2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_L2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_L2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_L2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S2(time, lndgrid) ;
		SMINN_TO_SOIL1N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL1" ;
		SMINN_TO_SOIL1N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S2:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL1N_S3(time, lndgrid) ;
		SMINN_TO_SOIL1N_S3:long_name = "mineral N flux for decomp. of SOIL3to SOIL1" ;
		SMINN_TO_SOIL1N_S3:units = "gN/m^2" ;
		SMINN_TO_SOIL1N_S3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL1N_S3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL1N_S3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_L3(time, lndgrid) ;
		SMINN_TO_SOIL2N_L3:long_name = "mineral N flux for decomp. of LITR3to SOIL2" ;
		SMINN_TO_SOIL2N_L3:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_L3:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_L3:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_L3:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL2N_S1(time, lndgrid) ;
		SMINN_TO_SOIL2N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL2" ;
		SMINN_TO_SOIL2N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL2N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL2N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL2N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S1(time, lndgrid) ;
		SMINN_TO_SOIL3N_S1:long_name = "mineral N flux for decomp. of SOIL1to SOIL3" ;
		SMINN_TO_SOIL3N_S1:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S1:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S1:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S1:missing_value = 1.e+36f ;
	float SMINN_TO_SOIL3N_S2(time, lndgrid) ;
		SMINN_TO_SOIL3N_S2:long_name = "mineral N flux for decomp. of SOIL2to SOIL3" ;
		SMINN_TO_SOIL3N_S2:units = "gN/m^2" ;
		SMINN_TO_SOIL3N_S2:cell_methods = "time: mean" ;
		SMINN_TO_SOIL3N_S2:_FillValue = 1.e+36f ;
		SMINN_TO_SOIL3N_S2:missing_value = 1.e+36f ;
	float SMIN_NH4(time, lndgrid) ;
		SMIN_NH4:long_name = "soil mineral NH4" ;
		SMIN_NH4:units = "gN/m^2" ;
		SMIN_NH4:cell_methods = "time: mean" ;
		SMIN_NH4:_FillValue = 1.e+36f ;
		SMIN_NH4:missing_value = 1.e+36f ;
	float SMIN_NH4_vr(time, levdcmp, lndgrid) ;
		SMIN_NH4_vr:long_name = "soil mineral NH4 (vert. res.)" ;
		SMIN_NH4_vr:units = "gN/m^3" ;
		SMIN_NH4_vr:cell_methods = "time: mean" ;
		SMIN_NH4_vr:_FillValue = 1.e+36f ;
		SMIN_NH4_vr:missing_value = 1.e+36f ;
	float SMIN_NO3(time, lndgrid) ;
		SMIN_NO3:long_name = "soil mineral NO3" ;
		SMIN_NO3:units = "gN/m^2" ;
		SMIN_NO3:cell_methods = "time: mean" ;
		SMIN_NO3:_FillValue = 1.e+36f ;
		SMIN_NO3:missing_value = 1.e+36f ;
	float SMIN_NO3_LEACHED(time, lndgrid) ;
		SMIN_NO3_LEACHED:long_name = "soil NO3 pool loss to leaching" ;
		SMIN_NO3_LEACHED:units = "gN/m^2/s" ;
		SMIN_NO3_LEACHED:cell_methods = "time: mean" ;
		SMIN_NO3_LEACHED:_FillValue = 1.e+36f ;
		SMIN_NO3_LEACHED:missing_value = 1.e+36f ;
	float SMIN_NO3_RUNOFF(time, lndgrid) ;
		SMIN_NO3_RUNOFF:long_name = "soil NO3 pool loss to runoff" ;
		SMIN_NO3_RUNOFF:units = "gN/m^2/s" ;
		SMIN_NO3_RUNOFF:cell_methods = "time: mean" ;
		SMIN_NO3_RUNOFF:_FillValue = 1.e+36f ;
		SMIN_NO3_RUNOFF:missing_value = 1.e+36f ;
	float SMIN_NO3_vr(time, levdcmp, lndgrid) ;
		SMIN_NO3_vr:long_name = "soil mineral NO3 (vert. res.)" ;
		SMIN_NO3_vr:units = "gN/m^3" ;
		SMIN_NO3_vr:cell_methods = "time: mean" ;
		SMIN_NO3_vr:_FillValue = 1.e+36f ;
		SMIN_NO3_vr:missing_value = 1.e+36f ;
	float SNOBCMCL(time, lndgrid) ;
		SNOBCMCL:long_name = "mass of BC in snow column" ;
		SNOBCMCL:units = "kg/m2" ;
		SNOBCMCL:cell_methods = "time: mean" ;
		SNOBCMCL:_FillValue = 1.e+36f ;
		SNOBCMCL:missing_value = 1.e+36f ;
	float SNOBCMSL(time, lndgrid) ;
		SNOBCMSL:long_name = "mass of BC in top snow layer" ;
		SNOBCMSL:units = "kg/m2" ;
		SNOBCMSL:cell_methods = "time: mean" ;
		SNOBCMSL:_FillValue = 1.e+36f ;
		SNOBCMSL:missing_value = 1.e+36f ;
	float SNODSTMCL(time, lndgrid) ;
		SNODSTMCL:long_name = "mass of dust in snow column" ;
		SNODSTMCL:units = "kg/m2" ;
		SNODSTMCL:cell_methods = "time: mean" ;
		SNODSTMCL:_FillValue = 1.e+36f ;
		SNODSTMCL:missing_value = 1.e+36f ;
	float SNODSTMSL(time, lndgrid) ;
		SNODSTMSL:long_name = "mass of dust in top snow layer" ;
		SNODSTMSL:units = "kg/m2" ;
		SNODSTMSL:cell_methods = "time: mean" ;
		SNODSTMSL:_FillValue = 1.e+36f ;
		SNODSTMSL:missing_value = 1.e+36f ;
	float SNOINTABS(time, lndgrid) ;
		SNOINTABS:long_name = "Percent of incoming solar absorbed by lower snow layers" ;
		SNOINTABS:units = "%" ;
		SNOINTABS:cell_methods = "time: mean" ;
		SNOINTABS:_FillValue = 1.e+36f ;
		SNOINTABS:missing_value = 1.e+36f ;
	float SNOOCMCL(time, lndgrid) ;
		SNOOCMCL:long_name = "mass of OC in snow column" ;
		SNOOCMCL:units = "kg/m2" ;
		SNOOCMCL:cell_methods = "time: mean" ;
		SNOOCMCL:_FillValue = 1.e+36f ;
		SNOOCMCL:missing_value = 1.e+36f ;
	float SNOOCMSL(time, lndgrid) ;
		SNOOCMSL:long_name = "mass of OC in top snow layer" ;
		SNOOCMSL:units = "kg/m2" ;
		SNOOCMSL:cell_methods = "time: mean" ;
		SNOOCMSL:_FillValue = 1.e+36f ;
		SNOOCMSL:missing_value = 1.e+36f ;
	float SNOW(time, lndgrid) ;
		SNOW:long_name = "atmospheric snow" ;
		SNOW:units = "mm/s" ;
		SNOW:cell_methods = "time: mean" ;
		SNOW:_FillValue = 1.e+36f ;
		SNOW:missing_value = 1.e+36f ;
	float SNOWDP(time, lndgrid) ;
		SNOWDP:long_name = "gridcell mean snow height" ;
		SNOWDP:units = "m" ;
		SNOWDP:cell_methods = "time: mean" ;
		SNOWDP:_FillValue = 1.e+36f ;
		SNOWDP:missing_value = 1.e+36f ;
	float SNOWICE(time, lndgrid) ;
		SNOWICE:long_name = "snow ice" ;
		SNOWICE:units = "kg/m2" ;
		SNOWICE:cell_methods = "time: mean" ;
		SNOWICE:_FillValue = 1.e+36f ;
		SNOWICE:missing_value = 1.e+36f ;
	float SNOWLIQ(time, lndgrid) ;
		SNOWLIQ:long_name = "snow liquid water" ;
		SNOWLIQ:units = "kg/m2" ;
		SNOWLIQ:cell_methods = "time: mean" ;
		SNOWLIQ:_FillValue = 1.e+36f ;
		SNOWLIQ:missing_value = 1.e+36f ;
	float SNOW_DEPTH(time, lndgrid) ;
		SNOW_DEPTH:long_name = "snow height of snow covered area" ;
		SNOW_DEPTH:units = "m" ;
		SNOW_DEPTH:cell_methods = "time: mean" ;
		SNOW_DEPTH:_FillValue = 1.e+36f ;
		SNOW_DEPTH:missing_value = 1.e+36f ;
	float SNOW_SINKS(time, lndgrid) ;
		SNOW_SINKS:long_name = "snow sinks (liquid water)" ;
		SNOW_SINKS:units = "mm/s" ;
		SNOW_SINKS:cell_methods = "time: mean" ;
		SNOW_SINKS:_FillValue = 1.e+36f ;
		SNOW_SINKS:missing_value = 1.e+36f ;
	float SNOW_SOURCES(time, lndgrid) ;
		SNOW_SOURCES:long_name = "snow sources (liquid water)" ;
		SNOW_SOURCES:units = "mm/s" ;
		SNOW_SOURCES:cell_methods = "time: mean" ;
		SNOW_SOURCES:_FillValue = 1.e+36f ;
		SNOW_SOURCES:missing_value = 1.e+36f ;
	float SOIL1C(time, lndgrid) ;
		SOIL1C:long_name = "SOIL1 C" ;
		SOIL1C:units = "gC/m^2" ;
		SOIL1C:cell_methods = "time: mean" ;
		SOIL1C:_FillValue = 1.e+36f ;
		SOIL1C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL2C(time, lndgrid) ;
		SOIL1C_TO_SOIL2C:long_name = "decomp. of soil 1 C to soil 2 C" ;
		SOIL1C_TO_SOIL2C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL2C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL2C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL2C:missing_value = 1.e+36f ;
	float SOIL1C_TO_SOIL3C(time, lndgrid) ;
		SOIL1C_TO_SOIL3C:long_name = "decomp. of soil 1 C to soil 3 C" ;
		SOIL1C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL1C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL1C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL1C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL1C_vr(time, levdcmp, lndgrid) ;
		SOIL1C_vr:long_name = "SOIL1 C (vertically resolved)" ;
		SOIL1C_vr:units = "gC/m^3" ;
		SOIL1C_vr:cell_methods = "time: mean" ;
		SOIL1C_vr:_FillValue = 1.e+36f ;
		SOIL1C_vr:missing_value = 1.e+36f ;
	float SOIL1N(time, lndgrid) ;
		SOIL1N:long_name = "SOIL1 N" ;
		SOIL1N:units = "gN/m^2" ;
		SOIL1N:cell_methods = "time: mean" ;
		SOIL1N:_FillValue = 1.e+36f ;
		SOIL1N:missing_value = 1.e+36f ;
	float SOIL1N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL1N_TNDNCY_VERT_TRANS:long_name = "soil 1 N tendency due to vertical transport" ;
		SOIL1N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL1N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL1N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL1N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL2N(time, lndgrid) ;
		SOIL1N_TO_SOIL2N:long_name = "decomp. of soil 1 N to soil 2 N" ;
		SOIL1N_TO_SOIL2N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL2N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL2N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL2N:missing_value = 1.e+36f ;
	float SOIL1N_TO_SOIL3N(time, lndgrid) ;
		SOIL1N_TO_SOIL3N:long_name = "decomp. of soil 1 N to soil 3 N" ;
		SOIL1N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL1N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL1N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL1N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL1N_vr(time, levdcmp, lndgrid) ;
		SOIL1N_vr:long_name = "SOIL1 N (vertically resolved)" ;
		SOIL1N_vr:units = "gN/m^3" ;
		SOIL1N_vr:cell_methods = "time: mean" ;
		SOIL1N_vr:_FillValue = 1.e+36f ;
		SOIL1N_vr:missing_value = 1.e+36f ;
	float SOIL1_HR_S2(time, lndgrid) ;
		SOIL1_HR_S2:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S2:units = "gC/m^2/s" ;
		SOIL1_HR_S2:cell_methods = "time: mean" ;
		SOIL1_HR_S2:_FillValue = 1.e+36f ;
		SOIL1_HR_S2:missing_value = 1.e+36f ;
	float SOIL1_HR_S3(time, lndgrid) ;
		SOIL1_HR_S3:long_name = "Het. Resp. from soil 1" ;
		SOIL1_HR_S3:units = "gC/m^2/s" ;
		SOIL1_HR_S3:cell_methods = "time: mean" ;
		SOIL1_HR_S3:_FillValue = 1.e+36f ;
		SOIL1_HR_S3:missing_value = 1.e+36f ;
	float SOIL2C(time, lndgrid) ;
		SOIL2C:long_name = "SOIL2 C" ;
		SOIL2C:units = "gC/m^2" ;
		SOIL2C:cell_methods = "time: mean" ;
		SOIL2C:_FillValue = 1.e+36f ;
		SOIL2C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL1C(time, lndgrid) ;
		SOIL2C_TO_SOIL1C:long_name = "decomp. of soil 2 C to soil 1 C" ;
		SOIL2C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL2C_TO_SOIL3C(time, lndgrid) ;
		SOIL2C_TO_SOIL3C:long_name = "decomp. of soil 2 C to soil 3 C" ;
		SOIL2C_TO_SOIL3C:units = "gC/m^2/s" ;
		SOIL2C_TO_SOIL3C:cell_methods = "time: mean" ;
		SOIL2C_TO_SOIL3C:_FillValue = 1.e+36f ;
		SOIL2C_TO_SOIL3C:missing_value = 1.e+36f ;
	float SOIL2C_vr(time, levdcmp, lndgrid) ;
		SOIL2C_vr:long_name = "SOIL2 C (vertically resolved)" ;
		SOIL2C_vr:units = "gC/m^3" ;
		SOIL2C_vr:cell_methods = "time: mean" ;
		SOIL2C_vr:_FillValue = 1.e+36f ;
		SOIL2C_vr:missing_value = 1.e+36f ;
	float SOIL2N(time, lndgrid) ;
		SOIL2N:long_name = "SOIL2 N" ;
		SOIL2N:units = "gN/m^2" ;
		SOIL2N:cell_methods = "time: mean" ;
		SOIL2N:_FillValue = 1.e+36f ;
		SOIL2N:missing_value = 1.e+36f ;
	float SOIL2N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL2N_TNDNCY_VERT_TRANS:long_name = "soil 2 N tendency due to vertical transport" ;
		SOIL2N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL2N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL2N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL2N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL1N(time, lndgrid) ;
		SOIL2N_TO_SOIL1N:long_name = "decomp. of soil 2 N to soil 1 N" ;
		SOIL2N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL2N_TO_SOIL3N(time, lndgrid) ;
		SOIL2N_TO_SOIL3N:long_name = "decomp. of soil 2 N to soil 3 N" ;
		SOIL2N_TO_SOIL3N:units = "gN/m^2" ;
		SOIL2N_TO_SOIL3N:cell_methods = "time: mean" ;
		SOIL2N_TO_SOIL3N:_FillValue = 1.e+36f ;
		SOIL2N_TO_SOIL3N:missing_value = 1.e+36f ;
	float SOIL2N_vr(time, levdcmp, lndgrid) ;
		SOIL2N_vr:long_name = "SOIL2 N (vertically resolved)" ;
		SOIL2N_vr:units = "gN/m^3" ;
		SOIL2N_vr:cell_methods = "time: mean" ;
		SOIL2N_vr:_FillValue = 1.e+36f ;
		SOIL2N_vr:missing_value = 1.e+36f ;
	float SOIL2_HR_S1(time, lndgrid) ;
		SOIL2_HR_S1:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S1:units = "gC/m^2/s" ;
		SOIL2_HR_S1:cell_methods = "time: mean" ;
		SOIL2_HR_S1:_FillValue = 1.e+36f ;
		SOIL2_HR_S1:missing_value = 1.e+36f ;
	float SOIL2_HR_S3(time, lndgrid) ;
		SOIL2_HR_S3:long_name = "Het. Resp. from soil 2" ;
		SOIL2_HR_S3:units = "gC/m^2/s" ;
		SOIL2_HR_S3:cell_methods = "time: mean" ;
		SOIL2_HR_S3:_FillValue = 1.e+36f ;
		SOIL2_HR_S3:missing_value = 1.e+36f ;
	float SOIL3C(time, lndgrid) ;
		SOIL3C:long_name = "SOIL3 C" ;
		SOIL3C:units = "gC/m^2" ;
		SOIL3C:cell_methods = "time: mean" ;
		SOIL3C:_FillValue = 1.e+36f ;
		SOIL3C:missing_value = 1.e+36f ;
	float SOIL3C_TO_SOIL1C(time, lndgrid) ;
		SOIL3C_TO_SOIL1C:long_name = "decomp. of soil 3 C to soil 1 C" ;
		SOIL3C_TO_SOIL1C:units = "gC/m^2/s" ;
		SOIL3C_TO_SOIL1C:cell_methods = "time: mean" ;
		SOIL3C_TO_SOIL1C:_FillValue = 1.e+36f ;
		SOIL3C_TO_SOIL1C:missing_value = 1.e+36f ;
	float SOIL3C_vr(time, levdcmp, lndgrid) ;
		SOIL3C_vr:long_name = "SOIL3 C (vertically resolved)" ;
		SOIL3C_vr:units = "gC/m^3" ;
		SOIL3C_vr:cell_methods = "time: mean" ;
		SOIL3C_vr:_FillValue = 1.e+36f ;
		SOIL3C_vr:missing_value = 1.e+36f ;
	float SOIL3N(time, lndgrid) ;
		SOIL3N:long_name = "SOIL3 N" ;
		SOIL3N:units = "gN/m^2" ;
		SOIL3N:cell_methods = "time: mean" ;
		SOIL3N:_FillValue = 1.e+36f ;
		SOIL3N:missing_value = 1.e+36f ;
	float SOIL3N_TNDNCY_VERT_TRANS(time, levdcmp, lndgrid) ;
		SOIL3N_TNDNCY_VERT_TRANS:long_name = "soil 3 N tendency due to vertical transport" ;
		SOIL3N_TNDNCY_VERT_TRANS:units = "gN/m^3/s" ;
		SOIL3N_TNDNCY_VERT_TRANS:cell_methods = "time: mean" ;
		SOIL3N_TNDNCY_VERT_TRANS:_FillValue = 1.e+36f ;
		SOIL3N_TNDNCY_VERT_TRANS:missing_value = 1.e+36f ;
	float SOIL3N_TO_SOIL1N(time, lndgrid) ;
		SOIL3N_TO_SOIL1N:long_name = "decomp. of soil 3 N to soil 1 N" ;
		SOIL3N_TO_SOIL1N:units = "gN/m^2" ;
		SOIL3N_TO_SOIL1N:cell_methods = "time: mean" ;
		SOIL3N_TO_SOIL1N:_FillValue = 1.e+36f ;
		SOIL3N_TO_SOIL1N:missing_value = 1.e+36f ;
	float SOIL3N_vr(time, levdcmp, lndgrid) ;
		SOIL3N_vr:long_name = "SOIL3 N (vertically resolved)" ;
		SOIL3N_vr:units = "gN/m^3" ;
		SOIL3N_vr:cell_methods = "time: mean" ;
		SOIL3N_vr:_FillValue = 1.e+36f ;
		SOIL3N_vr:missing_value = 1.e+36f ;
	float SOIL3_HR(time, lndgrid) ;
		SOIL3_HR:long_name = "Het. Resp. from soil 3" ;
		SOIL3_HR:units = "gC/m^2/s" ;
		SOIL3_HR:cell_methods = "time: mean" ;
		SOIL3_HR:_FillValue = 1.e+36f ;
		SOIL3_HR:missing_value = 1.e+36f ;
	float SOILC(time, lndgrid) ;
		SOILC:long_name = "soil C" ;
		SOILC:units = "gC/m^2" ;
		SOILC:cell_methods = "time: mean" ;
		SOILC:_FillValue = 1.e+36f ;
		SOILC:missing_value = 1.e+36f ;
	float SOILC_HR(time, lndgrid) ;
		SOILC_HR:long_name = "soil C heterotrophic respiration" ;
		SOILC_HR:units = "gC/m^2/s" ;
		SOILC_HR:cell_methods = "time: mean" ;
		SOILC_HR:_FillValue = 1.e+36f ;
		SOILC_HR:missing_value = 1.e+36f ;
	float SOILC_LOSS(time, lndgrid) ;
		SOILC_LOSS:long_name = "soil C loss" ;
		SOILC_LOSS:units = "gC/m^2/s" ;
		SOILC_LOSS:cell_methods = "time: mean" ;
		SOILC_LOSS:_FillValue = 1.e+36f ;
		SOILC_LOSS:missing_value = 1.e+36f ;
	float SOILICE(time, levgrnd, lndgrid) ;
		SOILICE:long_name = "soil ice (vegetated landunits only)" ;
		SOILICE:units = "kg/m2" ;
		SOILICE:cell_methods = "time: mean" ;
		SOILICE:_FillValue = 1.e+36f ;
		SOILICE:missing_value = 1.e+36f ;
	float SOILLIQ(time, levgrnd, lndgrid) ;
		SOILLIQ:long_name = "soil liquid water (vegetated landunits only)" ;
		SOILLIQ:units = "kg/m2" ;
		SOILLIQ:cell_methods = "time: mean" ;
		SOILLIQ:_FillValue = 1.e+36f ;
		SOILLIQ:missing_value = 1.e+36f ;
	float SOILPSI(time, levgrnd, lndgrid) ;
		SOILPSI:long_name = "soil water potential in each soil layer" ;
		SOILPSI:units = "MPa" ;
		SOILPSI:cell_methods = "time: mean" ;
		SOILPSI:_FillValue = 1.e+36f ;
		SOILPSI:missing_value = 1.e+36f ;
	float SOILWATER_10CM(time, lndgrid) ;
		SOILWATER_10CM:long_name = "soil liquid water + ice in top 10cm of soil (veg landunits only)" ;
		SOILWATER_10CM:units = "kg/m2" ;
		SOILWATER_10CM:cell_methods = "time: mean" ;
		SOILWATER_10CM:_FillValue = 1.e+36f ;
		SOILWATER_10CM:missing_value = 1.e+36f ;
	float SOMC_FIRE(time, lndgrid) ;
		SOMC_FIRE:long_name = "C loss due to peat burning" ;
		SOMC_FIRE:units = "gC/m^2/s" ;
		SOMC_FIRE:cell_methods = "time: mean" ;
		SOMC_FIRE:_FillValue = 1.e+36f ;
		SOMC_FIRE:missing_value = 1.e+36f ;
	float SOMHR(time, lndgrid) ;
		SOMHR:long_name = "soil organic matter heterotrophic respiration" ;
		SOMHR:units = "gC/m^2/s" ;
		SOMHR:cell_methods = "time: mean" ;
		SOMHR:_FillValue = 1.e+36f ;
		SOMHR:missing_value = 1.e+36f ;
	float SOM_C_LEACHED(time, lndgrid) ;
		SOM_C_LEACHED:long_name = "total flux of C from SOM pools due to leaching" ;
		SOM_C_LEACHED:units = "gC/m^2/s" ;
		SOM_C_LEACHED:cell_methods = "time: mean" ;
		SOM_C_LEACHED:_FillValue = 1.e+36f ;
		SOM_C_LEACHED:missing_value = 1.e+36f ;
	float SR(time, lndgrid) ;
		SR:long_name = "total soil respiration (HR + root resp)" ;
		SR:units = "gC/m^2/s" ;
		SR:cell_methods = "time: mean" ;
		SR:_FillValue = 1.e+36f ;
		SR:missing_value = 1.e+36f ;
	float STORVEGC(time, lndgrid) ;
		STORVEGC:long_name = "stored vegetation carbon, excluding cpool" ;
		STORVEGC:units = "gC/m^2" ;
		STORVEGC:cell_methods = "time: mean" ;
		STORVEGC:_FillValue = 1.e+36f ;
		STORVEGC:missing_value = 1.e+36f ;
	float STORVEGN(time, lndgrid) ;
		STORVEGN:long_name = "stored vegetation nitrogen" ;
		STORVEGN:units = "gN/m^2" ;
		STORVEGN:cell_methods = "time: mean" ;
		STORVEGN:_FillValue = 1.e+36f ;
		STORVEGN:missing_value = 1.e+36f ;
	float SUPPLEMENT_TO_SMINN(time, lndgrid) ;
		SUPPLEMENT_TO_SMINN:long_name = "supplemental N supply" ;
		SUPPLEMENT_TO_SMINN:units = "gN/m^2/s" ;
		SUPPLEMENT_TO_SMINN:cell_methods = "time: mean" ;
		SUPPLEMENT_TO_SMINN:_FillValue = 1.e+36f ;
		SUPPLEMENT_TO_SMINN:missing_value = 1.e+36f ;
	float SoilAlpha(time, lndgrid) ;
		SoilAlpha:long_name = "factor limiting ground evap" ;
		SoilAlpha:units = "unitless" ;
		SoilAlpha:cell_methods = "time: mean" ;
		SoilAlpha:_FillValue = 1.e+36f ;
		SoilAlpha:missing_value = 1.e+36f ;
	float SoilAlpha_U(time, lndgrid) ;
		SoilAlpha_U:long_name = "urban factor limiting ground evap" ;
		SoilAlpha_U:units = "unitless" ;
		SoilAlpha_U:cell_methods = "time: mean" ;
		SoilAlpha_U:_FillValue = 1.e+36f ;
		SoilAlpha_U:missing_value = 1.e+36f ;
	float TAUX(time, lndgrid) ;
		TAUX:long_name = "zonal surface stress" ;
		TAUX:units = "kg/m/s^2" ;
		TAUX:cell_methods = "time: mean" ;
		TAUX:_FillValue = 1.e+36f ;
		TAUX:missing_value = 1.e+36f ;
	float TAUY(time, lndgrid) ;
		TAUY:long_name = "meridional surface stress" ;
		TAUY:units = "kg/m/s^2" ;
		TAUY:cell_methods = "time: mean" ;
		TAUY:_FillValue = 1.e+36f ;
		TAUY:missing_value = 1.e+36f ;
	float TBOT(time, lndgrid) ;
		TBOT:long_name = "atmospheric air temperature" ;
		TBOT:units = "K" ;
		TBOT:cell_methods = "time: mean" ;
		TBOT:_FillValue = 1.e+36f ;
		TBOT:missing_value = 1.e+36f ;
	float TBUILD(time, lndgrid) ;
		TBUILD:long_name = "internal urban building temperature" ;
		TBUILD:units = "K" ;
		TBUILD:cell_methods = "time: mean" ;
		TBUILD:_FillValue = 1.e+36f ;
		TBUILD:missing_value = 1.e+36f ;
	float TG(time, lndgrid) ;
		TG:long_name = "ground temperature" ;
		TG:units = "K" ;
		TG:cell_methods = "time: mean" ;
		TG:_FillValue = 1.e+36f ;
		TG:missing_value = 1.e+36f ;
	float TG_R(time, lndgrid) ;
		TG_R:long_name = "Rural ground temperature" ;
		TG_R:units = "K" ;
		TG_R:cell_methods = "time: mean" ;
		TG_R:_FillValue = 1.e+36f ;
		TG_R:missing_value = 1.e+36f ;
	float TG_U(time, lndgrid) ;
		TG_U:long_name = "Urban ground temperature" ;
		TG_U:units = "K" ;
		TG_U:cell_methods = "time: mean" ;
		TG_U:_FillValue = 1.e+36f ;
		TG_U:missing_value = 1.e+36f ;
	float TH2OSFC(time, lndgrid) ;
		TH2OSFC:long_name = "surface water temperature" ;
		TH2OSFC:units = "K" ;
		TH2OSFC:cell_methods = "time: mean" ;
		TH2OSFC:_FillValue = 1.e+36f ;
		TH2OSFC:missing_value = 1.e+36f ;
	float THBOT(time, lndgrid) ;
		THBOT:long_name = "atmospheric air potential temperature" ;
		THBOT:units = "K" ;
		THBOT:cell_methods = "time: mean" ;
		THBOT:_FillValue = 1.e+36f ;
		THBOT:missing_value = 1.e+36f ;
	float TKE1(time, lndgrid) ;
		TKE1:long_name = "top lake level eddy thermal conductivity" ;
		TKE1:units = "W/(mK)" ;
		TKE1:cell_methods = "time: mean" ;
		TKE1:_FillValue = 1.e+36f ;
		TKE1:missing_value = 1.e+36f ;
	float TLAI(time, lndgrid) ;
		TLAI:long_name = "total projected leaf area index" ;
		TLAI:units = "none" ;
		TLAI:cell_methods = "time: mean" ;
		TLAI:_FillValue = 1.e+36f ;
		TLAI:missing_value = 1.e+36f ;
	float TLAKE(time, levlak, lndgrid) ;
		TLAKE:long_name = "lake temperature" ;
		TLAKE:units = "K" ;
		TLAKE:cell_methods = "time: mean" ;
		TLAKE:_FillValue = 1.e+36f ;
		TLAKE:missing_value = 1.e+36f ;
	float TOTCOLC(time, lndgrid) ;
		TOTCOLC:long_name = "total column carbon, incl veg and cpool" ;
		TOTCOLC:units = "gC/m^2" ;
		TOTCOLC:cell_methods = "time: mean" ;
		TOTCOLC:_FillValue = 1.e+36f ;
		TOTCOLC:missing_value = 1.e+36f ;
	float TOTCOLCH4(time, lndgrid) ;
		TOTCOLCH4:long_name = "total belowground CH4, (0 for non-lake special landunits)" ;
		TOTCOLCH4:units = "gC/m2" ;
		TOTCOLCH4:cell_methods = "time: mean" ;
		TOTCOLCH4:_FillValue = 1.e+36f ;
		TOTCOLCH4:missing_value = 1.e+36f ;
	float TOTCOLN(time, lndgrid) ;
		TOTCOLN:long_name = "total column-level N" ;
		TOTCOLN:units = "gN/m^2" ;
		TOTCOLN:cell_methods = "time: mean" ;
		TOTCOLN:_FillValue = 1.e+36f ;
		TOTCOLN:missing_value = 1.e+36f ;
	float TOTECOSYSC(time, lndgrid) ;
		TOTECOSYSC:long_name = "total ecosystem carbon, incl veg but excl cpool" ;
		TOTECOSYSC:units = "gC/m^2" ;
		TOTECOSYSC:cell_methods = "time: mean" ;
		TOTECOSYSC:_FillValue = 1.e+36f ;
		TOTECOSYSC:missing_value = 1.e+36f ;
	float TOTECOSYSN(time, lndgrid) ;
		TOTECOSYSN:long_name = "total ecosystem N" ;
		TOTECOSYSN:units = "gN/m^2" ;
		TOTECOSYSN:cell_methods = "time: mean" ;
		TOTECOSYSN:_FillValue = 1.e+36f ;
		TOTECOSYSN:missing_value = 1.e+36f ;
	float TOTLITC(time, lndgrid) ;
		TOTLITC:long_name = "total litter carbon" ;
		TOTLITC:units = "gC/m^2" ;
		TOTLITC:cell_methods = "time: mean" ;
		TOTLITC:_FillValue = 1.e+36f ;
		TOTLITC:missing_value = 1.e+36f ;
	float TOTLITC_1m(time, lndgrid) ;
		TOTLITC_1m:long_name = "total litter carbon to 1 meter depth" ;
		TOTLITC_1m:units = "gC/m^2" ;
		TOTLITC_1m:cell_methods = "time: mean" ;
		TOTLITC_1m:_FillValue = 1.e+36f ;
		TOTLITC_1m:missing_value = 1.e+36f ;
	float TOTLITN(time, lndgrid) ;
		TOTLITN:long_name = "total litter N" ;
		TOTLITN:units = "gN/m^2" ;
		TOTLITN:cell_methods = "time: mean" ;
		TOTLITN:_FillValue = 1.e+36f ;
		TOTLITN:missing_value = 1.e+36f ;
	float TOTLITN_1m(time, lndgrid) ;
		TOTLITN_1m:long_name = "total litter N to 1 meter" ;
		TOTLITN_1m:units = "gN/m^2" ;
		TOTLITN_1m:cell_methods = "time: mean" ;
		TOTLITN_1m:_FillValue = 1.e+36f ;
		TOTLITN_1m:missing_value = 1.e+36f ;
	float TOTPFTC(time, lndgrid) ;
		TOTPFTC:long_name = "total pft-level carbon, including cpool" ;
		TOTPFTC:units = "gC/m^2" ;
		TOTPFTC:cell_methods = "time: mean" ;
		TOTPFTC:_FillValue = 1.e+36f ;
		TOTPFTC:missing_value = 1.e+36f ;
	float TOTPFTN(time, lndgrid) ;
		TOTPFTN:long_name = "total PFT-level nitrogen" ;
		TOTPFTN:units = "gN/m^2" ;
		TOTPFTN:cell_methods = "time: mean" ;
		TOTPFTN:_FillValue = 1.e+36f ;
		TOTPFTN:missing_value = 1.e+36f ;
	float TOTPRODC(time, lndgrid) ;
		TOTPRODC:long_name = "total wood product C" ;
		TOTPRODC:units = "gC/m^2" ;
		TOTPRODC:cell_methods = "time: mean" ;
		TOTPRODC:_FillValue = 1.e+36f ;
		TOTPRODC:missing_value = 1.e+36f ;
	float TOTPRODN(time, lndgrid) ;
		TOTPRODN:long_name = "total wood product N" ;
		TOTPRODN:units = "gN/m^2" ;
		TOTPRODN:cell_methods = "time: mean" ;
		TOTPRODN:_FillValue = 1.e+36f ;
		TOTPRODN:missing_value = 1.e+36f ;
	float TOTSOMC(time, lndgrid) ;
		TOTSOMC:long_name = "total soil organic matter carbon" ;
		TOTSOMC:units = "gC/m^2" ;
		TOTSOMC:cell_methods = "time: mean" ;
		TOTSOMC:_FillValue = 1.e+36f ;
		TOTSOMC:missing_value = 1.e+36f ;
	float TOTSOMC_1m(time, lndgrid) ;
		TOTSOMC_1m:long_name = "total soil organic matter carbon to 1 meter depth" ;
		TOTSOMC_1m:units = "gC/m^2" ;
		TOTSOMC_1m:cell_methods = "time: mean" ;
		TOTSOMC_1m:_FillValue = 1.e+36f ;
		TOTSOMC_1m:missing_value = 1.e+36f ;
	float TOTSOMN(time, lndgrid) ;
		TOTSOMN:long_name = "total soil organic matter N" ;
		TOTSOMN:units = "gN/m^2" ;
		TOTSOMN:cell_methods = "time: mean" ;
		TOTSOMN:_FillValue = 1.e+36f ;
		TOTSOMN:missing_value = 1.e+36f ;
	float TOTSOMN_1m(time, lndgrid) ;
		TOTSOMN_1m:long_name = "total soil organic matter N to 1 meter" ;
		TOTSOMN_1m:units = "gN/m^2" ;
		TOTSOMN_1m:cell_methods = "time: mean" ;
		TOTSOMN_1m:_FillValue = 1.e+36f ;
		TOTSOMN_1m:missing_value = 1.e+36f ;
	float TOTVEGC(time, lndgrid) ;
		TOTVEGC:long_name = "total vegetation carbon, excluding cpool" ;
		TOTVEGC:units = "gC/m^2" ;
		TOTVEGC:cell_methods = "time: mean" ;
		TOTVEGC:_FillValue = 1.e+36f ;
		TOTVEGC:missing_value = 1.e+36f ;
	float TOTVEGN(time, lndgrid) ;
		TOTVEGN:long_name = "total vegetation nitrogen" ;
		TOTVEGN:units = "gN/m^2" ;
		TOTVEGN:cell_methods = "time: mean" ;
		TOTVEGN:_FillValue = 1.e+36f ;
		TOTVEGN:missing_value = 1.e+36f ;
	float TREFMNAV(time, lndgrid) ;
		TREFMNAV:long_name = "daily minimum of average 2-m temperature" ;
		TREFMNAV:units = "K" ;
		TREFMNAV:cell_methods = "time: mean" ;
		TREFMNAV:_FillValue = 1.e+36f ;
		TREFMNAV:missing_value = 1.e+36f ;
	float TREFMNAV_R(time, lndgrid) ;
		TREFMNAV_R:long_name = "Rural daily minimum of average 2-m temperature" ;
		TREFMNAV_R:units = "K" ;
		TREFMNAV_R:cell_methods = "time: mean" ;
		TREFMNAV_R:_FillValue = 1.e+36f ;
		TREFMNAV_R:missing_value = 1.e+36f ;
	float TREFMNAV_U(time, lndgrid) ;
		TREFMNAV_U:long_name = "Urban daily minimum of average 2-m temperature" ;
		TREFMNAV_U:units = "K" ;
		TREFMNAV_U:cell_methods = "time: mean" ;
		TREFMNAV_U:_FillValue = 1.e+36f ;
		TREFMNAV_U:missing_value = 1.e+36f ;
	float TREFMXAV(time, lndgrid) ;
		TREFMXAV:long_name = "daily maximum of average 2-m temperature" ;
		TREFMXAV:units = "K" ;
		TREFMXAV:cell_methods = "time: mean" ;
		TREFMXAV:_FillValue = 1.e+36f ;
		TREFMXAV:missing_value = 1.e+36f ;
	float TREFMXAV_R(time, lndgrid) ;
		TREFMXAV_R:long_name = "Rural daily maximum of average 2-m temperature" ;
		TREFMXAV_R:units = "K" ;
		TREFMXAV_R:cell_methods = "time: mean" ;
		TREFMXAV_R:_FillValue = 1.e+36f ;
		TREFMXAV_R:missing_value = 1.e+36f ;
	float TREFMXAV_U(time, lndgrid) ;
		TREFMXAV_U:long_name = "Urban daily maximum of average 2-m temperature" ;
		TREFMXAV_U:units = "K" ;
		TREFMXAV_U:cell_methods = "time: mean" ;
		TREFMXAV_U:_FillValue = 1.e+36f ;
		TREFMXAV_U:missing_value = 1.e+36f ;
	float TSA(time, lndgrid) ;
		TSA:long_name = "2m air temperature" ;
		TSA:units = "K" ;
		TSA:cell_methods = "time: mean" ;
		TSA:_FillValue = 1.e+36f ;
		TSA:missing_value = 1.e+36f ;
	float TSAI(time, lndgrid) ;
		TSAI:long_name = "total projected stem area index" ;
		TSAI:units = "none" ;
		TSAI:cell_methods = "time: mean" ;
		TSAI:_FillValue = 1.e+36f ;
		TSAI:missing_value = 1.e+36f ;
	float TSA_R(time, lndgrid) ;
		TSA_R:long_name = "Rural 2m air temperature" ;
		TSA_R:units = "K" ;
		TSA_R:cell_methods = "time: mean" ;
		TSA_R:_FillValue = 1.e+36f ;
		TSA_R:missing_value = 1.e+36f ;
	float TSA_U(time, lndgrid) ;
		TSA_U:long_name = "Urban 2m air temperature" ;
		TSA_U:units = "K" ;
		TSA_U:cell_methods = "time: mean" ;
		TSA_U:_FillValue = 1.e+36f ;
		TSA_U:missing_value = 1.e+36f ;
	float TSOI(time, levgrnd, lndgrid) ;
		TSOI:long_name = "soil temperature (vegetated landunits only)" ;
		TSOI:units = "K" ;
		TSOI:cell_methods = "time: mean" ;
		TSOI:_FillValue = 1.e+36f ;
		TSOI:missing_value = 1.e+36f ;
	float TSOI_10CM(time, lndgrid) ;
		TSOI_10CM:long_name = "soil temperature in top 10cm of soil" ;
		TSOI_10CM:units = "K" ;
		TSOI_10CM:cell_methods = "time: mean" ;
		TSOI_10CM:_FillValue = 1.e+36f ;
		TSOI_10CM:missing_value = 1.e+36f ;
	float TSOI_ICE(time, levgrnd, lndgrid) ;
		TSOI_ICE:long_name = "soil temperature (ice landunits only)" ;
		TSOI_ICE:units = "K" ;
		TSOI_ICE:cell_methods = "time: mean" ;
		TSOI_ICE:_FillValue = 1.e+36f ;
		TSOI_ICE:missing_value = 1.e+36f ;
	float TV(time, lndgrid) ;
		TV:long_name = "vegetation temperature" ;
		TV:units = "K" ;
		TV:cell_methods = "time: mean" ;
		TV:_FillValue = 1.e+36f ;
		TV:missing_value = 1.e+36f ;
	float TWS(time, lndgrid) ;
		TWS:long_name = "total water storage" ;
		TWS:units = "mm" ;
		TWS:cell_methods = "time: mean" ;
		TWS:_FillValue = 1.e+36f ;
		TWS:missing_value = 1.e+36f ;
	float T_SCALAR(time, levdcmp, lndgrid) ;
		T_SCALAR:long_name = "temperature inhibition of decomposition" ;
		T_SCALAR:units = "unitless" ;
		T_SCALAR:cell_methods = "time: mean" ;
		T_SCALAR:_FillValue = 1.e+36f ;
		T_SCALAR:missing_value = 1.e+36f ;
	float U10(time, lndgrid) ;
		U10:long_name = "10-m wind" ;
		U10:units = "m/s" ;
		U10:cell_methods = "time: mean" ;
		U10:_FillValue = 1.e+36f ;
		U10:missing_value = 1.e+36f ;
	float URBAN_AC(time, lndgrid) ;
		URBAN_AC:long_name = "urban air conditioning flux" ;
		URBAN_AC:units = "W/m^2" ;
		URBAN_AC:cell_methods = "time: mean" ;
		URBAN_AC:_FillValue = 1.e+36f ;
		URBAN_AC:missing_value = 1.e+36f ;
	float URBAN_HEAT(time, lndgrid) ;
		URBAN_HEAT:long_name = "urban heating flux" ;
		URBAN_HEAT:units = "W/m^2" ;
		URBAN_HEAT:cell_methods = "time: mean" ;
		URBAN_HEAT:_FillValue = 1.e+36f ;
		URBAN_HEAT:missing_value = 1.e+36f ;
	float VOCFLXT(time, lndgrid) ;
		VOCFLXT:long_name = "total VOC flux into atmosphere" ;
		VOCFLXT:units = "moles/m2/sec" ;
		VOCFLXT:cell_methods = "time: mean" ;
		VOCFLXT:_FillValue = 1.e+36f ;
		VOCFLXT:missing_value = 1.e+36f ;
	float VOLR(time, lndgrid) ;
		VOLR:long_name = "river channel water storage" ;
		VOLR:units = "m3" ;
		VOLR:cell_methods = "time: mean" ;
		VOLR:_FillValue = 1.e+36f ;
		VOLR:missing_value = 1.e+36f ;
	float WA(time, lndgrid) ;
		WA:long_name = "water in the unconfined aquifer (vegetated landunits only)" ;
		WA:units = "mm" ;
		WA:cell_methods = "time: mean" ;
		WA:_FillValue = 1.e+36f ;
		WA:missing_value = 1.e+36f ;
	float WASTEHEAT(time, lndgrid) ;
		WASTEHEAT:long_name = "sensible heat flux from heating/cooling sources of urban waste heat" ;
		WASTEHEAT:units = "W/m^2" ;
		WASTEHEAT:cell_methods = "time: mean" ;
		WASTEHEAT:_FillValue = 1.e+36f ;
		WASTEHEAT:missing_value = 1.e+36f ;
	float WF(time, lndgrid) ;
		WF:long_name = "soil water as frac. of whc for top 0.05 m" ;
		WF:units = "proportion" ;
		WF:cell_methods = "time: mean" ;
		WF:_FillValue = 1.e+36f ;
		WF:missing_value = 1.e+36f ;
	float WIND(time, lndgrid) ;
		WIND:long_name = "atmospheric wind velocity magnitude" ;
		WIND:units = "m/s" ;
		WIND:cell_methods = "time: mean" ;
		WIND:_FillValue = 1.e+36f ;
		WIND:missing_value = 1.e+36f ;
	float WOODC(time, lndgrid) ;
		WOODC:long_name = "wood C" ;
		WOODC:units = "gC/m^2" ;
		WOODC:cell_methods = "time: mean" ;
		WOODC:_FillValue = 1.e+36f ;
		WOODC:missing_value = 1.e+36f ;
	float WOODC_ALLOC(time, lndgrid) ;
		WOODC_ALLOC:long_name = "wood C allocation" ;
		WOODC_ALLOC:units = "gC/m^2/s" ;
		WOODC_ALLOC:cell_methods = "time: mean" ;
		WOODC_ALLOC:_FillValue = 1.e+36f ;
		WOODC_ALLOC:missing_value = 1.e+36f ;
	float WOODC_LOSS(time, lndgrid) ;
		WOODC_LOSS:long_name = "wood C loss" ;
		WOODC_LOSS:units = "gC/m^2/s" ;
		WOODC_LOSS:cell_methods = "time: mean" ;
		WOODC_LOSS:_FillValue = 1.e+36f ;
		WOODC_LOSS:missing_value = 1.e+36f ;
	float WOOD_HARVESTC(time, lndgrid) ;
		WOOD_HARVESTC:long_name = "wood harvest carbon (to product pools)" ;
		WOOD_HARVESTC:units = "gC/m^2/s" ;
		WOOD_HARVESTC:cell_methods = "time: mean" ;
		WOOD_HARVESTC:_FillValue = 1.e+36f ;
		WOOD_HARVESTC:missing_value = 1.e+36f ;
	float WOOD_HARVESTN(time, lndgrid) ;
		WOOD_HARVESTN:long_name = "wood harvest N (to product pools)" ;
		WOOD_HARVESTN:units = "gN/m^2/s" ;
		WOOD_HARVESTN:cell_methods = "time: mean" ;
		WOOD_HARVESTN:_FillValue = 1.e+36f ;
		WOOD_HARVESTN:missing_value = 1.e+36f ;
	float WTGQ(time, lndgrid) ;
		WTGQ:long_name = "surface tracer conductance" ;
		WTGQ:units = "m/s" ;
		WTGQ:cell_methods = "time: mean" ;
		WTGQ:_FillValue = 1.e+36f ;
		WTGQ:missing_value = 1.e+36f ;
	float W_SCALAR(time, levdcmp, lndgrid) ;
		W_SCALAR:long_name = "Moisture (dryness) inhibition of decomposition" ;
		W_SCALAR:units = "unitless" ;
		W_SCALAR:cell_methods = "time: mean" ;
		W_SCALAR:_FillValue = 1.e+36f ;
		W_SCALAR:missing_value = 1.e+36f ;
	float XSMRPOOL(time, lndgrid) ;
		XSMRPOOL:long_name = "temporary photosynthate C pool" ;
		XSMRPOOL:units = "gC/m^2" ;
		XSMRPOOL:cell_methods = "time: mean" ;
		XSMRPOOL:_FillValue = 1.e+36f ;
		XSMRPOOL:missing_value = 1.e+36f ;
	float XSMRPOOL_RECOVER(time, lndgrid) ;
		XSMRPOOL_RECOVER:long_name = "C flux assigned to recovery of negative xsmrpool" ;
		XSMRPOOL_RECOVER:units = "gC/m^2/s" ;
		XSMRPOOL_RECOVER:cell_methods = "time: mean" ;
		XSMRPOOL_RECOVER:_FillValue = 1.e+36f ;
		XSMRPOOL_RECOVER:missing_value = 1.e+36f ;
	float ZBOT(time, lndgrid) ;
		ZBOT:long_name = "atmospheric reference height" ;
		ZBOT:units = "m" ;
		ZBOT:cell_methods = "time: mean" ;
		ZBOT:_FillValue = 1.e+36f ;
		ZBOT:missing_value = 1.e+36f ;
	float ZWT(time, lndgrid) ;
		ZWT:long_name = "water table depth (vegetated landunits only)" ;
		ZWT:units = "m" ;
		ZWT:cell_methods = "time: mean" ;
		ZWT:_FillValue = 1.e+36f ;
		ZWT:missing_value = 1.e+36f ;
	float ZWT_CH4_UNSAT(time, lndgrid) ;
		ZWT_CH4_UNSAT:long_name = "depth of water table for methane production used in non-inundated area" ;
		ZWT_CH4_UNSAT:units = "m" ;
		ZWT_CH4_UNSAT:cell_methods = "time: mean" ;
		ZWT_CH4_UNSAT:_FillValue = 1.e+36f ;
		ZWT_CH4_UNSAT:missing_value = 1.e+36f ;
	float ZWT_PERCH(time, lndgrid) ;
		ZWT_PERCH:long_name = "perched water table depth (vegetated landunits only)" ;
		ZWT_PERCH:units = "m" ;
		ZWT_PERCH:cell_methods = "time: mean" ;
		ZWT_PERCH:_FillValue = 1.e+36f ;
		ZWT_PERCH:missing_value = 1.e+36f ;
	float o2_decomp_depth_unsat(time, levgrnd, lndgrid) ;
		o2_decomp_depth_unsat:long_name = "o2_decomp_depth_unsat" ;
		o2_decomp_depth_unsat:units = "mol/m3/2" ;
		o2_decomp_depth_unsat:cell_methods = "time: mean" ;
		o2_decomp_depth_unsat:_FillValue = 1.e+36f ;
		o2_decomp_depth_unsat:missing_value = 1.e+36f ;

// global attributes:
		:title = "CLM History file information" ;
		:comment = "NOTE: None of the variables are weighted by land fraction!" ;
		:Conventions = "CF-1.0" ;
		:history = "created on 09/25/14 13:24:56" ;
		:source = "Community Land Model CLM4.0" ;
		:hostname = "userdefined" ;
		:username = "gbisht" ;
		:version = "" ;
		:revision_id = "$Id: histFileMod.F90 42903 2012-12-21 15:32:10Z muszala $" ;
		:case_title = "UNSET" ;
		:case_id = "ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-4" ;
		:Surface_dataset = "surfdata_13x26pt_US-Brw_simyr1850.nc" ;
		:Initial_conditions_dataset = "arbitrary initialization" ;
		:PFT_physiological_constants_dataset = "clm_params.c140423.nc" ;
		:ltype_vegetated_or_bare_soil = 1 ;
		:ltype_crop = 2 ;
		:ltype_landice = 3 ;
		:ltype_landice_multiple_elevation_classes = 4 ;
		:ltype_deep_lake = 5 ;
		:ltype_wetland = 6 ;
		:ltype_urban_tbd = 7 ;
		:ltype_urban_hd = 8 ;
		:ltype_urban_md = 9 ;
		:natpft_not_vegetated = 1 ;
		:natpft_needleleaf_evergreen_temperate_tree = 2 ;
		:natpft_needleleaf_evergreen_boreal_tree = 3 ;
		:natpft_needleleaf_deciduous_boreal_tree = 4 ;
		:natpft_broadleaf_evergreen_tropical_tree = 5 ;
		:natpft_broadleaf_evergreen_temperate_tree = 6 ;
		:natpft_broadleaf_deciduous_tropical_tree = 7 ;
		:natpft_broadleaf_deciduous_temperate_tree = 8 ;
		:natpft_broadleaf_deciduous_boreal_tree = 9 ;
		:natpft_broadleaf_evergreen_shrub = 10 ;
		:natpft_broadleaf_deciduous_temperate_shrub = 11 ;
		:natpft_broadleaf_deciduous_boreal_shrub = 12 ;
		:natpft_c3_arctic_grass = 13 ;
		:natpft_c3_non-arctic_grass = 14 ;
		:natpft_c4_grass = 15 ;
		:natpft_c3_crop = 16 ;
		:natpft_c3_irrigated = 17 ;
		:Time_constant_3Dvars_filename = "./ugrid-13x26x10-subsurface-th-noice-dec-NGEE_SiteB-np-4.clm2.h0.0001-12-01-00000.nc" ;
		:Time_constant_3Dvars = "ZSOI:DZSOI:WATSAT:SUCSAT:BSW:HKSAT:ZLAKE:DZLAKE" ;
data:

 levgrnd = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 levlak = 0.05, 0.6, 2.1, 4.6, 8.1, 12.6, 18.6, 25.6, 34.325, 44.775 ;

 levdcmp = 0.007100635, 0.027925, 0.06225858, 0.1188651, 0.2121934, 
    0.3660658, 0.6197585, 1.038027, 1.727635, 2.864607, 4.739157, 7.829766, 
    12.92532, 21.32647, 35.17762 ;

 time = 1 ;

 mcdate = 11202 ;

 mcsec = 0 ;

 mdcur = 1 ;

 mscur = 0 ;

 nstep = 48 ;

 time_bounds =
  0, 1 ;

 date_written =
  "09/25/14" ;

 time_written =
  "13:24:56" ;

 lon = -156.6089, -156.6089, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6083, -156.6082, -156.608, -156.608, -156.6078, -156.6078, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, 
    -156.6069, -156.6069, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6063, -156.6062, -156.6089, -156.6089, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6083, -156.6082, -156.608, -156.608, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6074, -156.6073, 
    -156.6071, -156.6071, -156.6069, -156.6069, -156.6067, -156.6066, 
    -156.6065, -156.6064, -156.6063, -156.6062, -156.6089, -156.6089, 
    -156.6087, -156.6086, -156.6085, -156.6084, -156.6083, -156.6082, 
    -156.608, -156.608, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6074, -156.6073, -156.6071, -156.6071, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6065, -156.6064, -156.6062, -156.6062, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6085, -156.6084, 
    -156.6082, -156.6082, -156.608, -156.608, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6074, -156.6073, -156.6071, -156.6071, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6065, -156.6064, 
    -156.6062, -156.6062, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6085, -156.6084, -156.6082, -156.6082, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6076, -156.6075, -156.6073, -156.6073, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6067, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6062, -156.6089, -156.6088, 
    -156.6087, -156.6086, -156.6084, -156.6084, -156.6082, -156.6082, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6076, -156.6075, 
    -156.6073, -156.6073, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6067, -156.6066, -156.6064, -156.6064, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6087, -156.6086, -156.6084, -156.6084, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6078, -156.6077, 
    -156.6076, -156.6075, -156.6073, -156.6073, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6067, -156.6066, -156.6064, -156.6064, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6087, -156.6086, 
    -156.6084, -156.6084, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6078, -156.6077, -156.6075, -156.6075, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6069, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6064, -156.6062, -156.6061, -156.6089, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6084, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6078, -156.6077, -156.6075, -156.6075, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6069, -156.6068, 
    -156.6066, -156.6066, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6089, -156.6088, -156.6086, -156.6086, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.608, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6075, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6069, -156.6068, -156.6066, -156.6066, -156.6064, -156.6063, 
    -156.6062, -156.6061, -156.6089, -156.6088, -156.6086, -156.6086, 
    -156.6084, -156.6083, -156.6082, -156.6081, -156.608, -156.6079, 
    -156.6077, -156.6077, -156.6075, -156.6074, -156.6073, -156.6072, 
    -156.6071, -156.607, -156.6068, -156.6068, -156.6066, -156.6066, 
    -156.6064, -156.6063, -156.6062, -156.6061, -156.6088, -156.6088, 
    -156.6086, -156.6086, -156.6084, -156.6083, -156.6082, -156.6081, 
    -156.608, -156.6079, -156.6077, -156.6077, -156.6075, -156.6074, 
    -156.6073, -156.6072, -156.6071, -156.607, -156.6068, -156.6068, 
    -156.6066, -156.6065, -156.6064, -156.6063, -156.6062, -156.6061, 
    -156.6088, -156.6088, -156.6086, -156.6085, -156.6084, -156.6083, 
    -156.6082, -156.6081, -156.6079, -156.6079, -156.6077, -156.6077, 
    -156.6075, -156.6074, -156.6073, -156.6072, -156.6071, -156.607, 
    -156.6068, -156.6068, -156.6066, -156.6065, -156.6064, -156.6063, 
    -156.6062, -156.6061 ;

 lat = 71.27904, 71.27901, 71.27903, 71.27901, 71.27901, 71.27903, 71.27901, 
    71.27903, 71.279, 71.27902, 71.27902, 71.279, 71.27899, 71.27901, 
    71.27901, 71.27899, 71.27899, 71.27901, 71.27898, 71.27901, 71.27901, 
    71.27898, 71.27901, 71.27898, 71.27898, 71.279, 71.27911, 71.27908, 
    71.27911, 71.27908, 71.27908, 71.2791, 71.27908, 71.2791, 71.2791, 
    71.27907, 71.27907, 71.27909, 71.27909, 71.27907, 71.27909, 71.27906, 
    71.27906, 71.27908, 71.27906, 71.27908, 71.27905, 71.27908, 71.27908, 
    71.27905, 71.27908, 71.27905, 71.27915, 71.27918, 71.27915, 71.27917, 
    71.27917, 71.27915, 71.27917, 71.27914, 71.27914, 71.27917, 71.27914, 
    71.27917, 71.27916, 71.27914, 71.27914, 71.27916, 71.27914, 71.27916, 
    71.27913, 71.27915, 71.27913, 71.27915, 71.27915, 71.27912, 71.27914, 
    71.27912, 71.27923, 71.27925, 71.27923, 71.27925, 71.27924, 71.27922, 
    71.27922, 71.27924, 71.27921, 71.27924, 71.27921, 71.27924, 71.27924, 
    71.27921, 71.27921, 71.27923, 71.27923, 71.27921, 71.27923, 71.2792, 
    71.27922, 71.2792, 71.27922, 71.2792, 71.27922, 71.27919, 71.27932, 
    71.2793, 71.2793, 71.27932, 71.2793, 71.27932, 71.27931, 71.27929, 
    71.27929, 71.27931, 71.27931, 71.27928, 71.27928, 71.2793, 71.27928, 
    71.2793, 71.27927, 71.2793, 71.27927, 71.2793, 71.2793, 71.27927, 
    71.27929, 71.27927, 71.27927, 71.27929, 71.27937, 71.2794, 71.27937, 
    71.27939, 71.27939, 71.27937, 71.27937, 71.27939, 71.27938, 71.27936, 
    71.27936, 71.27938, 71.27935, 71.27937, 71.27935, 71.27937, 71.27935, 
    71.27937, 71.27934, 71.27937, 71.27937, 71.27934, 71.27937, 71.27934, 
    71.27934, 71.27936, 71.27944, 71.27946, 71.27946, 71.27944, 71.27946, 
    71.27943, 71.27943, 71.27946, 71.27946, 71.27943, 71.27945, 71.27943, 
    71.27943, 71.27945, 71.27942, 71.27944, 71.27942, 71.27944, 71.27942, 
    71.27944, 71.27943, 71.27941, 71.27943, 71.27941, 71.27943, 71.2794, 
    71.27951, 71.27953, 71.27951, 71.27953, 71.27953, 71.27951, 71.2795, 
    71.27953, 71.27953, 71.2795, 71.27953, 71.2795, 71.2795, 71.27952, 
    71.2795, 71.27952, 71.27949, 71.27951, 71.27949, 71.27951, 71.27951, 
    71.27949, 71.27951, 71.27948, 71.27948, 71.2795, 71.27959, 71.27961, 
    71.27961, 71.27958, 71.2796, 71.27958, 71.27958, 71.2796, 71.2796, 
    71.27957, 71.27957, 71.27959, 71.27957, 71.27959, 71.27959, 71.27956, 
    71.27959, 71.27956, 71.27956, 71.27959, 71.27958, 71.27956, 71.27958, 
    71.27956, 71.27958, 71.27955, 71.27966, 71.27968, 71.27968, 71.27966, 
    71.27968, 71.27965, 71.27967, 71.27965, 71.27967, 71.27965, 71.27967, 
    71.27964, 71.27966, 71.27964, 71.27964, 71.27966, 71.27963, 71.27966, 
    71.27966, 71.27963, 71.27963, 71.27966, 71.27962, 71.27965, 71.27962, 
    71.27965, 71.27973, 71.27975, 71.27975, 71.27972, 71.27975, 71.27972, 
    71.27972, 71.27975, 71.27974, 71.27972, 71.27974, 71.27972, 71.27974, 
    71.27971, 71.27973, 71.27971, 71.27973, 71.27971, 71.27972, 71.2797, 
    71.2797, 71.27972, 71.27972, 71.27969, 71.27972, 71.27969, 71.27982, 
    71.2798, 71.2798, 71.27982, 71.27982, 71.27979, 71.27982, 71.27979, 
    71.27982, 71.27979, 71.27979, 71.27981, 71.27981, 71.27979, 71.27981, 
    71.27978, 71.2798, 71.27978, 71.27978, 71.2798, 71.27977, 71.27979, 
    71.27977, 71.27979, 71.27977, 71.27979, 71.2799, 71.27987, 71.27987, 
    71.27989, 71.27987, 71.27989, 71.27988, 71.27986, 71.27986, 71.27988, 
    71.27988, 71.27985, 71.27988, 71.27985, 71.27985, 71.27988, 71.27988, 
    71.27985, 71.27987, 71.27985, 71.27985, 71.27987, 71.27984, 71.27986, 
    71.27984, 71.27985 ;

 area = 9.902211e-05, 9.902174e-05, 9.902174e-05, 9.902209e-05, 9.902172e-05, 
    9.902208e-05, 9.902207e-05, 9.902169e-05, 9.902168e-05, 9.902204e-05, 
    9.902203e-05, 9.902166e-05, 9.902201e-05, 9.902164e-05, 9.902163e-05, 
    9.902199e-05, 9.902198e-05, 9.902161e-05, 9.902196e-05, 9.902159e-05, 
    9.902158e-05, 9.902194e-05, 9.902156e-05, 9.902192e-05, 9.902155e-05, 
    4.951087e-05, 9.902174e-05, 9.902138e-05, 9.902137e-05, 9.902173e-05, 
    9.902172e-05, 9.902135e-05, 9.90217e-05, 9.902133e-05, 9.902168e-05, 
    9.902132e-05, 9.90213e-05, 9.902166e-05, 9.902164e-05, 9.902128e-05, 
    9.902163e-05, 9.902126e-05, 9.902161e-05, 9.902124e-05, 9.902123e-05, 
    9.902159e-05, 9.902121e-05, 9.902157e-05, 9.902119e-05, 9.902156e-05, 
    9.902118e-05, 9.902155e-05, 9.902102e-05, 9.902138e-05, 9.902137e-05, 
    9.9021e-05, 9.902135e-05, 9.902099e-05, 9.902097e-05, 9.902133e-05, 
    9.902132e-05, 9.902095e-05, 9.90213e-05, 9.902093e-05, 9.902128e-05, 
    9.902092e-05, 9.902126e-05, 9.90209e-05, 9.902124e-05, 9.902088e-05, 
    9.902123e-05, 9.902086e-05, 9.902084e-05, 9.902121e-05, 9.902119e-05, 
    9.902083e-05, 9.902118e-05, 9.902081e-05, 9.902065e-05, 9.902102e-05, 
    9.9021e-05, 9.902064e-05, 9.902099e-05, 9.902062e-05, 9.902097e-05, 
    9.90206e-05, 9.902095e-05, 9.902059e-05, 9.902094e-05, 9.902057e-05, 
    9.902092e-05, 9.902055e-05, 9.902054e-05, 9.90209e-05, 9.902052e-05, 
    9.902088e-05, 9.902086e-05, 9.90205e-05, 9.902048e-05, 9.902084e-05, 
    9.902046e-05, 9.902083e-05, 9.902046e-05, 9.902081e-05, 9.902029e-05, 
    9.902065e-05, 9.902064e-05, 9.902028e-05, 9.902062e-05, 9.902026e-05, 
    9.902024e-05, 9.90206e-05, 9.902059e-05, 9.902022e-05, 9.90202e-05, 
    9.902057e-05, 9.902019e-05, 9.902055e-05, 9.902054e-05, 9.902017e-05, 
    9.902052e-05, 9.902015e-05, 9.902014e-05, 9.90205e-05, 9.902048e-05, 
    9.902012e-05, 9.902046e-05, 9.90201e-05, 9.902046e-05, 9.902009e-05, 
    9.901992e-05, 9.902028e-05, 9.901991e-05, 9.902028e-05, 9.902026e-05, 
    9.901989e-05, 9.901988e-05, 9.902024e-05, 9.902022e-05, 9.901986e-05, 
    9.90202e-05, 9.901984e-05, 9.901982e-05, 9.902019e-05, 9.90198e-05, 
    9.902017e-05, 9.901979e-05, 9.902015e-05, 9.901977e-05, 9.902013e-05, 
    9.902012e-05, 9.901975e-05, 9.90201e-05, 9.901973e-05, 9.901972e-05, 
    9.902009e-05, 9.901955e-05, 9.901992e-05, 9.901991e-05, 9.901955e-05, 
    9.90199e-05, 9.901953e-05, 9.901951e-05, 9.901988e-05, 9.901986e-05, 
    9.901949e-05, 9.901984e-05, 9.901947e-05, 9.901946e-05, 9.901982e-05, 
    9.901944e-05, 9.90198e-05, 9.901942e-05, 9.901979e-05, 9.90194e-05, 
    9.901977e-05, 9.901975e-05, 9.901939e-05, 9.901974e-05, 9.901937e-05, 
    9.901972e-05, 9.901936e-05, 9.901919e-05, 9.901955e-05, 9.901918e-05, 
    9.901955e-05, 9.901953e-05, 9.901916e-05, 9.901915e-05, 9.901951e-05, 
    9.90195e-05, 9.901913e-05, 9.901911e-05, 9.901947e-05, 9.90191e-05, 
    9.901946e-05, 9.901907e-05, 9.901944e-05, 9.901906e-05, 9.901942e-05, 
    9.901904e-05, 9.90194e-05, 9.901939e-05, 9.901902e-05, 9.901937e-05, 
    9.9019e-05, 9.901899e-05, 9.901936e-05, 9.901919e-05, 9.901883e-05, 
    9.901882e-05, 9.901918e-05, 9.90188e-05, 9.901916e-05, 9.901915e-05, 
    9.901878e-05, 9.901877e-05, 9.901913e-05, 9.901911e-05, 9.901875e-05, 
    9.901873e-05, 9.90191e-05, 9.901871e-05, 9.901907e-05, 9.90187e-05, 
    9.901906e-05, 9.901867e-05, 9.901904e-05, 9.901902e-05, 9.901866e-05, 
    9.901901e-05, 9.901864e-05, 9.901863e-05, 9.901899e-05, 9.901846e-05, 
    9.901883e-05, 9.901846e-05, 9.901882e-05, 9.90188e-05, 9.901843e-05, 
    9.901842e-05, 9.901878e-05, 9.90184e-05, 9.901876e-05, 9.901838e-05, 
    9.901875e-05, 9.901873e-05, 9.901836e-05, 9.901835e-05, 9.901871e-05, 
    9.90187e-05, 9.901833e-05, 9.901867e-05, 9.901831e-05, 9.901866e-05, 
    9.90183e-05, 9.901864e-05, 9.901827e-05, 9.901863e-05, 9.901827e-05, 
    9.90181e-05, 9.901846e-05, 9.901809e-05, 9.901846e-05, 9.901843e-05, 
    9.901807e-05, 9.901842e-05, 9.901806e-05, 9.901803e-05, 9.90184e-05, 
    9.901802e-05, 9.901838e-05, 9.901837e-05, 9.9018e-05, 9.901798e-05, 
    9.901835e-05, 9.901797e-05, 9.901833e-05, 9.901795e-05, 9.901831e-05, 
    9.901793e-05, 9.90183e-05, 9.901827e-05, 9.901791e-05, 9.901827e-05, 
    9.90179e-05, 9.90181e-05, 9.901774e-05, 9.901809e-05, 9.901772e-05, 
    9.901771e-05, 9.901807e-05, 9.901769e-05, 9.901806e-05, 9.901803e-05, 
    9.901767e-05, 9.901766e-05, 9.901802e-05, 9.9018e-05, 9.901763e-05, 
    9.901798e-05, 9.901762e-05, 9.90176e-05, 9.901796e-05, 9.901758e-05, 
    9.901795e-05, 9.901757e-05, 9.901793e-05, 9.901791e-05, 9.901755e-05, 
    9.90179e-05, 9.901754e-05, 9.901774e-05, 9.901737e-05, 9.901773e-05, 
    9.901736e-05, 9.901734e-05, 9.901771e-05, 9.901733e-05, 9.901768e-05, 
    9.901731e-05, 9.901767e-05, 9.901766e-05, 9.901728e-05, 9.901727e-05, 
    9.901763e-05, 9.901762e-05, 9.901726e-05, 9.901723e-05, 9.90176e-05, 
    9.901722e-05, 9.901758e-05, 9.901757e-05, 9.90172e-05, 9.901755e-05, 
    9.901718e-05, 9.901718e-05, 9.901754e-05 ;

 topo = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0 ;

 landfrac = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 landmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 pftmask = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1 ;

 ACTUAL_IMMOB =
  5.00767e-14, 5.021391e-14, 5.018725e-14, 5.029783e-14, 5.023652e-14, 
    5.03089e-14, 5.010455e-14, 5.021933e-14, 5.014608e-14, 5.008909e-14, 
    5.051216e-14, 5.030277e-14, 5.072961e-14, 5.059623e-14, 5.093115e-14, 
    5.070883e-14, 5.097595e-14, 5.092479e-14, 5.107884e-14, 5.103473e-14, 
    5.123149e-14, 5.10992e-14, 5.133348e-14, 5.119994e-14, 5.122082e-14, 
    5.109482e-14, 5.034498e-14, 5.048609e-14, 5.03366e-14, 5.035673e-14, 
    5.034771e-14, 5.023776e-14, 5.01823e-14, 5.006624e-14, 5.008733e-14, 
    5.017259e-14, 5.036579e-14, 5.030026e-14, 5.046545e-14, 5.046172e-14, 
    5.064542e-14, 5.056262e-14, 5.08711e-14, 5.07835e-14, 5.103657e-14, 
    5.097296e-14, 5.103357e-14, 5.10152e-14, 5.103381e-14, 5.094051e-14, 
    5.098049e-14, 5.089838e-14, 5.057812e-14, 5.067229e-14, 5.039125e-14, 
    5.022198e-14, 5.010957e-14, 5.002974e-14, 5.004103e-14, 5.006253e-14, 
    5.017309e-14, 5.027701e-14, 5.035615e-14, 5.040906e-14, 5.046119e-14, 
    5.061875e-14, 5.070219e-14, 5.088879e-14, 5.085517e-14, 5.091215e-14, 
    5.096663e-14, 5.105799e-14, 5.104296e-14, 5.108319e-14, 5.091068e-14, 
    5.102534e-14, 5.083601e-14, 5.088781e-14, 5.047519e-14, 5.031795e-14, 
    5.025093e-14, 5.019237e-14, 5.00497e-14, 5.014823e-14, 5.010939e-14, 
    5.020181e-14, 5.026049e-14, 5.023147e-14, 5.041051e-14, 5.034092e-14, 
    5.070713e-14, 5.054949e-14, 5.096027e-14, 5.086208e-14, 5.098381e-14, 
    5.092171e-14, 5.102808e-14, 5.093235e-14, 5.109817e-14, 5.113424e-14, 
    5.110959e-14, 5.12043e-14, 5.092704e-14, 5.103356e-14, 5.023065e-14, 
    5.023538e-14, 5.025744e-14, 5.016046e-14, 5.015453e-14, 5.006566e-14, 
    5.014476e-14, 5.017841e-14, 5.02639e-14, 5.031441e-14, 5.036243e-14, 
    5.046796e-14, 5.058571e-14, 5.075028e-14, 5.086844e-14, 5.094759e-14, 
    5.089907e-14, 5.094191e-14, 5.089402e-14, 5.087157e-14, 5.112071e-14, 
    5.098085e-14, 5.119068e-14, 5.117909e-14, 5.108414e-14, 5.118039e-14, 
    5.023871e-14, 5.021148e-14, 5.011685e-14, 5.019091e-14, 5.005598e-14, 
    5.01315e-14, 5.017489e-14, 5.034234e-14, 5.037914e-14, 5.041322e-14, 
    5.048053e-14, 5.056685e-14, 5.071818e-14, 5.084976e-14, 5.09698e-14, 
    5.096101e-14, 5.096411e-14, 5.09909e-14, 5.092451e-14, 5.100179e-14, 
    5.101474e-14, 5.098085e-14, 5.117753e-14, 5.112137e-14, 5.117884e-14, 
    5.114228e-14, 5.022034e-14, 5.026616e-14, 5.024139e-14, 5.028795e-14, 
    5.025514e-14, 5.040092e-14, 5.044461e-14, 5.064893e-14, 5.056515e-14, 
    5.069851e-14, 5.057871e-14, 5.059994e-14, 5.070279e-14, 5.05852e-14, 
    5.084247e-14, 5.066803e-14, 5.099194e-14, 5.081783e-14, 5.100284e-14, 
    5.096928e-14, 5.102485e-14, 5.107458e-14, 5.113715e-14, 5.125249e-14, 
    5.12258e-14, 5.132223e-14, 5.033446e-14, 5.039384e-14, 5.038864e-14, 
    5.045079e-14, 5.049672e-14, 5.059628e-14, 5.075581e-14, 5.069585e-14, 
    5.080595e-14, 5.082803e-14, 5.066078e-14, 5.076346e-14, 5.043359e-14, 
    5.048689e-14, 5.045518e-14, 5.033913e-14, 5.070963e-14, 5.051957e-14, 
    5.087039e-14, 5.076756e-14, 5.106749e-14, 5.091836e-14, 5.12111e-14, 
    5.133598e-14, 5.145358e-14, 5.159071e-14, 5.042627e-14, 5.038593e-14, 
    5.045818e-14, 5.055804e-14, 5.065073e-14, 5.077382e-14, 5.078643e-14, 
    5.080947e-14, 5.086918e-14, 5.091934e-14, 5.081673e-14, 5.093192e-14, 
    5.049919e-14, 5.072613e-14, 5.037065e-14, 5.047773e-14, 5.055217e-14, 
    5.051955e-14, 5.0689e-14, 5.07289e-14, 5.089095e-14, 5.080722e-14, 
    5.130514e-14, 5.108504e-14, 5.169514e-14, 5.152488e-14, 5.037183e-14, 
    5.042615e-14, 5.061502e-14, 5.052519e-14, 5.078206e-14, 5.084521e-14, 
    5.089656e-14, 5.096212e-14, 5.096922e-14, 5.100806e-14, 5.094441e-14, 
    5.100556e-14, 5.077409e-14, 5.087757e-14, 5.059348e-14, 5.066265e-14, 
    5.063085e-14, 5.059593e-14, 5.070367e-14, 5.081833e-14, 5.082084e-14, 
    5.085757e-14, 5.096097e-14, 5.07831e-14, 5.133343e-14, 5.09937e-14, 
    5.048536e-14, 5.058984e-14, 5.060481e-14, 5.056434e-14, 5.083888e-14, 
    5.073945e-14, 5.100712e-14, 5.093483e-14, 5.105327e-14, 5.099442e-14, 
    5.098576e-14, 5.091016e-14, 5.086305e-14, 5.0744e-14, 5.064708e-14, 
    5.057022e-14, 5.05881e-14, 5.067253e-14, 5.082536e-14, 5.096984e-14, 
    5.09382e-14, 5.104427e-14, 5.076344e-14, 5.088123e-14, 5.08357e-14, 
    5.095441e-14, 5.069424e-14, 5.091566e-14, 5.063758e-14, 5.066199e-14, 
    5.073748e-14, 5.088918e-14, 5.092281e-14, 5.09586e-14, 5.093653e-14, 
    5.082924e-14, 5.081168e-14, 5.073565e-14, 5.071463e-14, 5.065668e-14, 
    5.060867e-14, 5.065253e-14, 5.069856e-14, 5.082931e-14, 5.094702e-14, 
    5.107528e-14, 5.110667e-14, 5.125624e-14, 5.113442e-14, 5.133531e-14, 
    5.116443e-14, 5.146017e-14, 5.092856e-14, 5.115951e-14, 5.074093e-14, 
    5.078609e-14, 5.086768e-14, 5.105478e-14, 5.095385e-14, 5.10719e-14, 
    5.0811e-14, 5.067541e-14, 5.064038e-14, 5.057488e-14, 5.064187e-14, 
    5.063643e-14, 5.07005e-14, 5.067992e-14, 5.083365e-14, 5.075109e-14, 
    5.098553e-14, 5.107098e-14, 5.131211e-14, 5.145971e-14, 5.160989e-14, 
    5.167611e-14, 5.169627e-14, 5.170469e-14 ;

 AGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ALTMAX_LASTYEAR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 AR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_CROP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BAF_PEATF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BCDEP =
  9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 9.571682e-15, 
    9.571682e-15, 9.571682e-15, 9.571682e-15 ;

 BGNPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BTRAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 BUILDHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4PROD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_AERE_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_DIFF_SAT =
  -7.207679e-15, -7.196442e-15, -7.198626e-15, -7.189572e-15, -7.194594e-15, 
    -7.188667e-15, -7.2054e-15, -7.195995e-15, -7.201998e-15, -7.206668e-15, 
    -7.172033e-15, -7.189168e-15, -7.154298e-15, -7.165188e-15, 
    -7.137872e-15, -7.155989e-15, -7.134226e-15, -7.138398e-15, -7.12586e-15, 
    -7.129449e-15, -7.113433e-15, -7.124204e-15, -7.105153e-15, 
    -7.116005e-15, -7.114305e-15, -7.124559e-15, -7.18572e-15, -7.174162e-15, 
    -7.186405e-15, -7.184755e-15, -7.185496e-15, -7.194489e-15, 
    -7.199023e-15, -7.20854e-15, -7.206812e-15, -7.199824e-15, -7.184013e-15, 
    -7.189378e-15, -7.175873e-15, -7.176178e-15, -7.161174e-15, 
    -7.167934e-15, -7.142771e-15, -7.149914e-15, -7.1293e-15, -7.134477e-15, 
    -7.129542e-15, -7.131038e-15, -7.129523e-15, -7.137117e-15, 
    -7.133862e-15, -7.14055e-15, -7.166667e-15, -7.158979e-15, -7.181934e-15, 
    -7.195771e-15, -7.204987e-15, -7.211532e-15, -7.210606e-15, 
    -7.208841e-15, -7.199783e-15, -7.191281e-15, -7.184808e-15, 
    -7.180482e-15, -7.176222e-15, -7.163336e-15, -7.156535e-15, 
    -7.141326e-15, -7.144072e-15, -7.139424e-15, -7.134992e-15, 
    -7.127554e-15, -7.128778e-15, -7.125503e-15, -7.139549e-15, 
    -7.130209e-15, -7.145634e-15, -7.141412e-15, -7.175052e-15, 
    -7.187932e-15, -7.193403e-15, -7.198205e-15, -7.209894e-15, 
    -7.201819e-15, -7.205001e-15, -7.197436e-15, -7.192633e-15, 
    -7.195009e-15, -7.180364e-15, -7.186053e-15, -7.156132e-15, 
    -7.169002e-15, -7.135509e-15, -7.143508e-15, -7.133594e-15, 
    -7.138651e-15, -7.129987e-15, -7.137784e-15, -7.124286e-15, 
    -7.121349e-15, -7.123356e-15, -7.115655e-15, -7.138217e-15, 
    -7.129541e-15, -7.195075e-15, -7.194687e-15, -7.192883e-15, 
    -7.200817e-15, -7.201303e-15, -7.208588e-15, -7.202107e-15, 
    -7.199348e-15, -7.192355e-15, -7.188221e-15, -7.184293e-15, 
    -7.175666e-15, -7.166044e-15, -7.152616e-15, -7.142989e-15, 
    -7.136544e-15, -7.140496e-15, -7.137006e-15, -7.140907e-15, 
    -7.142737e-15, -7.122448e-15, -7.133831e-15, -7.116762e-15, 
    -7.117706e-15, -7.125425e-15, -7.1176e-15, -7.194415e-15, -7.196645e-15, 
    -7.204392e-15, -7.198329e-15, -7.209381e-15, -7.203191e-15, 
    -7.199633e-15, -7.185931e-15, -7.182927e-15, -7.18014e-15, -7.17464e-15, 
    -7.167589e-15, -7.155235e-15, -7.144509e-15, -7.134735e-15, 
    -7.135451e-15, -7.135199e-15, -7.133016e-15, -7.138423e-15, 
    -7.132129e-15, -7.131072e-15, -7.133834e-15, -7.117832e-15, 
    -7.122399e-15, -7.117726e-15, -7.1207e-15, -7.195921e-15, -7.192169e-15, 
    -7.194196e-15, -7.190384e-15, -7.193068e-15, -7.181139e-15, 
    -7.177567e-15, -7.16088e-15, -7.167727e-15, -7.156838e-15, -7.16662e-15, 
    -7.164885e-15, -7.156478e-15, -7.166092e-15, -7.145097e-15, 
    -7.159319e-15, -7.132931e-15, -7.1471e-15, -7.132045e-15, -7.134777e-15, 
    -7.130254e-15, -7.126204e-15, -7.121115e-15, -7.111734e-15, 
    -7.113905e-15, -7.10607e-15, -7.186582e-15, -7.181721e-15, -7.182152e-15, 
    -7.177071e-15, -7.173315e-15, -7.165186e-15, -7.152168e-15, 
    -7.157062e-15, -7.148084e-15, -7.146282e-15, -7.159924e-15, 
    -7.151542e-15, -7.178473e-15, -7.174112e-15, -7.176709e-15, 
    -7.186196e-15, -7.15593e-15, -7.171443e-15, -7.14283e-15, -7.151212e-15, 
    -7.126781e-15, -7.138916e-15, -7.1151e-15, -7.104942e-15, -7.095408e-15, 
    -7.084272e-15, -7.179073e-15, -7.182374e-15, -7.176467e-15, 
    -7.168302e-15, -7.160741e-15, -7.1507e-15, -7.149675e-15, -7.147795e-15, 
    -7.142931e-15, -7.138844e-15, -7.147198e-15, -7.13782e-15, -7.173095e-15, 
    -7.154587e-15, -7.18362e-15, -7.174859e-15, -7.168784e-15, -7.171451e-15, 
    -7.157622e-15, -7.154366e-15, -7.141152e-15, -7.147981e-15, 
    -7.107445e-15, -7.125345e-15, -7.075816e-15, -7.089614e-15, 
    -7.183526e-15, -7.179085e-15, -7.163652e-15, -7.170991e-15, 
    -7.150031e-15, -7.144881e-15, -7.1407e-15, -7.135356e-15, -7.134781e-15, 
    -7.131618e-15, -7.136802e-15, -7.131823e-15, -7.150678e-15, 
    -7.142245e-15, -7.165417e-15, -7.159768e-15, -7.162367e-15, 
    -7.165217e-15, -7.156424e-15, -7.147066e-15, -7.14687e-15, -7.143872e-15, 
    -7.135423e-15, -7.149947e-15, -7.105132e-15, -7.132763e-15, 
    -7.174247e-15, -7.165704e-15, -7.164489e-15, -7.167795e-15, 
    -7.145397e-15, -7.153503e-15, -7.131696e-15, -7.137582e-15, 
    -7.127941e-15, -7.13273e-15, -7.133435e-15, -7.139592e-15, -7.143428e-15, 
    -7.153131e-15, -7.161038e-15, -7.167317e-15, -7.165856e-15, 
    -7.158961e-15, -7.146495e-15, -7.134728e-15, -7.137303e-15, 
    -7.128672e-15, -7.151548e-15, -7.141944e-15, -7.145653e-15, 
    -7.135987e-15, -7.15719e-15, -7.139118e-15, -7.161817e-15, -7.159825e-15, 
    -7.153664e-15, -7.14129e-15, -7.138562e-15, -7.135643e-15, -7.137444e-15, 
    -7.14618e-15, -7.147614e-15, -7.153815e-15, -7.155527e-15, -7.160258e-15, 
    -7.164177e-15, -7.160595e-15, -7.156836e-15, -7.146177e-15, 
    -7.136585e-15, -7.126146e-15, -7.123595e-15, -7.111416e-15, 
    -7.121324e-15, -7.104977e-15, -7.118864e-15, -7.09485e-15, -7.138078e-15, 
    -7.119281e-15, -7.153386e-15, -7.149703e-15, -7.143044e-15, 
    -7.127807e-15, -7.136032e-15, -7.126416e-15, -7.14767e-15, -7.158721e-15, 
    -7.161588e-15, -7.166934e-15, -7.161466e-15, -7.161911e-15, 
    -7.156683e-15, -7.158363e-15, -7.145824e-15, -7.152556e-15, 
    -7.133451e-15, -7.126492e-15, -7.106889e-15, -7.094901e-15, 
    -7.082729e-15, -7.077361e-15, -7.075728e-15, -7.075046e-15 ;

 CH4_SURF_DIFF_UNSAT =
  1.579902e-14, 1.537487e-14, 1.545734e-14, 1.511517e-14, 1.5305e-14, 
    1.508093e-14, 1.571304e-14, 1.535802e-14, 1.558467e-14, 1.576085e-14, 
    1.445096e-14, 1.509991e-14, 1.377671e-14, 1.419076e-14, 1.315047e-14, 
    1.384113e-14, 1.301117e-14, 1.317042e-14, 1.269112e-14, 1.282845e-14, 
    1.221515e-14, 1.262773e-14, 1.189716e-14, 1.231371e-14, 1.224855e-14, 
    1.264134e-14, 1.496936e-14, 1.453175e-14, 1.499527e-14, 1.493288e-14, 
    1.496088e-14, 1.530107e-14, 1.547246e-14, 1.583145e-14, 1.576628e-14, 
    1.550263e-14, 1.490482e-14, 1.510779e-14, 1.459628e-14, 1.460783e-14, 
    1.403819e-14, 1.429505e-14, 1.333734e-14, 1.36096e-14, 1.282272e-14, 
    1.302065e-14, 1.283201e-14, 1.288922e-14, 1.283127e-14, 1.312154e-14, 
    1.299718e-14, 1.325259e-14, 1.424694e-14, 1.395476e-14, 1.482602e-14, 
    1.534967e-14, 1.569747e-14, 1.594422e-14, 1.590934e-14, 1.584283e-14, 
    1.550108e-14, 1.517974e-14, 1.493481e-14, 1.477096e-14, 1.460949e-14, 
    1.41206e-14, 1.386184e-14, 1.328226e-14, 1.33869e-14, 1.320965e-14, 
    1.304034e-14, 1.2756e-14, 1.28028e-14, 1.267751e-14, 1.321435e-14, 
    1.285758e-14, 1.344649e-14, 1.328544e-14, 1.456551e-14, 1.505304e-14, 
    1.526015e-14, 1.544148e-14, 1.588251e-14, 1.557795e-14, 1.569802e-14, 
    1.541238e-14, 1.523086e-14, 1.532064e-14, 1.476647e-14, 1.498194e-14, 
    1.384651e-14, 1.433567e-14, 1.306009e-14, 1.336542e-14, 1.298689e-14, 
    1.318007e-14, 1.284906e-14, 1.314697e-14, 1.263089e-14, 1.251847e-14, 
    1.259529e-14, 1.230021e-14, 1.316348e-14, 1.283201e-14, 1.532315e-14, 
    1.530851e-14, 1.52403e-14, 1.554013e-14, 1.555847e-14, 1.583323e-14, 
    1.558876e-14, 1.548464e-14, 1.522034e-14, 1.506397e-14, 1.491533e-14, 
    1.458846e-14, 1.422331e-14, 1.371262e-14, 1.334563e-14, 1.309958e-14, 
    1.325047e-14, 1.311725e-14, 1.326617e-14, 1.333596e-14, 1.256059e-14, 
    1.299602e-14, 1.234266e-14, 1.237882e-14, 1.267453e-14, 1.237475e-14, 
    1.529823e-14, 1.538249e-14, 1.5675e-14, 1.544609e-14, 1.586315e-14, 
    1.56297e-14, 1.549545e-14, 1.497741e-14, 1.48636e-14, 1.475803e-14, 
    1.454953e-14, 1.428191e-14, 1.381232e-14, 1.340365e-14, 1.303049e-14, 
    1.305784e-14, 1.304821e-14, 1.296483e-14, 1.317135e-14, 1.293092e-14, 
    1.289056e-14, 1.299608e-14, 1.238367e-14, 1.255866e-14, 1.237959e-14, 
    1.249353e-14, 1.535511e-14, 1.521332e-14, 1.528993e-14, 1.514586e-14, 
    1.524736e-14, 1.479597e-14, 1.466061e-14, 1.402714e-14, 1.428717e-14, 
    1.387334e-14, 1.424514e-14, 1.417926e-14, 1.38598e-14, 1.422506e-14, 
    1.342616e-14, 1.39678e-14, 1.296159e-14, 1.350259e-14, 1.292768e-14, 
    1.30321e-14, 1.285921e-14, 1.270433e-14, 1.250948e-14, 1.214985e-14, 
    1.223314e-14, 1.193234e-14, 1.500193e-14, 1.481799e-14, 1.48342e-14, 
    1.464169e-14, 1.449931e-14, 1.419067e-14, 1.369552e-14, 1.388174e-14, 
    1.353987e-14, 1.347123e-14, 1.399061e-14, 1.367172e-14, 1.469488e-14, 
    1.45296e-14, 1.462802e-14, 1.498741e-14, 1.383881e-14, 1.442836e-14, 
    1.333956e-14, 1.365907e-14, 1.272641e-14, 1.31903e-14, 1.227898e-14, 
    1.188916e-14, 1.152225e-14, 1.109323e-14, 1.471761e-14, 1.48426e-14, 
    1.46188e-14, 1.430909e-14, 1.402172e-14, 1.363958e-14, 1.360048e-14, 
    1.352888e-14, 1.33434e-14, 1.318742e-14, 1.350622e-14, 1.314832e-14, 
    1.449123e-14, 1.378763e-14, 1.488984e-14, 1.455799e-14, 1.432735e-14, 
    1.442855e-14, 1.390303e-14, 1.377914e-14, 1.327559e-14, 1.353593e-14, 
    1.198537e-14, 1.267159e-14, 1.076651e-14, 1.12992e-14, 1.488627e-14, 
    1.471804e-14, 1.413242e-14, 1.441109e-14, 1.361407e-14, 1.341782e-14, 
    1.325828e-14, 1.305429e-14, 1.303227e-14, 1.291139e-14, 1.310947e-14, 
    1.291922e-14, 1.363877e-14, 1.331726e-14, 1.419939e-14, 1.398472e-14, 
    1.408349e-14, 1.41918e-14, 1.385748e-14, 1.35012e-14, 1.349361e-14, 
    1.337934e-14, 1.305726e-14, 1.361085e-14, 1.189672e-14, 1.295552e-14, 
    1.453459e-14, 1.421045e-14, 1.416418e-14, 1.428975e-14, 1.34375e-14, 
    1.374635e-14, 1.291434e-14, 1.313926e-14, 1.277073e-14, 1.295387e-14, 
    1.298081e-14, 1.321599e-14, 1.336238e-14, 1.373218e-14, 1.403301e-14, 
    1.427154e-14, 1.421608e-14, 1.395405e-14, 1.347941e-14, 1.303027e-14, 
    1.312866e-14, 1.279874e-14, 1.367188e-14, 1.33058e-14, 1.344729e-14, 
    1.307834e-14, 1.388668e-14, 1.319828e-14, 1.406259e-14, 1.398683e-14, 
    1.375248e-14, 1.328095e-14, 1.317665e-14, 1.306523e-14, 1.313399e-14, 
    1.346736e-14, 1.352198e-14, 1.375818e-14, 1.382338e-14, 1.400333e-14, 
    1.415228e-14, 1.401618e-14, 1.387323e-14, 1.346723e-14, 1.310124e-14, 
    1.270212e-14, 1.260444e-14, 1.213786e-14, 1.251765e-14, 1.189082e-14, 
    1.242371e-14, 1.150113e-14, 1.315842e-14, 1.243943e-14, 1.374182e-14, 
    1.360157e-14, 1.334784e-14, 1.276579e-14, 1.308008e-14, 1.271252e-14, 
    1.352412e-14, 1.3945e-14, 1.405391e-14, 1.425703e-14, 1.404927e-14, 
    1.406617e-14, 1.386733e-14, 1.393123e-14, 1.345375e-14, 1.371025e-14, 
    1.298148e-14, 1.271543e-14, 1.196385e-14, 1.150287e-14, 1.103348e-14, 
    1.082618e-14, 1.076308e-14, 1.073669e-14 ;

 CH4_SURF_EBUL_SAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CH4_SURF_EBUL_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_CTRUNC =
  1.931953e-23, 1.931952e-23, 1.931953e-23, 1.931952e-23, 1.931952e-23, 
    1.931952e-23, 1.931953e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 
    1.93195e-23, 1.931952e-23, 1.931949e-23, 1.93195e-23, 1.931947e-23, 
    1.931949e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 
    1.931945e-23, 1.931946e-23, 1.931944e-23, 1.931945e-23, 1.931945e-23, 
    1.931946e-23, 1.931951e-23, 1.93195e-23, 1.931951e-23, 1.931951e-23, 
    1.931951e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931951e-23, 1.931952e-23, 1.93195e-23, 1.93195e-23, 
    1.931949e-23, 1.93195e-23, 1.931948e-23, 1.931948e-23, 1.931946e-23, 
    1.931947e-23, 1.931946e-23, 1.931947e-23, 1.931946e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.93195e-23, 1.931949e-23, 1.931951e-23, 
    1.931952e-23, 1.931953e-23, 1.931954e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931952e-23, 1.931951e-23, 1.931951e-23, 1.93195e-23, 
    1.931949e-23, 1.931949e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931946e-23, 1.931947e-23, 
    1.931947e-23, 1.931948e-23, 1.931947e-23, 1.93195e-23, 1.931952e-23, 
    1.931952e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931952e-23, 1.931952e-23, 1.931952e-23, 1.931951e-23, 1.931951e-23, 
    1.931949e-23, 1.93195e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 
    1.931946e-23, 1.931945e-23, 1.931947e-23, 1.931946e-23, 1.931952e-23, 
    1.931952e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931953e-23, 1.931952e-23, 1.931952e-23, 1.931951e-23, 
    1.93195e-23, 1.93195e-23, 1.931948e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931946e-23, 
    1.931947e-23, 1.931945e-23, 1.931945e-23, 1.931946e-23, 1.931945e-23, 
    1.931952e-23, 1.931952e-23, 1.931953e-23, 1.931953e-23, 1.931953e-23, 
    1.931953e-23, 1.931953e-23, 1.931951e-23, 1.931951e-23, 1.931951e-23, 
    1.93195e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931945e-23, 1.931946e-23, 1.931945e-23, 
    1.931946e-23, 1.931952e-23, 1.931952e-23, 1.931952e-23, 1.931952e-23, 
    1.931952e-23, 1.931951e-23, 1.931951e-23, 1.931949e-23, 1.93195e-23, 
    1.931949e-23, 1.93195e-23, 1.93195e-23, 1.931949e-23, 1.93195e-23, 
    1.931948e-23, 1.931949e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931946e-23, 1.931945e-23, 
    1.931945e-23, 1.931944e-23, 1.931951e-23, 1.931951e-23, 1.931951e-23, 
    1.931951e-23, 1.93195e-23, 1.93195e-23, 1.931948e-23, 1.931949e-23, 
    1.931948e-23, 1.931948e-23, 1.931949e-23, 1.931948e-23, 1.931951e-23, 
    1.93195e-23, 1.931951e-23, 1.931951e-23, 1.931949e-23, 1.93195e-23, 
    1.931948e-23, 1.931948e-23, 1.931946e-23, 1.931947e-23, 1.931945e-23, 
    1.931944e-23, 1.931943e-23, 1.931942e-23, 1.931951e-23, 1.931951e-23, 
    1.931951e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931948e-23, 1.931948e-23, 1.931947e-23, 1.931948e-23, 1.931947e-23, 
    1.93195e-23, 1.931949e-23, 1.931951e-23, 1.93195e-23, 1.93195e-23, 
    1.93195e-23, 1.931949e-23, 1.931949e-23, 1.931947e-23, 1.931948e-23, 
    1.931944e-23, 1.931946e-23, 1.931942e-23, 1.931943e-23, 1.931951e-23, 
    1.931951e-23, 1.931949e-23, 1.93195e-23, 1.931948e-23, 1.931948e-23, 
    1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931947e-23, 1.931948e-23, 1.931948e-23, 1.93195e-23, 1.931949e-23, 
    1.931949e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931948e-23, 1.931947e-23, 1.931948e-23, 1.931944e-23, 1.931947e-23, 
    1.93195e-23, 1.93195e-23, 1.93195e-23, 1.93195e-23, 1.931948e-23, 
    1.931949e-23, 1.931947e-23, 1.931947e-23, 1.931946e-23, 1.931947e-23, 
    1.931947e-23, 1.931947e-23, 1.931948e-23, 1.931949e-23, 1.931949e-23, 
    1.93195e-23, 1.93195e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 
    1.931947e-23, 1.931946e-23, 1.931948e-23, 1.931947e-23, 1.931948e-23, 
    1.931947e-23, 1.931949e-23, 1.931947e-23, 1.931949e-23, 1.931949e-23, 
    1.931949e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 1.931947e-23, 
    1.931948e-23, 1.931948e-23, 1.931949e-23, 1.931949e-23, 1.931949e-23, 
    1.93195e-23, 1.931949e-23, 1.931949e-23, 1.931948e-23, 1.931947e-23, 
    1.931946e-23, 1.931946e-23, 1.931945e-23, 1.931946e-23, 1.931944e-23, 
    1.931945e-23, 1.931943e-23, 1.931947e-23, 1.931946e-23, 1.931949e-23, 
    1.931948e-23, 1.931948e-23, 1.931946e-23, 1.931947e-23, 1.931946e-23, 
    1.931948e-23, 1.931949e-23, 1.931949e-23, 1.93195e-23, 1.931949e-23, 
    1.931949e-23, 1.931949e-23, 1.931949e-23, 1.931948e-23, 1.931948e-23, 
    1.931947e-23, 1.931946e-23, 1.931944e-23, 1.931943e-23, 1.931942e-23, 
    1.931942e-23, 1.931942e-23, 1.931942e-23 ;

 COL_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 COL_NTRUNC =
  1.975388e-24, 1.975387e-24, 1.975387e-24, 1.975386e-24, 1.975386e-24, 
    1.975386e-24, 1.975388e-24, 1.975387e-24, 1.975387e-24, 1.975388e-24, 
    1.975384e-24, 1.975386e-24, 1.975381e-24, 1.975383e-24, 1.975379e-24, 
    1.975382e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975379e-24, 
    1.975376e-24, 1.975378e-24, 1.975375e-24, 1.975377e-24, 1.975377e-24, 
    1.975378e-24, 1.975385e-24, 1.975384e-24, 1.975385e-24, 1.975385e-24, 
    1.975385e-24, 1.975386e-24, 1.975387e-24, 1.975388e-24, 1.975388e-24, 
    1.975387e-24, 1.975385e-24, 1.975386e-24, 1.975384e-24, 1.975384e-24, 
    1.975382e-24, 1.975383e-24, 1.97538e-24, 1.975381e-24, 1.975378e-24, 
    1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.97538e-24, 1.975383e-24, 1.975382e-24, 1.975385e-24, 
    1.975387e-24, 1.975388e-24, 1.975388e-24, 1.975388e-24, 1.975388e-24, 
    1.975387e-24, 1.975386e-24, 1.975385e-24, 1.975385e-24, 1.975384e-24, 
    1.975383e-24, 1.975382e-24, 1.97538e-24, 1.97538e-24, 1.97538e-24, 
    1.975379e-24, 1.975378e-24, 1.975378e-24, 1.975378e-24, 1.97538e-24, 
    1.975379e-24, 1.97538e-24, 1.97538e-24, 1.975384e-24, 1.975386e-24, 
    1.975386e-24, 1.975387e-24, 1.975388e-24, 1.975387e-24, 1.975388e-24, 
    1.975387e-24, 1.975386e-24, 1.975386e-24, 1.975385e-24, 1.975385e-24, 
    1.975382e-24, 1.975383e-24, 1.975379e-24, 1.97538e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975377e-24, 
    1.975378e-24, 1.975377e-24, 1.975379e-24, 1.975379e-24, 1.975386e-24, 
    1.975386e-24, 1.975386e-24, 1.975387e-24, 1.975387e-24, 1.975388e-24, 
    1.975387e-24, 1.975387e-24, 1.975386e-24, 1.975386e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975381e-24, 1.97538e-24, 1.975379e-24, 
    1.97538e-24, 1.975379e-24, 1.97538e-24, 1.97538e-24, 1.975378e-24, 
    1.975379e-24, 1.975377e-24, 1.975377e-24, 1.975378e-24, 1.975377e-24, 
    1.975386e-24, 1.975387e-24, 1.975388e-24, 1.975387e-24, 1.975388e-24, 
    1.975387e-24, 1.975387e-24, 1.975385e-24, 1.975385e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975382e-24, 1.97538e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975377e-24, 1.975378e-24, 1.975377e-24, 
    1.975377e-24, 1.975387e-24, 1.975386e-24, 1.975386e-24, 1.975386e-24, 
    1.975386e-24, 1.975385e-24, 1.975384e-24, 1.975382e-24, 1.975383e-24, 
    1.975382e-24, 1.975383e-24, 1.975383e-24, 1.975382e-24, 1.975383e-24, 
    1.97538e-24, 1.975382e-24, 1.975379e-24, 1.975381e-24, 1.975379e-24, 
    1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975377e-24, 1.975376e-24, 
    1.975377e-24, 1.975376e-24, 1.975385e-24, 1.975385e-24, 1.975385e-24, 
    1.975384e-24, 1.975384e-24, 1.975383e-24, 1.975381e-24, 1.975382e-24, 
    1.975381e-24, 1.97538e-24, 1.975382e-24, 1.975381e-24, 1.975384e-24, 
    1.975384e-24, 1.975384e-24, 1.975385e-24, 1.975382e-24, 1.975384e-24, 
    1.97538e-24, 1.975381e-24, 1.975378e-24, 1.975379e-24, 1.975377e-24, 
    1.975375e-24, 1.975374e-24, 1.975373e-24, 1.975384e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975382e-24, 1.975381e-24, 1.975381e-24, 
    1.975381e-24, 1.97538e-24, 1.975379e-24, 1.975381e-24, 1.975379e-24, 
    1.975384e-24, 1.975381e-24, 1.975385e-24, 1.975384e-24, 1.975383e-24, 
    1.975384e-24, 1.975382e-24, 1.975381e-24, 1.97538e-24, 1.975381e-24, 
    1.975376e-24, 1.975378e-24, 1.975372e-24, 1.975373e-24, 1.975385e-24, 
    1.975384e-24, 1.975383e-24, 1.975383e-24, 1.975381e-24, 1.97538e-24, 
    1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.975379e-24, 1.975381e-24, 1.97538e-24, 1.975383e-24, 1.975382e-24, 
    1.975382e-24, 1.975383e-24, 1.975382e-24, 1.975381e-24, 1.97538e-24, 
    1.97538e-24, 1.975379e-24, 1.975381e-24, 1.975375e-24, 1.975379e-24, 
    1.975384e-24, 1.975383e-24, 1.975383e-24, 1.975383e-24, 1.97538e-24, 
    1.975381e-24, 1.975379e-24, 1.975379e-24, 1.975378e-24, 1.975379e-24, 
    1.975379e-24, 1.97538e-24, 1.97538e-24, 1.975381e-24, 1.975382e-24, 
    1.975383e-24, 1.975383e-24, 1.975382e-24, 1.97538e-24, 1.975379e-24, 
    1.975379e-24, 1.975378e-24, 1.975381e-24, 1.97538e-24, 1.97538e-24, 
    1.975379e-24, 1.975382e-24, 1.97538e-24, 1.975382e-24, 1.975382e-24, 
    1.975381e-24, 1.97538e-24, 1.975379e-24, 1.975379e-24, 1.975379e-24, 
    1.97538e-24, 1.975381e-24, 1.975381e-24, 1.975382e-24, 1.975382e-24, 
    1.975383e-24, 1.975382e-24, 1.975382e-24, 1.97538e-24, 1.975379e-24, 
    1.975378e-24, 1.975378e-24, 1.975376e-24, 1.975377e-24, 1.975375e-24, 
    1.975377e-24, 1.975374e-24, 1.975379e-24, 1.975377e-24, 1.975381e-24, 
    1.975381e-24, 1.97538e-24, 1.975378e-24, 1.975379e-24, 1.975378e-24, 
    1.975381e-24, 1.975382e-24, 1.975382e-24, 1.975383e-24, 1.975382e-24, 
    1.975382e-24, 1.975382e-24, 1.975382e-24, 1.97538e-24, 1.975381e-24, 
    1.975379e-24, 1.975378e-24, 1.975376e-24, 1.975374e-24, 1.975373e-24, 
    1.975372e-24, 1.975372e-24, 1.975372e-24 ;

 CONC_CH4_SAT =
  3.297007e-08, 3.294845e-08, 3.295266e-08, 3.293521e-08, 3.29449e-08, 
    3.293347e-08, 3.29657e-08, 3.294758e-08, 3.295916e-08, 3.296815e-08, 
    3.290132e-08, 3.293444e-08, 3.286712e-08, 3.288819e-08, 3.283536e-08, 
    3.287038e-08, 3.282831e-08, 3.28364e-08, 3.281214e-08, 3.281909e-08, 
    3.278798e-08, 3.280892e-08, 3.277194e-08, 3.2793e-08, 3.278969e-08, 
    3.280961e-08, 3.292781e-08, 3.290543e-08, 3.292912e-08, 3.292593e-08, 
    3.292737e-08, 3.294469e-08, 3.295339e-08, 3.297176e-08, 3.296843e-08, 
    3.295496e-08, 3.29245e-08, 3.293486e-08, 3.290883e-08, 3.290942e-08, 
    3.288044e-08, 3.28935e-08, 3.284487e-08, 3.285869e-08, 3.28188e-08, 
    3.282882e-08, 3.281926e-08, 3.282216e-08, 3.281922e-08, 3.283392e-08, 
    3.282762e-08, 3.284057e-08, 3.289105e-08, 3.287619e-08, 3.29205e-08, 
    3.294712e-08, 3.296491e-08, 3.29775e-08, 3.297572e-08, 3.297232e-08, 
    3.295488e-08, 3.293853e-08, 3.292606e-08, 3.291771e-08, 3.29095e-08, 
    3.288456e-08, 3.287145e-08, 3.284205e-08, 3.284739e-08, 3.283838e-08, 
    3.282982e-08, 3.281541e-08, 3.281778e-08, 3.281143e-08, 3.283864e-08, 
    3.282054e-08, 3.285042e-08, 3.284224e-08, 3.290714e-08, 3.293207e-08, 
    3.294256e-08, 3.295185e-08, 3.297435e-08, 3.29588e-08, 3.296493e-08, 
    3.295039e-08, 3.294113e-08, 3.294571e-08, 3.291749e-08, 3.292845e-08, 
    3.287067e-08, 3.289555e-08, 3.283082e-08, 3.28463e-08, 3.282711e-08, 
    3.28369e-08, 3.282011e-08, 3.283523e-08, 3.280908e-08, 3.280337e-08, 
    3.280726e-08, 3.279235e-08, 3.283606e-08, 3.281925e-08, 3.294583e-08, 
    3.294508e-08, 3.294162e-08, 3.295687e-08, 3.295781e-08, 3.297184e-08, 
    3.295937e-08, 3.295405e-08, 3.29406e-08, 3.293263e-08, 3.292506e-08, 
    3.290842e-08, 3.288983e-08, 3.286389e-08, 3.284529e-08, 3.283283e-08, 
    3.284048e-08, 3.283372e-08, 3.284127e-08, 3.284481e-08, 3.28055e-08, 
    3.282756e-08, 3.279449e-08, 3.279633e-08, 3.281127e-08, 3.279612e-08, 
    3.294456e-08, 3.294886e-08, 3.296376e-08, 3.295211e-08, 3.297337e-08, 
    3.296145e-08, 3.295458e-08, 3.29282e-08, 3.292243e-08, 3.291705e-08, 
    3.290645e-08, 3.289283e-08, 3.286896e-08, 3.284822e-08, 3.282933e-08, 
    3.283071e-08, 3.283022e-08, 3.282599e-08, 3.283646e-08, 3.282427e-08, 
    3.282221e-08, 3.282758e-08, 3.279657e-08, 3.280542e-08, 3.279636e-08, 
    3.280213e-08, 3.294747e-08, 3.294024e-08, 3.294414e-08, 3.293679e-08, 
    3.294196e-08, 3.291895e-08, 3.291205e-08, 3.287985e-08, 3.289309e-08, 
    3.287205e-08, 3.289097e-08, 3.288761e-08, 3.287131e-08, 3.288995e-08, 
    3.284934e-08, 3.287682e-08, 3.282582e-08, 3.285319e-08, 3.282411e-08, 
    3.282941e-08, 3.282065e-08, 3.281279e-08, 3.280293e-08, 3.278472e-08, 
    3.278894e-08, 3.277373e-08, 3.292947e-08, 3.292009e-08, 3.292094e-08, 
    3.291114e-08, 3.290388e-08, 3.28882e-08, 3.286304e-08, 3.287251e-08, 
    3.285516e-08, 3.285166e-08, 3.287804e-08, 3.286182e-08, 3.291382e-08, 
    3.290539e-08, 3.291043e-08, 3.292872e-08, 3.287029e-08, 3.290024e-08, 
    3.284498e-08, 3.286119e-08, 3.281391e-08, 3.283739e-08, 3.279126e-08, 
    3.27715e-08, 3.275303e-08, 3.273132e-08, 3.291499e-08, 3.292137e-08, 
    3.290998e-08, 3.289418e-08, 3.28796e-08, 3.28602e-08, 3.285823e-08, 
    3.285459e-08, 3.284519e-08, 3.283728e-08, 3.285341e-08, 3.28353e-08, 
    3.290338e-08, 3.28677e-08, 3.292375e-08, 3.290683e-08, 3.289512e-08, 
    3.290029e-08, 3.287359e-08, 3.28673e-08, 3.284172e-08, 3.285496e-08, 
    3.277635e-08, 3.281109e-08, 3.271488e-08, 3.274172e-08, 3.292359e-08, 
    3.291503e-08, 3.288521e-08, 3.28994e-08, 3.285892e-08, 3.284895e-08, 
    3.284087e-08, 3.283051e-08, 3.282941e-08, 3.282328e-08, 3.283333e-08, 
    3.282369e-08, 3.286016e-08, 3.284386e-08, 3.288865e-08, 3.287773e-08, 
    3.288276e-08, 3.288827e-08, 3.287128e-08, 3.285315e-08, 3.285281e-08, 
    3.284699e-08, 3.283053e-08, 3.285875e-08, 3.277179e-08, 3.282539e-08, 
    3.290569e-08, 3.288916e-08, 3.288685e-08, 3.289324e-08, 3.284995e-08, 
    3.286562e-08, 3.282343e-08, 3.283484e-08, 3.281616e-08, 3.282544e-08, 
    3.28268e-08, 3.283873e-08, 3.284614e-08, 3.28649e-08, 3.288018e-08, 
    3.289232e-08, 3.28895e-08, 3.287616e-08, 3.285205e-08, 3.282929e-08, 
    3.283427e-08, 3.281758e-08, 3.286185e-08, 3.284326e-08, 3.285043e-08, 
    3.283174e-08, 3.287275e-08, 3.28377e-08, 3.28817e-08, 3.287785e-08, 
    3.286593e-08, 3.284197e-08, 3.283673e-08, 3.283107e-08, 3.283457e-08, 
    3.285145e-08, 3.285423e-08, 3.286623e-08, 3.286953e-08, 3.287869e-08, 
    3.288626e-08, 3.287933e-08, 3.287206e-08, 3.285146e-08, 3.283289e-08, 
    3.281267e-08, 3.280774e-08, 3.278404e-08, 3.280328e-08, 3.277149e-08, 
    3.279843e-08, 3.275185e-08, 3.283573e-08, 3.27993e-08, 3.28654e-08, 
    3.285829e-08, 3.284537e-08, 3.281586e-08, 3.283183e-08, 3.281317e-08, 
    3.285435e-08, 3.287568e-08, 3.288126e-08, 3.289157e-08, 3.288102e-08, 
    3.288188e-08, 3.287178e-08, 3.287503e-08, 3.285077e-08, 3.28638e-08, 
    3.282682e-08, 3.281333e-08, 3.277531e-08, 3.2752e-08, 3.272836e-08, 
    3.271791e-08, 3.271473e-08, 3.27134e-08,
  5.410123e-11, 5.412475e-11, 5.412022e-11, 5.413908e-11, 5.412868e-11, 
    5.414098e-11, 5.410608e-11, 5.412562e-11, 5.411319e-11, 5.410345e-11, 
    5.41754e-11, 5.413994e-11, 5.421283e-11, 5.419017e-11, 5.424724e-11, 
    5.420921e-11, 5.425493e-11, 5.424631e-11, 5.427263e-11, 5.42651e-11, 
    5.429836e-11, 5.42761e-11, 5.431584e-11, 5.429314e-11, 5.429663e-11, 
    5.427534e-11, 5.414724e-11, 5.417094e-11, 5.41458e-11, 5.414919e-11, 
    5.41477e-11, 5.412884e-11, 5.411922e-11, 5.409954e-11, 5.410315e-11, 
    5.411766e-11, 5.415072e-11, 5.413961e-11, 5.41679e-11, 5.416727e-11, 
    5.419859e-11, 5.418447e-11, 5.423715e-11, 5.422223e-11, 5.426542e-11, 
    5.425455e-11, 5.426488e-11, 5.426177e-11, 5.426492e-11, 5.424898e-11, 
    5.42558e-11, 5.424182e-11, 5.418709e-11, 5.420315e-11, 5.415512e-11, 
    5.412593e-11, 5.410691e-11, 5.409327e-11, 5.40952e-11, 5.409884e-11, 
    5.411774e-11, 5.413563e-11, 5.41492e-11, 5.415824e-11, 5.416717e-11, 
    5.419375e-11, 5.420815e-11, 5.424008e-11, 5.423446e-11, 5.424408e-11, 
    5.425347e-11, 5.426903e-11, 5.426649e-11, 5.42733e-11, 5.424393e-11, 
    5.426341e-11, 5.423123e-11, 5.424002e-11, 5.416905e-11, 5.414263e-11, 
    5.413092e-11, 5.412107e-11, 5.409667e-11, 5.411349e-11, 5.410685e-11, 
    5.412277e-11, 5.41328e-11, 5.412786e-11, 5.415849e-11, 5.414657e-11, 
    5.4209e-11, 5.418215e-11, 5.425238e-11, 5.423563e-11, 5.425641e-11, 
    5.424583e-11, 5.42639e-11, 5.424764e-11, 5.427589e-11, 5.428196e-11, 
    5.42778e-11, 5.429398e-11, 5.424673e-11, 5.426483e-11, 5.41277e-11, 
    5.41285e-11, 5.41323e-11, 5.411558e-11, 5.411459e-11, 5.409942e-11, 
    5.411297e-11, 5.411869e-11, 5.413342e-11, 5.414202e-11, 5.415023e-11, 
    5.416828e-11, 5.418831e-11, 5.421644e-11, 5.423671e-11, 5.425025e-11, 
    5.424198e-11, 5.424928e-11, 5.42411e-11, 5.423729e-11, 5.427965e-11, 
    5.425583e-11, 5.429165e-11, 5.428969e-11, 5.427345e-11, 5.428992e-11, 
    5.412907e-11, 5.412444e-11, 5.410817e-11, 5.41209e-11, 5.409777e-11, 
    5.411066e-11, 5.411802e-11, 5.41467e-11, 5.415313e-11, 5.415891e-11, 
    5.417046e-11, 5.418519e-11, 5.421098e-11, 5.423346e-11, 5.425404e-11, 
    5.425254e-11, 5.425306e-11, 5.42576e-11, 5.424629e-11, 5.425946e-11, 
    5.426162e-11, 5.425589e-11, 5.428943e-11, 5.427986e-11, 5.428965e-11, 
    5.428344e-11, 5.412596e-11, 5.413377e-11, 5.412954e-11, 5.413747e-11, 
    5.413184e-11, 5.415669e-11, 5.416413e-11, 5.419906e-11, 5.418487e-11, 
    5.42076e-11, 5.418723e-11, 5.419081e-11, 5.42081e-11, 5.418837e-11, 
    5.423212e-11, 5.420226e-11, 5.425778e-11, 5.422779e-11, 5.425964e-11, 
    5.425395e-11, 5.426343e-11, 5.427185e-11, 5.428254e-11, 5.430209e-11, 
    5.429759e-11, 5.4314e-11, 5.414547e-11, 5.415554e-11, 5.415476e-11, 
    5.416537e-11, 5.417319e-11, 5.419025e-11, 5.421745e-11, 5.420726e-11, 
    5.422608e-11, 5.422981e-11, 5.420129e-11, 5.421871e-11, 5.416236e-11, 
    5.417137e-11, 5.416608e-11, 5.41462e-11, 5.420947e-11, 5.417697e-11, 
    5.423702e-11, 5.421948e-11, 5.427064e-11, 5.424511e-11, 5.429508e-11, 
    5.431612e-11, 5.434032e-11, 5.436961e-11, 5.416115e-11, 5.41543e-11, 
    5.416666e-11, 5.418356e-11, 5.419951e-11, 5.422053e-11, 5.422274e-11, 
    5.422664e-11, 5.423688e-11, 5.424542e-11, 5.422778e-11, 5.424758e-11, 
    5.417325e-11, 5.421233e-11, 5.415161e-11, 5.416978e-11, 5.418261e-11, 
    5.417709e-11, 5.420612e-11, 5.421292e-11, 5.424047e-11, 5.42263e-11, 
    5.431084e-11, 5.427348e-11, 5.439223e-11, 5.43555e-11, 5.415188e-11, 
    5.416118e-11, 5.419335e-11, 5.417806e-11, 5.422199e-11, 5.423273e-11, 
    5.424155e-11, 5.425265e-11, 5.425392e-11, 5.426051e-11, 5.424971e-11, 
    5.426012e-11, 5.422058e-11, 5.423828e-11, 5.41898e-11, 5.420155e-11, 
    5.419618e-11, 5.419021e-11, 5.420861e-11, 5.422802e-11, 5.422861e-11, 
    5.42348e-11, 5.425193e-11, 5.422217e-11, 5.431534e-11, 5.425758e-11, 
    5.41713e-11, 5.418896e-11, 5.419168e-11, 5.418481e-11, 5.423165e-11, 
    5.421467e-11, 5.426037e-11, 5.424807e-11, 5.426826e-11, 5.425822e-11, 
    5.425673e-11, 5.424386e-11, 5.423579e-11, 5.421542e-11, 5.419887e-11, 
    5.418583e-11, 5.418887e-11, 5.420321e-11, 5.422925e-11, 5.425396e-11, 
    5.424853e-11, 5.426673e-11, 5.42188e-11, 5.423883e-11, 5.423104e-11, 
    5.425138e-11, 5.420695e-11, 5.424429e-11, 5.419733e-11, 5.420149e-11, 
    5.421434e-11, 5.424008e-11, 5.424601e-11, 5.425205e-11, 5.424836e-11, 
    5.422994e-11, 5.4227e-11, 5.421407e-11, 5.421041e-11, 5.42006e-11, 
    5.419239e-11, 5.419985e-11, 5.420764e-11, 5.423002e-11, 5.425006e-11, 
    5.427194e-11, 5.427736e-11, 5.430245e-11, 5.42818e-11, 5.431563e-11, 
    5.428652e-11, 5.434128e-11, 5.424669e-11, 5.428601e-11, 5.421498e-11, 
    5.422269e-11, 5.423644e-11, 5.42683e-11, 5.425129e-11, 5.427126e-11, 
    5.42269e-11, 5.420362e-11, 5.41978e-11, 5.418659e-11, 5.419806e-11, 
    5.419713e-11, 5.420808e-11, 5.420457e-11, 5.423077e-11, 5.421671e-11, 
    5.425665e-11, 5.427115e-11, 5.431222e-11, 5.434146e-11, 5.437397e-11, 
    5.43882e-11, 5.439255e-11, 5.439435e-11,
  2.415411e-14, 2.419185e-14, 2.418454e-14, 2.421494e-14, 2.419812e-14, 
    2.421799e-14, 2.416181e-14, 2.419331e-14, 2.417323e-14, 2.415758e-14, 
    2.427383e-14, 2.421631e-14, 2.433416e-14, 2.429734e-14, 2.439003e-14, 
    2.432835e-14, 2.44025e-14, 2.438837e-14, 2.443119e-14, 2.441893e-14, 
    2.447348e-14, 2.443686e-14, 2.450197e-14, 2.44648e-14, 2.447057e-14, 
    2.443563e-14, 2.4228e-14, 2.426663e-14, 2.422568e-14, 2.423119e-14, 
    2.422875e-14, 2.419843e-14, 2.418308e-14, 2.41513e-14, 2.415709e-14, 
    2.418047e-14, 2.423368e-14, 2.421569e-14, 2.426127e-14, 2.426024e-14, 
    2.431095e-14, 2.428808e-14, 2.437348e-14, 2.434922e-14, 2.441945e-14, 
    2.440176e-14, 2.441859e-14, 2.44135e-14, 2.441866e-14, 2.439273e-14, 
    2.440383e-14, 2.438106e-14, 2.429234e-14, 2.431836e-14, 2.424073e-14, 
    2.419393e-14, 2.416317e-14, 2.414126e-14, 2.414436e-14, 2.415024e-14, 
    2.418061e-14, 2.420928e-14, 2.423111e-14, 2.42457e-14, 2.426009e-14, 
    2.430338e-14, 2.432657e-14, 2.437832e-14, 2.436908e-14, 2.438482e-14, 
    2.44e-14, 2.442537e-14, 2.442121e-14, 2.443236e-14, 2.438448e-14, 
    2.441626e-14, 2.436379e-14, 2.437812e-14, 2.42636e-14, 2.422056e-14, 
    2.420193e-14, 2.418593e-14, 2.414673e-14, 2.417378e-14, 2.41631e-14, 
    2.418858e-14, 2.420473e-14, 2.419676e-14, 2.42461e-14, 2.422689e-14, 
    2.432794e-14, 2.428439e-14, 2.439823e-14, 2.437099e-14, 2.440478e-14, 
    2.438755e-14, 2.441704e-14, 2.43905e-14, 2.443654e-14, 2.444653e-14, 
    2.44397e-14, 2.446608e-14, 2.438902e-14, 2.441856e-14, 2.419652e-14, 
    2.419781e-14, 2.42039e-14, 2.417713e-14, 2.417552e-14, 2.415113e-14, 
    2.417287e-14, 2.41821e-14, 2.420569e-14, 2.421958e-14, 2.423281e-14, 
    2.426192e-14, 2.429439e-14, 2.433994e-14, 2.437275e-14, 2.439474e-14, 
    2.438128e-14, 2.439315e-14, 2.437986e-14, 2.437365e-14, 2.444276e-14, 
    2.440391e-14, 2.446229e-14, 2.445907e-14, 2.443261e-14, 2.445943e-14, 
    2.419873e-14, 2.419125e-14, 2.416518e-14, 2.418559e-14, 2.414848e-14, 
    2.416919e-14, 2.418108e-14, 2.422721e-14, 2.423744e-14, 2.424681e-14, 
    2.426541e-14, 2.428925e-14, 2.433106e-14, 2.436753e-14, 2.440091e-14, 
    2.439847e-14, 2.439932e-14, 2.440674e-14, 2.438831e-14, 2.440976e-14, 
    2.441333e-14, 2.440395e-14, 2.445864e-14, 2.444301e-14, 2.4459e-14, 
    2.444884e-14, 2.41937e-14, 2.420629e-14, 2.419948e-14, 2.421227e-14, 
    2.420323e-14, 2.424334e-14, 2.425537e-14, 2.431183e-14, 2.428875e-14, 
    2.43256e-14, 2.429253e-14, 2.429836e-14, 2.432663e-14, 2.429434e-14, 
    2.436544e-14, 2.431707e-14, 2.440703e-14, 2.435853e-14, 2.441006e-14, 
    2.440076e-14, 2.441619e-14, 2.442998e-14, 2.44474e-14, 2.447943e-14, 
    2.447203e-14, 2.44989e-14, 2.422512e-14, 2.424143e-14, 2.424007e-14, 
    2.42572e-14, 2.426986e-14, 2.42974e-14, 2.434151e-14, 2.432494e-14, 
    2.435545e-14, 2.436155e-14, 2.431525e-14, 2.43436e-14, 2.425241e-14, 
    2.426705e-14, 2.425839e-14, 2.422636e-14, 2.432865e-14, 2.427608e-14, 
    2.437327e-14, 2.434478e-14, 2.4428e-14, 2.438652e-14, 2.446794e-14, 
    2.450257e-14, 2.453786e-14, 2.457966e-14, 2.425042e-14, 2.423932e-14, 
    2.425926e-14, 2.428672e-14, 2.431243e-14, 2.434651e-14, 2.435003e-14, 
    2.43564e-14, 2.437298e-14, 2.438689e-14, 2.435834e-14, 2.439038e-14, 
    2.42703e-14, 2.433326e-14, 2.423506e-14, 2.426451e-14, 2.428514e-14, 
    2.427616e-14, 2.432307e-14, 2.43341e-14, 2.437894e-14, 2.43558e-14, 
    2.449396e-14, 2.443278e-14, 2.461175e-14, 2.455955e-14, 2.423543e-14, 
    2.425042e-14, 2.430251e-14, 2.427773e-14, 2.434882e-14, 2.43663e-14, 
    2.438058e-14, 2.439872e-14, 2.440073e-14, 2.441149e-14, 2.439385e-14, 
    2.441082e-14, 2.434658e-14, 2.437529e-14, 2.429664e-14, 2.431573e-14, 
    2.430697e-14, 2.429732e-14, 2.432712e-14, 2.435877e-14, 2.435957e-14, 
    2.43697e-14, 2.439804e-14, 2.434911e-14, 2.450163e-14, 2.440717e-14, 
    2.426676e-14, 2.429548e-14, 2.429974e-14, 2.428858e-14, 2.436454e-14, 
    2.433699e-14, 2.441124e-14, 2.439119e-14, 2.442408e-14, 2.440773e-14, 
    2.440531e-14, 2.438434e-14, 2.437126e-14, 2.433823e-14, 2.431141e-14, 
    2.429021e-14, 2.429515e-14, 2.431844e-14, 2.436073e-14, 2.440086e-14, 
    2.439205e-14, 2.442158e-14, 2.434366e-14, 2.437626e-14, 2.436361e-14, 
    2.439661e-14, 2.432448e-14, 2.438552e-14, 2.430884e-14, 2.431558e-14, 
    2.433645e-14, 2.437839e-14, 2.438785e-14, 2.439774e-14, 2.439166e-14, 
    2.436183e-14, 2.4357e-14, 2.433597e-14, 2.43301e-14, 2.431412e-14, 
    2.430084e-14, 2.431295e-14, 2.432564e-14, 2.436189e-14, 2.439452e-14, 
    2.443015e-14, 2.443893e-14, 2.448029e-14, 2.444645e-14, 2.450213e-14, 
    2.445453e-14, 2.453957e-14, 2.438924e-14, 2.445338e-14, 2.433744e-14, 
    2.434995e-14, 2.437245e-14, 2.442435e-14, 2.439645e-14, 2.442914e-14, 
    2.435682e-14, 2.431918e-14, 2.43096e-14, 2.429148e-14, 2.431002e-14, 
    2.430851e-14, 2.432625e-14, 2.432056e-14, 2.43631e-14, 2.434025e-14, 
    2.440522e-14, 2.442891e-14, 2.449604e-14, 2.453962e-14, 2.458569e-14, 
    2.460596e-14, 2.461215e-14, 2.461473e-14,
  3.238497e-18, 3.246673e-18, 3.245087e-18, 3.251938e-18, 3.248038e-18, 
    3.252645e-18, 3.240162e-18, 3.246989e-18, 3.242635e-18, 3.239245e-18, 
    3.26561e-18, 3.252254e-18, 3.279617e-18, 3.27105e-18, 3.29263e-18, 
    3.27827e-18, 3.295536e-18, 3.292237e-18, 3.302226e-18, 3.299363e-18, 
    3.31212e-18, 3.303548e-18, 3.318783e-18, 3.310083e-18, 3.311435e-18, 
    3.303262e-18, 3.254958e-18, 3.263938e-18, 3.254422e-18, 3.255702e-18, 
    3.255132e-18, 3.248111e-18, 3.244774e-18, 3.237887e-18, 3.23914e-18, 
    3.244206e-18, 3.256278e-18, 3.252105e-18, 3.262671e-18, 3.262433e-18, 
    3.274214e-18, 3.268897e-18, 3.288764e-18, 3.283113e-18, 3.299483e-18, 
    3.295357e-18, 3.299285e-18, 3.298096e-18, 3.2993e-18, 3.293252e-18, 
    3.295841e-18, 3.29053e-18, 3.269888e-18, 3.275937e-18, 3.257912e-18, 
    3.24713e-18, 3.240458e-18, 3.235715e-18, 3.236385e-18, 3.237659e-18, 
    3.244236e-18, 3.250621e-18, 3.255677e-18, 3.25906e-18, 3.262398e-18, 
    3.272466e-18, 3.27785e-18, 3.289898e-18, 3.287739e-18, 3.291411e-18, 
    3.294947e-18, 3.300867e-18, 3.299895e-18, 3.302501e-18, 3.291327e-18, 
    3.298743e-18, 3.286505e-18, 3.289847e-18, 3.263236e-18, 3.253234e-18, 
    3.248931e-18, 3.245389e-18, 3.236899e-18, 3.242756e-18, 3.240444e-18, 
    3.245961e-18, 3.249567e-18, 3.247732e-18, 3.259152e-18, 3.254702e-18, 
    3.27817e-18, 3.268045e-18, 3.294535e-18, 3.288183e-18, 3.296061e-18, 
    3.292043e-18, 3.298924e-18, 3.292731e-18, 3.303477e-18, 3.305812e-18, 
    3.304214e-18, 3.310378e-18, 3.292386e-18, 3.299278e-18, 3.247681e-18, 
    3.247967e-18, 3.249376e-18, 3.243483e-18, 3.243133e-18, 3.237849e-18, 
    3.242557e-18, 3.244557e-18, 3.249789e-18, 3.253007e-18, 3.256074e-18, 
    3.262826e-18, 3.270368e-18, 3.280958e-18, 3.288594e-18, 3.293717e-18, 
    3.29058e-18, 3.293349e-18, 3.29025e-18, 3.288802e-18, 3.304932e-18, 
    3.295861e-18, 3.309491e-18, 3.308738e-18, 3.30256e-18, 3.308823e-18, 
    3.248179e-18, 3.246539e-18, 3.240893e-18, 3.245311e-18, 3.237275e-18, 
    3.241762e-18, 3.24434e-18, 3.254779e-18, 3.257146e-18, 3.25932e-18, 
    3.263634e-18, 3.269169e-18, 3.278891e-18, 3.287381e-18, 3.295156e-18, 
    3.294587e-18, 3.294787e-18, 3.296518e-18, 3.292221e-18, 3.297225e-18, 
    3.298058e-18, 3.295869e-18, 3.308637e-18, 3.304986e-18, 3.308722e-18, 
    3.306347e-18, 3.247068e-18, 3.24993e-18, 3.248352e-18, 3.251316e-18, 
    3.249222e-18, 3.258521e-18, 3.261313e-18, 3.274424e-18, 3.269056e-18, 
    3.277622e-18, 3.269931e-18, 3.271288e-18, 3.277872e-18, 3.27035e-18, 
    3.286899e-18, 3.275646e-18, 3.296586e-18, 3.285294e-18, 3.297293e-18, 
    3.295122e-18, 3.298723e-18, 3.301943e-18, 3.306011e-18, 3.313505e-18, 
    3.311772e-18, 3.318058e-18, 3.25429e-18, 3.258075e-18, 3.257755e-18, 
    3.261729e-18, 3.264668e-18, 3.271061e-18, 3.281321e-18, 3.277464e-18, 
    3.284562e-18, 3.285984e-18, 3.275209e-18, 3.281809e-18, 3.26062e-18, 
    3.264023e-18, 3.262006e-18, 3.254581e-18, 3.278335e-18, 3.266118e-18, 
    3.288718e-18, 3.282081e-18, 3.301482e-18, 3.291809e-18, 3.310814e-18, 
    3.31893e-18, 3.326872e-18, 3.336192e-18, 3.260157e-18, 3.257582e-18, 
    3.262206e-18, 3.268588e-18, 3.274556e-18, 3.282483e-18, 3.283303e-18, 
    3.284786e-18, 3.288646e-18, 3.291889e-18, 3.285242e-18, 3.292703e-18, 
    3.264786e-18, 3.279403e-18, 3.256596e-18, 3.263432e-18, 3.268217e-18, 
    3.266131e-18, 3.277027e-18, 3.279595e-18, 3.29004e-18, 3.284645e-18, 
    3.316914e-18, 3.302605e-18, 3.343346e-18, 3.331709e-18, 3.256679e-18, 
    3.260154e-18, 3.272254e-18, 3.266494e-18, 3.28302e-18, 3.287092e-18, 
    3.290417e-18, 3.294649e-18, 3.295117e-18, 3.297628e-18, 3.293512e-18, 
    3.297471e-18, 3.2825e-18, 3.289185e-18, 3.270885e-18, 3.275323e-18, 
    3.273285e-18, 3.271041e-18, 3.27797e-18, 3.285343e-18, 3.285522e-18, 
    3.287886e-18, 3.294515e-18, 3.283088e-18, 3.318724e-18, 3.296644e-18, 
    3.263946e-18, 3.270625e-18, 3.271606e-18, 3.269012e-18, 3.286683e-18, 
    3.280269e-18, 3.29757e-18, 3.292891e-18, 3.300565e-18, 3.296748e-18, 
    3.296186e-18, 3.291295e-18, 3.288246e-18, 3.280559e-18, 3.27432e-18, 
    3.269391e-18, 3.270538e-18, 3.275955e-18, 3.2858e-18, 3.295149e-18, 
    3.293096e-18, 3.299982e-18, 3.281819e-18, 3.289414e-18, 3.28647e-18, 
    3.294155e-18, 3.277357e-18, 3.291593e-18, 3.273719e-18, 3.275287e-18, 
    3.280142e-18, 3.289915e-18, 3.292113e-18, 3.294422e-18, 3.293001e-18, 
    3.286054e-18, 3.284926e-18, 3.280029e-18, 3.278667e-18, 3.274947e-18, 
    3.27186e-18, 3.274675e-18, 3.27763e-18, 3.286066e-18, 3.293671e-18, 
    3.301986e-18, 3.304032e-18, 3.313718e-18, 3.305802e-18, 3.318843e-18, 
    3.307709e-18, 3.327269e-18, 3.292451e-18, 3.307425e-18, 3.28037e-18, 
    3.283281e-18, 3.28853e-18, 3.300638e-18, 3.294119e-18, 3.301754e-18, 
    3.284884e-18, 3.276132e-18, 3.273897e-18, 3.269687e-18, 3.273993e-18, 
    3.273644e-18, 3.277767e-18, 3.276443e-18, 3.286346e-18, 3.281025e-18, 
    3.296166e-18, 3.3017e-18, 3.317391e-18, 3.327269e-18, 3.337528e-18, 
    3.342052e-18, 3.343431e-18, 3.344007e-18,
  1.367581e-22, 1.372659e-22, 1.371673e-22, 1.375947e-22, 1.373507e-22, 
    1.376389e-22, 1.368614e-22, 1.372857e-22, 1.370149e-22, 1.368043e-22, 
    1.384511e-22, 1.376144e-22, 1.393391e-22, 1.387912e-22, 1.401877e-22, 
    1.392515e-22, 1.403773e-22, 1.401617e-22, 1.40814e-22, 1.406269e-22, 
    1.414619e-22, 1.409004e-22, 1.41898e-22, 1.413282e-22, 1.414168e-22, 
    1.408818e-22, 1.377834e-22, 1.383464e-22, 1.377499e-22, 1.378301e-22, 
    1.377943e-22, 1.373554e-22, 1.371482e-22, 1.3672e-22, 1.367978e-22, 
    1.371127e-22, 1.378662e-22, 1.376049e-22, 1.38266e-22, 1.382511e-22, 
    1.389896e-22, 1.386562e-22, 1.399351e-22, 1.395665e-22, 1.406348e-22, 
    1.403653e-22, 1.406219e-22, 1.405442e-22, 1.406229e-22, 1.40228e-22, 
    1.40397e-22, 1.400502e-22, 1.387184e-22, 1.390992e-22, 1.379683e-22, 
    1.372948e-22, 1.368798e-22, 1.365853e-22, 1.366269e-22, 1.36706e-22, 
    1.371145e-22, 1.375122e-22, 1.378283e-22, 1.3804e-22, 1.382489e-22, 
    1.388806e-22, 1.39224e-22, 1.400093e-22, 1.398681e-22, 1.401079e-22, 
    1.403386e-22, 1.407253e-22, 1.406617e-22, 1.408321e-22, 1.401022e-22, 
    1.405867e-22, 1.397876e-22, 1.400057e-22, 1.383025e-22, 1.376755e-22, 
    1.37407e-22, 1.371861e-22, 1.366588e-22, 1.370226e-22, 1.36879e-22, 
    1.372215e-22, 1.374463e-22, 1.373316e-22, 1.380458e-22, 1.377673e-22, 
    1.392448e-22, 1.386029e-22, 1.403116e-22, 1.398971e-22, 1.404113e-22, 
    1.401489e-22, 1.405984e-22, 1.401938e-22, 1.408959e-22, 1.410487e-22, 
    1.409442e-22, 1.413473e-22, 1.401713e-22, 1.406216e-22, 1.373284e-22, 
    1.373463e-22, 1.374342e-22, 1.370678e-22, 1.37046e-22, 1.367177e-22, 
    1.370101e-22, 1.371345e-22, 1.374601e-22, 1.376614e-22, 1.378532e-22, 
    1.382758e-22, 1.387486e-22, 1.394263e-22, 1.399239e-22, 1.402582e-22, 
    1.400534e-22, 1.402342e-22, 1.400319e-22, 1.399374e-22, 1.409912e-22, 
    1.403984e-22, 1.412893e-22, 1.4124e-22, 1.408361e-22, 1.412455e-22, 
    1.373595e-22, 1.372574e-22, 1.369068e-22, 1.371811e-22, 1.366821e-22, 
    1.369608e-22, 1.371211e-22, 1.377724e-22, 1.379202e-22, 1.380564e-22, 
    1.383264e-22, 1.386732e-22, 1.392916e-22, 1.398449e-22, 1.403521e-22, 
    1.40315e-22, 1.40328e-22, 1.404412e-22, 1.401606e-22, 1.404873e-22, 
    1.405419e-22, 1.403987e-22, 1.412333e-22, 1.409945e-22, 1.412389e-22, 
    1.410835e-22, 1.372903e-22, 1.374689e-22, 1.373703e-22, 1.375556e-22, 
    1.374248e-22, 1.380066e-22, 1.381814e-22, 1.39003e-22, 1.386662e-22, 
    1.39209e-22, 1.387209e-22, 1.388062e-22, 1.392258e-22, 1.387472e-22, 
    1.398137e-22, 1.390806e-22, 1.404456e-22, 1.397094e-22, 1.404917e-22, 
    1.403499e-22, 1.405851e-22, 1.407957e-22, 1.410616e-22, 1.415522e-22, 
    1.414386e-22, 1.418503e-22, 1.377415e-22, 1.379785e-22, 1.379583e-22, 
    1.382071e-22, 1.383912e-22, 1.387918e-22, 1.394498e-22, 1.391984e-22, 
    1.396609e-22, 1.397537e-22, 1.390519e-22, 1.394817e-22, 1.381378e-22, 
    1.383511e-22, 1.382245e-22, 1.377599e-22, 1.392555e-22, 1.384823e-22, 
    1.399321e-22, 1.394993e-22, 1.407656e-22, 1.40134e-22, 1.41376e-22, 
    1.41908e-22, 1.424196e-22, 1.430185e-22, 1.381087e-22, 1.379474e-22, 
    1.382369e-22, 1.386371e-22, 1.39011e-22, 1.395256e-22, 1.395788e-22, 
    1.396756e-22, 1.399273e-22, 1.401389e-22, 1.397056e-22, 1.40192e-22, 
    1.383993e-22, 1.393249e-22, 1.378859e-22, 1.383142e-22, 1.386137e-22, 
    1.384829e-22, 1.391699e-22, 1.393372e-22, 1.400185e-22, 1.396663e-22, 
    1.417759e-22, 1.408393e-22, 1.434779e-22, 1.427304e-22, 1.37891e-22, 
    1.381085e-22, 1.388668e-22, 1.385056e-22, 1.395604e-22, 1.39826e-22, 
    1.400428e-22, 1.403192e-22, 1.403496e-22, 1.405137e-22, 1.402448e-22, 
    1.405033e-22, 1.395266e-22, 1.399625e-22, 1.387806e-22, 1.390592e-22, 
    1.389312e-22, 1.387905e-22, 1.392313e-22, 1.397122e-22, 1.397235e-22, 
    1.398779e-22, 1.403117e-22, 1.395648e-22, 1.418953e-22, 1.404505e-22, 
    1.383459e-22, 1.387648e-22, 1.38826e-22, 1.386633e-22, 1.397993e-22, 
    1.393812e-22, 1.405099e-22, 1.402043e-22, 1.407055e-22, 1.404562e-22, 
    1.404195e-22, 1.401001e-22, 1.399013e-22, 1.394002e-22, 1.389963e-22, 
    1.38687e-22, 1.38759e-22, 1.391003e-22, 1.397419e-22, 1.403519e-22, 
    1.402179e-22, 1.406674e-22, 1.394821e-22, 1.399776e-22, 1.397856e-22, 
    1.402869e-22, 1.391915e-22, 1.401208e-22, 1.389584e-22, 1.390568e-22, 
    1.393729e-22, 1.400106e-22, 1.401535e-22, 1.403044e-22, 1.402115e-22, 
    1.397584e-22, 1.396848e-22, 1.393655e-22, 1.392769e-22, 1.390354e-22, 
    1.388418e-22, 1.390184e-22, 1.392094e-22, 1.397591e-22, 1.402554e-22, 
    1.407985e-22, 1.409321e-22, 1.415668e-22, 1.410486e-22, 1.419032e-22, 
    1.411742e-22, 1.424461e-22, 1.401763e-22, 1.411549e-22, 1.393877e-22, 
    1.395774e-22, 1.399201e-22, 1.407108e-22, 1.402845e-22, 1.407837e-22, 
    1.39682e-22, 1.39112e-22, 1.389696e-22, 1.387056e-22, 1.389756e-22, 
    1.389537e-22, 1.392181e-22, 1.391318e-22, 1.397773e-22, 1.394303e-22, 
    1.404183e-22, 1.4078e-22, 1.418067e-22, 1.424454e-22, 1.431037e-22, 
    1.433946e-22, 1.434832e-22, 1.435203e-22,
  1.875917e-27, 1.885557e-27, 1.883683e-27, 1.891701e-27, 1.887163e-27, 
    1.892523e-27, 1.877874e-27, 1.885936e-27, 1.880789e-27, 1.876791e-27, 
    1.907654e-27, 1.892068e-27, 1.924248e-27, 1.913985e-27, 1.940217e-27, 
    1.922605e-27, 1.943788e-27, 1.939721e-27, 1.952018e-27, 1.948489e-27, 
    1.964261e-27, 1.953648e-27, 1.972503e-27, 1.96173e-27, 1.963406e-27, 
    1.953297e-27, 1.895209e-27, 1.905703e-27, 1.894585e-27, 1.896079e-27, 
    1.895412e-27, 1.887252e-27, 1.883325e-27, 1.875192e-27, 1.876668e-27, 
    1.882648e-27, 1.896751e-27, 1.891889e-27, 1.904192e-27, 1.903914e-27, 
    1.917685e-27, 1.911465e-27, 1.935455e-27, 1.928517e-27, 1.948636e-27, 
    1.943557e-27, 1.948395e-27, 1.946929e-27, 1.948414e-27, 1.940971e-27, 
    1.944156e-27, 1.937622e-27, 1.912626e-27, 1.919738e-27, 1.89865e-27, 
    1.886112e-27, 1.878224e-27, 1.872653e-27, 1.873425e-27, 1.874927e-27, 
    1.882683e-27, 1.890164e-27, 1.896043e-27, 1.899983e-27, 1.903874e-27, 
    1.91566e-27, 1.922086e-27, 1.936853e-27, 1.934193e-27, 1.938711e-27, 
    1.943053e-27, 1.950346e-27, 1.949146e-27, 1.952362e-27, 1.938601e-27, 
    1.947732e-27, 1.932676e-27, 1.936783e-27, 1.904886e-27, 1.893202e-27, 
    1.888215e-27, 1.884041e-27, 1.874031e-27, 1.880936e-27, 1.87821e-27, 
    1.884711e-27, 1.888939e-27, 1.886802e-27, 1.900091e-27, 1.894909e-27, 
    1.922476e-27, 1.910475e-27, 1.942546e-27, 1.93474e-27, 1.944423e-27, 
    1.939479e-27, 1.947954e-27, 1.940326e-27, 1.953564e-27, 1.956451e-27, 
    1.954476e-27, 1.962087e-27, 1.939902e-27, 1.948391e-27, 1.886743e-27, 
    1.88708e-27, 1.888715e-27, 1.881795e-27, 1.88138e-27, 1.875149e-27, 
    1.880696e-27, 1.88306e-27, 1.889195e-27, 1.892939e-27, 1.896508e-27, 
    1.904376e-27, 1.913191e-27, 1.925885e-27, 1.935245e-27, 1.941538e-27, 
    1.93768e-27, 1.941086e-27, 1.937277e-27, 1.935496e-27, 1.955365e-27, 
    1.944183e-27, 1.960991e-27, 1.960059e-27, 1.952436e-27, 1.960165e-27, 
    1.887326e-27, 1.885393e-27, 1.878736e-27, 1.883944e-27, 1.874472e-27, 
    1.879763e-27, 1.882808e-27, 1.895007e-27, 1.897754e-27, 1.900289e-27, 
    1.905318e-27, 1.911782e-27, 1.923353e-27, 1.933759e-27, 1.943308e-27, 
    1.942608e-27, 1.942854e-27, 1.944987e-27, 1.9397e-27, 1.945857e-27, 
    1.946888e-27, 1.944187e-27, 1.959934e-27, 1.955425e-27, 1.96004e-27, 
    1.957103e-27, 1.886017e-27, 1.88936e-27, 1.887526e-27, 1.890973e-27, 
    1.88854e-27, 1.899366e-27, 1.902622e-27, 1.917941e-27, 1.911652e-27, 
    1.921801e-27, 1.912673e-27, 1.914264e-27, 1.922124e-27, 1.913162e-27, 
    1.933175e-27, 1.919393e-27, 1.945071e-27, 1.931215e-27, 1.945941e-27, 
    1.943267e-27, 1.9477e-27, 1.951673e-27, 1.956691e-27, 1.965963e-27, 
    1.963815e-27, 1.971599e-27, 1.894429e-27, 1.898842e-27, 1.898462e-27, 
    1.903095e-27, 1.906526e-27, 1.913994e-27, 1.926326e-27, 1.921599e-27, 
    1.930294e-27, 1.932041e-27, 1.918847e-27, 1.926927e-27, 1.901807e-27, 
    1.905782e-27, 1.903421e-27, 1.894772e-27, 1.922675e-27, 1.908228e-27, 
    1.935398e-27, 1.927255e-27, 1.951105e-27, 1.939203e-27, 1.96263e-27, 
    1.972697e-27, 1.982358e-27, 1.993937e-27, 1.901264e-27, 1.89826e-27, 
    1.903649e-27, 1.911113e-27, 1.918086e-27, 1.92775e-27, 1.92875e-27, 
    1.930571e-27, 1.935306e-27, 1.93929e-27, 1.931138e-27, 1.940291e-27, 
    1.906688e-27, 1.92398e-27, 1.897117e-27, 1.905095e-27, 1.910676e-27, 
    1.908235e-27, 1.921062e-27, 1.924206e-27, 1.937027e-27, 1.930395e-27, 
    1.9702e-27, 1.952501e-27, 2.002823e-27, 1.988366e-27, 1.897209e-27, 
    1.901258e-27, 1.915395e-27, 1.908658e-27, 1.928404e-27, 1.933401e-27, 
    1.937481e-27, 1.942691e-27, 1.943261e-27, 1.946356e-27, 1.941285e-27, 
    1.946159e-27, 1.92777e-27, 1.93597e-27, 1.913785e-27, 1.918984e-27, 
    1.916594e-27, 1.913969e-27, 1.922217e-27, 1.931264e-27, 1.931472e-27, 
    1.934379e-27, 1.942565e-27, 1.928486e-27, 1.972467e-27, 1.945179e-27, 
    1.90568e-27, 1.913497e-27, 1.914633e-27, 1.911597e-27, 1.932899e-27, 
    1.925035e-27, 1.946282e-27, 1.940523e-27, 1.949971e-27, 1.94527e-27, 
    1.944578e-27, 1.93856e-27, 1.934817e-27, 1.925392e-27, 1.917811e-27, 
    1.912039e-27, 1.913381e-27, 1.919758e-27, 1.931822e-27, 1.943306e-27, 
    1.940783e-27, 1.949252e-27, 1.926932e-27, 1.936256e-27, 1.932643e-27, 
    1.942079e-27, 1.92147e-27, 1.938964e-27, 1.917101e-27, 1.918938e-27, 
    1.924879e-27, 1.93688e-27, 1.939566e-27, 1.942411e-27, 1.940658e-27, 
    1.932132e-27, 1.930745e-27, 1.924738e-27, 1.923076e-27, 1.918539e-27, 
    1.914926e-27, 1.918224e-27, 1.921807e-27, 1.932141e-27, 1.941488e-27, 
    1.951728e-27, 1.954247e-27, 1.966247e-27, 1.956453e-27, 1.972617e-27, 
    1.958838e-27, 1.982884e-27, 1.940004e-27, 1.958463e-27, 1.925155e-27, 
    1.928723e-27, 1.935176e-27, 1.950077e-27, 1.942035e-27, 1.95145e-27, 
    1.930691e-27, 1.91998e-27, 1.91731e-27, 1.912387e-27, 1.917423e-27, 
    1.917014e-27, 1.921968e-27, 1.920347e-27, 1.932485e-27, 1.925957e-27, 
    1.944557e-27, 1.95138e-27, 1.970777e-27, 1.982864e-27, 1.995579e-27, 
    2.001207e-27, 2.002924e-27, 2.003641e-27,
  8.265279e-33, 8.322252e-33, 8.31116e-33, 8.35812e-33, 8.331727e-33, 
    8.3629e-33, 8.276825e-33, 8.324498e-33, 8.294049e-33, 8.270429e-33, 
    8.452032e-33, 8.360255e-33, 8.550994e-33, 8.489875e-33, 8.64565e-33, 
    8.54128e-33, 8.666852e-33, 8.642685e-33, 8.715767e-33, 8.694775e-33, 
    8.788752e-33, 8.725472e-33, 8.837945e-33, 8.773634e-33, 8.783642e-33, 
    8.723381e-33, 8.378517e-33, 8.440362e-33, 8.374892e-33, 8.383591e-33, 
    8.3797e-33, 8.332251e-33, 8.309062e-33, 8.260981e-33, 8.2697e-33, 
    8.305047e-33, 8.387508e-33, 8.359198e-33, 8.43126e-33, 8.429596e-33, 
    8.512047e-33, 8.474774e-33, 8.617371e-33, 8.576243e-33, 8.695651e-33, 
    8.665465e-33, 8.69422e-33, 8.685499e-33, 8.694334e-33, 8.650107e-33, 
    8.669026e-33, 8.630224e-33, 8.481732e-33, 8.524297e-33, 8.398559e-33, 
    8.325562e-33, 8.278899e-33, 8.246023e-33, 8.250557e-33, 8.25943e-33, 
    8.305253e-33, 8.349168e-33, 8.383367e-33, 8.406309e-33, 8.429355e-33, 
    8.499947e-33, 8.5382e-33, 8.625679e-33, 8.609882e-33, 8.636701e-33, 
    8.66247e-33, 8.705826e-33, 8.698684e-33, 8.717822e-33, 8.63603e-33, 
    8.690289e-33, 8.600884e-33, 8.625243e-33, 8.43548e-33, 8.366836e-33, 
    8.337869e-33, 8.313283e-33, 8.254135e-33, 8.294926e-33, 8.278817e-33, 
    8.317235e-33, 8.342046e-33, 8.329603e-33, 8.406938e-33, 8.376769e-33, 
    8.540507e-33, 8.468859e-33, 8.659461e-33, 8.613126e-33, 8.670609e-33, 
    8.641243e-33, 8.691601e-33, 8.646267e-33, 8.724972e-33, 8.742176e-33, 
    8.730412e-33, 8.775754e-33, 8.643755e-33, 8.6942e-33, 8.329255e-33, 
    8.331242e-33, 8.340741e-33, 8.300004e-33, 8.297548e-33, 8.260732e-33, 
    8.293501e-33, 8.307478e-33, 8.343527e-33, 8.365307e-33, 8.386076e-33, 
    8.432366e-33, 8.485127e-33, 8.560671e-33, 8.616121e-33, 8.653469e-33, 
    8.630563e-33, 8.650782e-33, 8.628175e-33, 8.617608e-33, 8.735712e-33, 
    8.66919e-33, 8.769219e-33, 8.763663e-33, 8.71827e-33, 8.76429e-33, 
    8.332672e-33, 8.321266e-33, 8.28192e-33, 8.312697e-33, 8.256736e-33, 
    8.287988e-33, 8.305996e-33, 8.377354e-33, 8.393328e-33, 8.408102e-33, 
    8.437992e-33, 8.476677e-33, 8.545682e-33, 8.607317e-33, 8.66398e-33, 
    8.659821e-33, 8.661283e-33, 8.673964e-33, 8.642556e-33, 8.679132e-33, 
    8.685265e-33, 8.669207e-33, 8.762918e-33, 8.736051e-33, 8.763545e-33, 
    8.746047e-33, 8.324959e-33, 8.344491e-33, 8.333832e-33, 8.353875e-33, 
    8.339733e-33, 8.402736e-33, 8.421903e-33, 8.513599e-33, 8.475903e-33, 
    8.536505e-33, 8.482008e-33, 8.491544e-33, 8.538444e-33, 8.484932e-33, 
    8.603868e-33, 8.522277e-33, 8.674457e-33, 8.592265e-33, 8.679628e-33, 
    8.663734e-33, 8.690084e-33, 8.713724e-33, 8.743591e-33, 8.798889e-33, 
    8.786064e-33, 8.832532e-33, 8.373977e-33, 8.399677e-33, 8.39745e-33, 
    8.424705e-33, 8.445225e-33, 8.489917e-33, 8.563272e-33, 8.535293e-33, 
    8.586768e-33, 8.597123e-33, 8.519e-33, 8.566838e-33, 8.417017e-33, 
    8.440795e-33, 8.426659e-33, 8.375979e-33, 8.541679e-33, 8.455423e-33, 
    8.617033e-33, 8.568773e-33, 8.710345e-33, 8.639624e-33, 8.779001e-33, 
    8.839122e-33, 8.896747e-33, 8.966275e-33, 8.413778e-33, 8.396274e-33, 
    8.428014e-33, 8.472685e-33, 8.514446e-33, 8.571702e-33, 8.577619e-33, 
    8.588412e-33, 8.616477e-33, 8.640122e-33, 8.59179e-33, 8.646063e-33, 
    8.446241e-33, 8.549391e-33, 8.38963e-33, 8.43669e-33, 8.470062e-33, 
    8.455446e-33, 8.53211e-33, 8.550716e-33, 8.626703e-33, 8.587365e-33, 
    8.824213e-33, 8.71867e-33, 9.020414e-33, 8.932812e-33, 8.390157e-33, 
    8.413735e-33, 8.498328e-33, 8.457976e-33, 8.575569e-33, 8.605192e-33, 
    8.629378e-33, 8.660325e-33, 8.663702e-33, 8.682098e-33, 8.651967e-33, 
    8.680922e-33, 8.571825e-33, 8.620423e-33, 8.488663e-33, 8.519832e-33, 
    8.505493e-33, 8.489762e-33, 8.538944e-33, 8.592538e-33, 8.59375e-33, 
    8.610994e-33, 8.659649e-33, 8.576058e-33, 8.837803e-33, 8.67517e-33, 
    8.440156e-33, 8.486967e-33, 8.49375e-33, 8.47556e-33, 8.602215e-33, 
    8.555629e-33, 8.681659e-33, 8.647439e-33, 8.703591e-33, 8.67564e-33, 
    8.671531e-33, 8.635787e-33, 8.613586e-33, 8.557748e-33, 8.512799e-33, 
    8.478203e-33, 8.48624e-33, 8.524414e-33, 8.595842e-33, 8.663979e-33, 
    8.649001e-33, 8.699312e-33, 8.566854e-33, 8.62213e-33, 8.600705e-33, 
    8.656686e-33, 8.534536e-33, 8.638258e-33, 8.508532e-33, 8.519548e-33, 
    8.554707e-33, 8.625849e-33, 8.641758e-33, 8.658661e-33, 8.64824e-33, 
    8.597674e-33, 8.589444e-33, 8.553866e-33, 8.544037e-33, 8.517154e-33, 
    8.495499e-33, 8.515266e-33, 8.536536e-33, 8.597721e-33, 8.65318e-33, 
    8.714052e-33, 8.729034e-33, 8.800623e-33, 8.742217e-33, 8.838704e-33, 
    8.756475e-33, 8.899968e-33, 8.644399e-33, 8.754198e-33, 8.556332e-33, 
    8.57746e-33, 8.61573e-33, 8.704254e-33, 8.656423e-33, 8.712416e-33, 
    8.589128e-33, 8.525737e-33, 8.509789e-33, 8.480291e-33, 8.510464e-33, 
    8.508009e-33, 8.537469e-33, 8.52788e-33, 8.599761e-33, 8.561082e-33, 
    8.671411e-33, 8.711988e-33, 8.827628e-33, 8.899804e-33, 8.976109e-33, 
    9.010455e-33, 9.021023e-33, 9.02544e-33,
  1.190679e-38, 1.202235e-38, 1.19998e-38, 1.20946e-38, 1.204157e-38, 
    1.21042e-38, 1.193015e-38, 1.202693e-38, 1.196507e-38, 1.191719e-38, 
    1.228438e-38, 1.209888e-38, 1.248528e-38, 1.236126e-38, 1.268109e-38, 
    1.246568e-38, 1.27253e-38, 1.267487e-38, 1.282758e-38, 1.278362e-38, 
    1.29811e-38, 1.284793e-38, 1.308503e-38, 1.29492e-38, 1.297031e-38, 
    1.284355e-38, 1.21356e-38, 1.226068e-38, 1.21283e-38, 1.214583e-38, 
    1.213798e-38, 1.204264e-38, 1.199558e-38, 1.189806e-38, 1.191571e-38, 
    1.19874e-38, 1.215372e-38, 1.209673e-38, 1.224209e-38, 1.223871e-38, 
    1.240646e-38, 1.233051e-38, 1.262218e-38, 1.253679e-38, 1.278546e-38, 
    1.272237e-38, 1.278247e-38, 1.276422e-38, 1.278271e-38, 1.269034e-38, 
    1.272982e-38, 1.264891e-38, 1.234468e-38, 1.243137e-38, 1.217598e-38, 
    1.202913e-38, 1.193436e-38, 1.186773e-38, 1.187698e-38, 1.189494e-38, 
    1.198782e-38, 1.207658e-38, 1.214535e-38, 1.219159e-38, 1.223822e-38, 
    1.238186e-38, 1.245944e-38, 1.263949e-38, 1.26066e-38, 1.266242e-38, 
    1.271612e-38, 1.280677e-38, 1.279181e-38, 1.283191e-38, 1.2661e-38, 
    1.277426e-38, 1.25879e-38, 1.263855e-38, 1.225078e-38, 1.211209e-38, 
    1.205395e-38, 1.200412e-38, 1.188422e-38, 1.196686e-38, 1.19342e-38, 
    1.201213e-38, 1.206228e-38, 1.203727e-38, 1.219285e-38, 1.213207e-38, 
    1.24641e-38, 1.231849e-38, 1.270985e-38, 1.261335e-38, 1.273311e-38, 
    1.267185e-38, 1.2777e-38, 1.268232e-38, 1.28469e-38, 1.288303e-38, 
    1.285832e-38, 1.295364e-38, 1.267709e-38, 1.278244e-38, 1.203657e-38, 
    1.20406e-38, 1.205966e-38, 1.197717e-38, 1.197218e-38, 1.189756e-38, 
    1.196396e-38, 1.199233e-38, 1.206524e-38, 1.210902e-38, 1.215082e-38, 
    1.224434e-38, 1.235161e-38, 1.250482e-38, 1.261958e-38, 1.269734e-38, 
    1.264961e-38, 1.269173e-38, 1.264464e-38, 1.262266e-38, 1.286946e-38, 
    1.273017e-38, 1.293988e-38, 1.292818e-38, 1.283285e-38, 1.29295e-38, 
    1.204347e-38, 1.202032e-38, 1.194048e-38, 1.200291e-38, 1.188947e-38, 
    1.195278e-38, 1.198934e-38, 1.213328e-38, 1.216542e-38, 1.219521e-38, 
    1.225575e-38, 1.233438e-38, 1.247453e-38, 1.260129e-38, 1.271927e-38, 
    1.271059e-38, 1.271364e-38, 1.274012e-38, 1.267459e-38, 1.275092e-38, 
    1.276375e-38, 1.273019e-38, 1.292661e-38, 1.287014e-38, 1.292793e-38, 
    1.289113e-38, 1.202783e-38, 1.206719e-38, 1.204579e-38, 1.208605e-38, 
    1.205765e-38, 1.218442e-38, 1.222316e-38, 1.240967e-38, 1.233281e-38, 
    1.245601e-38, 1.234523e-38, 1.236466e-38, 1.245997e-38, 1.235118e-38, 
    1.259416e-38, 1.242734e-38, 1.274115e-38, 1.25701e-38, 1.275195e-38, 
    1.271875e-38, 1.277381e-38, 1.282332e-38, 1.288598e-38, 1.300245e-38, 
    1.297538e-38, 1.307355e-38, 1.212645e-38, 1.217824e-38, 1.217372e-38, 
    1.22288e-38, 1.227044e-38, 1.236133e-38, 1.251007e-38, 1.245353e-38, 
    1.255861e-38, 1.258011e-38, 1.242064e-38, 1.251733e-38, 1.221323e-38, 
    1.226148e-38, 1.223277e-38, 1.21305e-38, 1.246646e-38, 1.229119e-38, 
    1.262148e-38, 1.252132e-38, 1.281624e-38, 1.266852e-38, 1.29605e-38, 
    1.308756e-38, 1.320936e-38, 1.335713e-38, 1.220666e-38, 1.217135e-38, 
    1.22355e-38, 1.232629e-38, 1.241136e-38, 1.252739e-38, 1.253964e-38, 
    1.256203e-38, 1.262031e-38, 1.266952e-38, 1.256907e-38, 1.26819e-38, 
    1.22726e-38, 1.248202e-38, 1.215798e-38, 1.225316e-38, 1.232094e-38, 
    1.229121e-38, 1.24471e-38, 1.248467e-38, 1.264161e-38, 1.255985e-38, 
    1.305601e-38, 1.283372e-38, 1.347445e-38, 1.328519e-38, 1.215903e-38, 
    1.220657e-38, 1.23785e-38, 1.229635e-38, 1.253539e-38, 1.259687e-38, 
    1.264714e-38, 1.271166e-38, 1.271869e-38, 1.275713e-38, 1.26942e-38, 
    1.275466e-38, 1.252765e-38, 1.262852e-38, 1.235877e-38, 1.242235e-38, 
    1.239308e-38, 1.236101e-38, 1.24609e-38, 1.257063e-38, 1.25731e-38, 
    1.260893e-38, 1.271039e-38, 1.25364e-38, 1.308486e-38, 1.274277e-38, 
    1.226014e-38, 1.235537e-38, 1.236915e-38, 1.233209e-38, 1.259068e-38, 
    1.249461e-38, 1.27562e-38, 1.268477e-38, 1.280208e-38, 1.274362e-38, 
    1.273504e-38, 1.266049e-38, 1.261431e-38, 1.24989e-38, 1.2408e-38, 
    1.233747e-38, 1.235384e-38, 1.24316e-38, 1.257747e-38, 1.271929e-38, 
    1.268805e-38, 1.279312e-38, 1.251734e-38, 1.263209e-38, 1.258757e-38, 
    1.270406e-38, 1.245201e-38, 1.266577e-38, 1.239927e-38, 1.242176e-38, 
    1.249275e-38, 1.263986e-38, 1.267293e-38, 1.270819e-38, 1.268644e-38, 
    1.258127e-38, 1.256418e-38, 1.249104e-38, 1.24712e-38, 1.241687e-38, 
    1.23727e-38, 1.241302e-38, 1.245606e-38, 1.258135e-38, 1.269676e-38, 
    1.282401e-38, 1.285541e-38, 1.300619e-38, 1.288317e-38, 1.308678e-38, 
    1.291325e-38, 1.321624e-38, 1.267851e-38, 1.290837e-38, 1.249602e-38, 
    1.253931e-38, 1.26188e-38, 1.280352e-38, 1.270351e-38, 1.282061e-38, 
    1.256352e-38, 1.243429e-38, 1.240184e-38, 1.234173e-38, 1.240322e-38, 
    1.239821e-38, 1.245792e-38, 1.243857e-38, 1.258559e-38, 1.250562e-38, 
    1.27348e-38, 1.28197e-38, 1.306318e-38, 1.321583e-38, 1.337831e-38, 
    1.345278e-38, 1.347575e-38, 1.348536e-38,
  5.605194e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 5.605194e-45, 7.006492e-45, 7.006492e-45, 5.605194e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 5.605194e-45, 5.605194e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 5.605194e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 5.605194e-45, 7.006492e-45, 5.605194e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 5.605194e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 5.605194e-45, 7.006492e-45, 5.605194e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 7.006492e-45, 
    7.006492e-45, 7.006492e-45, 7.006492e-45,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_CH4_UNSAT =
  9.109084e-06, 8.948252e-06, 8.979536e-06, 8.849694e-06, 8.921738e-06, 
    8.836692e-06, 9.076496e-06, 8.941861e-06, 9.027827e-06, 9.094617e-06, 
    8.597322e-06, 8.843898e-06, 8.340689e-06, 8.49833e-06, 8.101944e-06, 
    8.36523e-06, 8.048787e-06, 8.109554e-06, 7.926582e-06, 7.97903e-06, 
    7.744675e-06, 7.902368e-06, 7.623016e-06, 7.782357e-06, 7.757442e-06, 
    7.907565e-06, 8.794321e-06, 8.628045e-06, 8.804164e-06, 8.780469e-06, 
    8.791103e-06, 8.920249e-06, 8.985277e-06, 9.121371e-06, 9.096676e-06, 
    8.996714e-06, 8.769813e-06, 8.846886e-06, 8.652563e-06, 8.656954e-06, 
    8.440259e-06, 8.53801e-06, 8.173221e-06, 8.277013e-06, 7.976841e-06, 
    8.052401e-06, 7.98039e-06, 8.002231e-06, 7.980106e-06, 8.090904e-06, 
    8.043445e-06, 8.140896e-06, 8.519708e-06, 8.408499e-06, 8.739877e-06, 
    8.938697e-06, 9.070593e-06, 9.1641e-06, 9.150885e-06, 9.125688e-06, 
    8.99613e-06, 8.874201e-06, 8.7812e-06, 8.718951e-06, 8.657586e-06, 
    8.471638e-06, 8.373117e-06, 8.152218e-06, 8.192119e-06, 8.124522e-06, 
    8.059916e-06, 7.951361e-06, 7.969236e-06, 7.921385e-06, 8.12631e-06, 
    7.990154e-06, 8.214839e-06, 8.153426e-06, 8.640878e-06, 8.826099e-06, 
    8.904725e-06, 8.973522e-06, 9.140724e-06, 9.02528e-06, 9.070801e-06, 
    8.962481e-06, 8.893602e-06, 8.927675e-06, 8.717248e-06, 8.799097e-06, 
    8.367274e-06, 8.553462e-06, 8.067453e-06, 8.183931e-06, 8.039518e-06, 
    8.113231e-06, 7.986899e-06, 8.100603e-06, 7.903573e-06, 7.860624e-06, 
    7.889975e-06, 7.777194e-06, 8.106903e-06, 7.980389e-06, 8.928628e-06, 
    8.923072e-06, 8.897185e-06, 9.010938e-06, 9.017894e-06, 9.122048e-06, 
    9.029378e-06, 8.989893e-06, 8.889609e-06, 8.830251e-06, 8.7738e-06, 
    8.64959e-06, 8.510719e-06, 8.31627e-06, 8.176384e-06, 8.082523e-06, 
    8.140087e-06, 8.089267e-06, 8.146076e-06, 8.172694e-06, 7.876717e-06, 
    8.043001e-06, 7.793422e-06, 7.807247e-06, 7.920246e-06, 7.805689e-06, 
    8.91917e-06, 8.951141e-06, 9.062076e-06, 8.975268e-06, 9.133386e-06, 
    9.044901e-06, 8.993994e-06, 8.797383e-06, 8.754149e-06, 8.714041e-06, 
    8.634792e-06, 8.533008e-06, 8.354252e-06, 8.198506e-06, 8.056157e-06, 
    8.066592e-06, 8.062919e-06, 8.031095e-06, 8.109905e-06, 8.018152e-06, 
    8.002744e-06, 8.043023e-06, 7.809098e-06, 7.875976e-06, 7.807541e-06, 
    7.851091e-06, 8.94075e-06, 8.886946e-06, 8.916022e-06, 8.861339e-06, 
    8.899865e-06, 8.728459e-06, 8.677022e-06, 8.436056e-06, 8.535012e-06, 
    8.377491e-06, 8.519022e-06, 8.493954e-06, 8.372341e-06, 8.511379e-06, 
    8.207095e-06, 8.413465e-06, 8.029858e-06, 8.236236e-06, 8.016913e-06, 
    8.056772e-06, 7.990773e-06, 7.931629e-06, 7.857185e-06, 7.719694e-06, 
    7.751547e-06, 7.636475e-06, 8.806693e-06, 8.736823e-06, 8.74298e-06, 
    8.669826e-06, 8.615695e-06, 8.498293e-06, 8.309755e-06, 8.380689e-06, 
    8.250438e-06, 8.224271e-06, 8.422145e-06, 8.300688e-06, 8.690045e-06, 
    8.627218e-06, 8.664631e-06, 8.80118e-06, 8.364342e-06, 8.58872e-06, 
    8.174069e-06, 8.295865e-06, 7.940063e-06, 8.117137e-06, 7.769077e-06, 
    7.619957e-06, 7.479458e-06, 7.315024e-06, 8.698679e-06, 8.746172e-06, 
    8.661124e-06, 8.543354e-06, 8.43399e-06, 8.288439e-06, 8.273539e-06, 
    8.246247e-06, 8.175531e-06, 8.116039e-06, 8.237613e-06, 8.101121e-06, 
    8.612636e-06, 8.344848e-06, 8.764119e-06, 8.638013e-06, 8.550301e-06, 
    8.588789e-06, 8.388794e-06, 8.341609e-06, 8.149674e-06, 8.248933e-06, 
    7.656776e-06, 7.919127e-06, 7.189679e-06, 7.39399e-06, 8.76276e-06, 
    8.698844e-06, 8.47613e-06, 8.582148e-06, 8.278718e-06, 8.203911e-06, 
    8.143068e-06, 8.06524e-06, 8.056837e-06, 8.010697e-06, 8.086296e-06, 
    8.013686e-06, 8.288129e-06, 8.165564e-06, 8.501612e-06, 8.419904e-06, 
    8.4575e-06, 8.498724e-06, 8.371449e-06, 8.235699e-06, 8.232803e-06, 
    8.18924e-06, 8.066386e-06, 8.277488e-06, 7.622858e-06, 8.027556e-06, 
    8.629109e-06, 8.505825e-06, 8.488213e-06, 8.53599e-06, 8.211413e-06, 
    8.329119e-06, 8.011823e-06, 8.097662e-06, 7.956987e-06, 8.026911e-06, 
    8.037195e-06, 8.126935e-06, 8.18277e-06, 8.323723e-06, 8.438288e-06, 
    8.529063e-06, 8.507962e-06, 8.408228e-06, 8.227392e-06, 8.056073e-06, 
    8.093622e-06, 7.967684e-06, 8.300744e-06, 8.161195e-06, 8.215148e-06, 
    8.074418e-06, 8.382573e-06, 8.120191e-06, 8.449545e-06, 8.420706e-06, 
    8.331454e-06, 8.151719e-06, 8.111929e-06, 8.069416e-06, 8.095652e-06, 
    8.222799e-06, 8.24362e-06, 8.333625e-06, 8.358461e-06, 8.426986e-06, 
    8.483686e-06, 8.431881e-06, 8.377451e-06, 8.222748e-06, 8.083159e-06, 
    7.930786e-06, 7.89347e-06, 7.715113e-06, 7.860314e-06, 7.620599e-06, 
    7.824419e-06, 7.471376e-06, 8.104979e-06, 7.830421e-06, 8.327394e-06, 
    8.273953e-06, 8.17723e-06, 7.955105e-06, 8.075081e-06, 7.93476e-06, 
    8.244436e-06, 8.404782e-06, 8.446242e-06, 8.523545e-06, 8.444474e-06, 
    8.450907e-06, 8.3752e-06, 8.399535e-06, 8.217608e-06, 8.315365e-06, 
    8.037451e-06, 7.935871e-06, 7.648538e-06, 7.472038e-06, 7.292106e-06, 
    7.212576e-06, 7.18836e-06, 7.178234e-06,
  3.808703e-06, 3.674137e-06, 3.700163e-06, 3.592628e-06, 3.652142e-06, 
    3.581932e-06, 3.781286e-06, 3.668825e-06, 3.74048e-06, 3.796525e-06, 
    3.387302e-06, 3.58786e-06, 3.183708e-06, 3.308159e-06, 2.999129e-06, 
    3.202945e-06, 2.958684e-06, 3.004946e-06, 2.86662e-06, 2.905978e-06, 
    2.73195e-06, 2.84853e-06, 2.643523e-06, 2.759613e-06, 2.74131e-06, 
    2.852408e-06, 3.547165e-06, 3.41203e-06, 3.55523e-06, 3.535825e-06, 
    3.54453e-06, 3.650904e-06, 3.704937e-06, 3.819069e-06, 3.798258e-06, 
    3.714481e-06, 3.527112e-06, 3.590324e-06, 3.431845e-06, 3.435394e-06, 
    3.262084e-06, 3.339801e-06, 3.053744e-06, 3.134026e-06, 2.904331e-06, 
    2.961433e-06, 2.907001e-06, 2.923464e-06, 2.906787e-06, 2.990716e-06, 
    2.954637e-06, 3.028927e-06, 3.325189e-06, 3.236996e-06, 3.502687e-06, 
    3.66619e-06, 3.776325e-06, 3.855178e-06, 3.843995e-06, 3.822706e-06, 
    3.713993e-06, 3.612833e-06, 3.536429e-06, 3.485658e-06, 3.435905e-06, 
    3.286931e-06, 3.209142e-06, 3.037605e-06, 3.068296e-06, 3.016384e-06, 
    2.967138e-06, 2.885184e-06, 2.89861e-06, 2.86273e-06, 3.017757e-06, 
    2.914352e-06, 3.085831e-06, 3.038537e-06, 3.42238e-06, 3.573232e-06, 
    3.63804e-06, 3.695153e-06, 3.835404e-06, 3.738345e-06, 3.776499e-06, 
    3.68597e-06, 3.628855e-06, 3.657064e-06, 3.484274e-06, 3.55108e-06, 
    3.204554e-06, 3.352151e-06, 2.972865e-06, 3.061988e-06, 2.951663e-06, 
    3.007758e-06, 2.911901e-06, 2.998115e-06, 2.849427e-06, 2.817456e-06, 
    2.839287e-06, 2.755821e-06, 3.002923e-06, 2.906997e-06, 3.657854e-06, 
    3.653247e-06, 3.631818e-06, 3.726355e-06, 3.73217e-06, 3.819637e-06, 
    3.741777e-06, 3.708793e-06, 3.625558e-06, 3.576643e-06, 3.530375e-06, 
    3.42944e-06, 3.31802e-06, 3.164617e-06, 3.056178e-06, 2.984333e-06, 
    3.028309e-06, 2.989471e-06, 3.032899e-06, 3.053342e-06, 2.829415e-06, 
    2.954299e-06, 2.767762e-06, 2.777954e-06, 2.861878e-06, 2.776805e-06, 
    3.650014e-06, 3.676543e-06, 3.769177e-06, 3.696612e-06, 3.829207e-06, 
    3.754773e-06, 3.712209e-06, 3.549669e-06, 3.514329e-06, 3.481663e-06, 
    3.417496e-06, 3.335806e-06, 3.19434e-06, 3.073217e-06, 2.964285e-06, 
    2.972214e-06, 2.969421e-06, 2.945281e-06, 3.005216e-06, 2.935489e-06, 
    2.923848e-06, 2.954319e-06, 2.779321e-06, 2.828869e-06, 2.778171e-06, 
    2.810387e-06, 3.667913e-06, 3.623355e-06, 3.647407e-06, 3.602225e-06, 
    3.634031e-06, 3.493384e-06, 3.45162e-06, 3.258752e-06, 3.337404e-06, 
    3.212584e-06, 3.324644e-06, 3.304677e-06, 3.208525e-06, 3.318554e-06, 
    3.079839e-06, 3.240906e-06, 2.944345e-06, 3.102364e-06, 2.934553e-06, 
    2.964753e-06, 2.914823e-06, 2.870395e-06, 2.814907e-06, 2.713691e-06, 
    2.736993e-06, 2.653245e-06, 3.557305e-06, 3.500199e-06, 3.505221e-06, 
    3.445804e-06, 3.402106e-06, 3.308133e-06, 3.159533e-06, 3.215104e-06, 
    3.113387e-06, 3.09312e-06, 3.24777e-06, 3.152458e-06, 3.46218e-06, 
    3.41138e-06, 3.441598e-06, 3.552783e-06, 3.202253e-06, 3.38041e-06, 
    3.054397e-06, 3.148702e-06, 2.876712e-06, 3.010736e-06, 2.749855e-06, 
    2.64131e-06, 2.540882e-06, 2.425606e-06, 3.469187e-06, 3.507823e-06, 
    3.438766e-06, 3.344064e-06, 3.257127e-06, 3.142916e-06, 3.131325e-06, 
    3.110136e-06, 3.055525e-06, 3.009903e-06, 3.10344e-06, 2.998511e-06, 
    3.399622e-06, 3.18697e-06, 3.522464e-06, 3.420084e-06, 3.349622e-06, 
    3.380472e-06, 3.221482e-06, 3.184439e-06, 3.035654e-06, 3.11222e-06, 
    2.667922e-06, 2.861035e-06, 2.339425e-06, 2.480653e-06, 3.521358e-06, 
    3.469324e-06, 3.29051e-06, 3.375142e-06, 3.135353e-06, 3.077389e-06, 
    3.030594e-06, 2.971181e-06, 2.964801e-06, 2.929855e-06, 2.987207e-06, 
    2.932115e-06, 3.142674e-06, 3.047859e-06, 3.310776e-06, 3.245998e-06, 
    3.27574e-06, 3.308478e-06, 3.207843e-06, 3.101956e-06, 3.099722e-06, 
    3.066074e-06, 2.972026e-06, 3.134396e-06, 2.643387e-06, 2.942578e-06, 
    3.412915e-06, 3.314118e-06, 3.300114e-06, 3.338189e-06, 3.083181e-06, 
    3.174662e-06, 2.930706e-06, 2.995871e-06, 2.889408e-06, 2.942115e-06, 
    2.949901e-06, 3.018237e-06, 3.061095e-06, 3.170442e-06, 3.260525e-06, 
    3.332658e-06, 3.315832e-06, 3.236784e-06, 3.095528e-06, 2.964217e-06, 
    2.992784e-06, 2.897444e-06, 3.152507e-06, 3.044499e-06, 3.086063e-06, 
    2.978163e-06, 3.216583e-06, 3.013052e-06, 3.269438e-06, 3.246634e-06, 
    3.176489e-06, 3.037218e-06, 3.006762e-06, 2.974356e-06, 2.994339e-06, 
    3.091977e-06, 3.108098e-06, 3.17819e-06, 3.197644e-06, 3.251595e-06, 
    3.296519e-06, 3.25546e-06, 3.212554e-06, 3.091941e-06, 2.984813e-06, 
    2.869763e-06, 2.841894e-06, 2.710336e-06, 2.817217e-06, 2.641756e-06, 
    2.790605e-06, 2.53514e-06, 3.00144e-06, 2.79506e-06, 3.173316e-06, 
    3.131648e-06, 3.056822e-06, 2.887984e-06, 2.978667e-06, 2.872733e-06, 
    3.108731e-06, 3.234063e-06, 3.266822e-06, 3.328253e-06, 3.265422e-06, 
    3.270516e-06, 3.210791e-06, 3.229938e-06, 3.087968e-06, 3.163917e-06, 
    2.950094e-06, 2.873567e-06, 2.661966e-06, 2.53562e-06, 2.409748e-06, 
    2.355062e-06, 2.338528e-06, 2.331631e-06,
  1.765086e-06, 1.695146e-06, 1.708644e-06, 1.652961e-06, 1.683749e-06, 
    1.647436e-06, 1.750807e-06, 1.692393e-06, 1.729582e-06, 1.758742e-06, 
    1.547309e-06, 1.650498e-06, 1.443446e-06, 1.506827e-06, 1.350086e-06, 
    1.453221e-06, 1.329734e-06, 1.353017e-06, 1.283552e-06, 1.30327e-06, 
    1.216364e-06, 1.2745e-06, 1.172491e-06, 1.230129e-06, 1.221019e-06, 
    1.27644e-06, 1.629492e-06, 1.559986e-06, 1.633652e-06, 1.623644e-06, 
    1.628133e-06, 1.683108e-06, 1.711121e-06, 1.770489e-06, 1.759645e-06, 
    1.716076e-06, 1.619153e-06, 1.651771e-06, 1.570154e-06, 1.571976e-06, 
    1.483322e-06, 1.522996e-06, 1.377629e-06, 1.418241e-06, 1.302444e-06, 
    1.331116e-06, 1.303783e-06, 1.312043e-06, 1.303676e-06, 1.345849e-06, 
    1.3277e-06, 1.365105e-06, 1.515527e-06, 1.470543e-06, 1.606573e-06, 
    1.691027e-06, 1.748225e-06, 1.789325e-06, 1.783489e-06, 1.772385e-06, 
    1.715823e-06, 1.663406e-06, 1.623956e-06, 1.597809e-06, 1.572238e-06, 
    1.495991e-06, 1.456371e-06, 1.369483e-06, 1.38498e-06, 1.35878e-06, 
    1.333985e-06, 1.292847e-06, 1.299576e-06, 1.281604e-06, 1.359473e-06, 
    1.30747e-06, 1.393843e-06, 1.369953e-06, 1.565295e-06, 1.642943e-06, 
    1.676447e-06, 1.706045e-06, 1.779007e-06, 1.728472e-06, 1.748315e-06, 
    1.701282e-06, 1.671694e-06, 1.686299e-06, 1.597097e-06, 1.631511e-06, 
    1.454039e-06, 1.529313e-06, 1.336866e-06, 1.381793e-06, 1.326205e-06, 
    1.354433e-06, 1.306241e-06, 1.349576e-06, 1.274949e-06, 1.258972e-06, 
    1.269879e-06, 1.228241e-06, 1.351998e-06, 1.303781e-06, 1.686708e-06, 
    1.684322e-06, 1.673227e-06, 1.722243e-06, 1.725263e-06, 1.770785e-06, 
    1.730256e-06, 1.713124e-06, 1.669988e-06, 1.644705e-06, 1.620835e-06, 
    1.56892e-06, 1.511864e-06, 1.433754e-06, 1.378858e-06, 1.342637e-06, 
    1.364794e-06, 1.345223e-06, 1.367109e-06, 1.377427e-06, 1.264945e-06, 
    1.32753e-06, 1.234188e-06, 1.239266e-06, 1.281178e-06, 1.238693e-06, 
    1.682647e-06, 1.696394e-06, 1.744505e-06, 1.706802e-06, 1.775775e-06, 
    1.737012e-06, 1.714897e-06, 1.630783e-06, 1.612568e-06, 1.595754e-06, 
    1.562791e-06, 1.520954e-06, 1.448848e-06, 1.387466e-06, 1.33255e-06, 
    1.336538e-06, 1.335133e-06, 1.322999e-06, 1.353152e-06, 1.31808e-06, 
    1.312235e-06, 1.32754e-06, 1.239947e-06, 1.264673e-06, 1.239374e-06, 
    1.255443e-06, 1.69192e-06, 1.668848e-06, 1.681297e-06, 1.657921e-06, 
    1.674372e-06, 1.601784e-06, 1.580309e-06, 1.481624e-06, 1.521771e-06, 
    1.458122e-06, 1.515249e-06, 1.50505e-06, 1.456057e-06, 1.512137e-06, 
    1.390813e-06, 1.472533e-06, 1.322528e-06, 1.402206e-06, 1.31761e-06, 
    1.332786e-06, 1.307707e-06, 1.285441e-06, 1.257699e-06, 1.207289e-06, 
    1.218872e-06, 1.177305e-06, 1.634723e-06, 1.605291e-06, 1.607877e-06, 
    1.577322e-06, 1.554898e-06, 1.506814e-06, 1.431175e-06, 1.459404e-06, 
    1.407786e-06, 1.397529e-06, 1.47603e-06, 1.427586e-06, 1.585736e-06, 
    1.559653e-06, 1.575162e-06, 1.63239e-06, 1.452869e-06, 1.543779e-06, 
    1.377959e-06, 1.425681e-06, 1.288604e-06, 1.355934e-06, 1.225271e-06, 
    1.171396e-06, 1.121816e-06, 1.065229e-06, 1.589338e-06, 1.609217e-06, 
    1.573707e-06, 1.525176e-06, 1.480796e-06, 1.422747e-06, 1.416872e-06, 
    1.40614e-06, 1.378528e-06, 1.355514e-06, 1.402751e-06, 1.349775e-06, 
    1.553624e-06, 1.445103e-06, 1.616758e-06, 1.564118e-06, 1.528019e-06, 
    1.543811e-06, 1.462648e-06, 1.443818e-06, 1.368498e-06, 1.407196e-06, 
    1.184577e-06, 1.280756e-06, 1.023158e-06, 1.092207e-06, 1.616189e-06, 
    1.589408e-06, 1.497818e-06, 1.541081e-06, 1.418913e-06, 1.389575e-06, 
    1.365946e-06, 1.336018e-06, 1.33281e-06, 1.315251e-06, 1.344083e-06, 
    1.316385e-06, 1.422625e-06, 1.374658e-06, 1.508164e-06, 1.475127e-06, 
    1.490284e-06, 1.50699e-06, 1.455712e-06, 1.402e-06, 1.40087e-06, 
    1.383857e-06, 1.336442e-06, 1.418428e-06, 1.172423e-06, 1.321639e-06, 
    1.560441e-06, 1.509871e-06, 1.50272e-06, 1.522173e-06, 1.392503e-06, 
    1.438853e-06, 1.315678e-06, 1.348445e-06, 1.294964e-06, 1.321408e-06, 
    1.32532e-06, 1.359715e-06, 1.381341e-06, 1.436711e-06, 1.482528e-06, 
    1.519345e-06, 1.510747e-06, 1.470435e-06, 1.398747e-06, 1.332516e-06, 
    1.346891e-06, 1.298991e-06, 1.427611e-06, 1.372962e-06, 1.39396e-06, 
    1.339531e-06, 1.460156e-06, 1.3571e-06, 1.487071e-06, 1.475451e-06, 
    1.439781e-06, 1.369287e-06, 1.353932e-06, 1.337616e-06, 1.347674e-06, 
    1.396951e-06, 1.405109e-06, 1.440644e-06, 1.450527e-06, 1.477978e-06, 
    1.500885e-06, 1.479947e-06, 1.458107e-06, 1.396933e-06, 1.342878e-06, 
    1.285124e-06, 1.271182e-06, 1.205622e-06, 1.258852e-06, 1.171616e-06, 
    1.245572e-06, 1.118988e-06, 1.35125e-06, 1.247794e-06, 1.43817e-06, 
    1.417036e-06, 1.379183e-06, 1.29425e-06, 1.339785e-06, 1.286611e-06, 
    1.405429e-06, 1.46905e-06, 1.485737e-06, 1.517093e-06, 1.485024e-06, 
    1.48762e-06, 1.45721e-06, 1.466951e-06, 1.394924e-06, 1.433399e-06, 
    1.325416e-06, 1.287029e-06, 1.181626e-06, 1.119225e-06, 1.057473e-06, 
    1.030777e-06, 1.022722e-06, 1.019363e-06,
  4.452763e-07, 4.240201e-07, 4.281064e-07, 4.113005e-07, 4.205762e-07, 
    4.096401e-07, 4.409198e-07, 4.231876e-07, 4.3446e-07, 4.433398e-07, 
    3.797864e-07, 4.1056e-07, 3.492983e-07, 3.678441e-07, 3.223266e-07, 
    3.521461e-07, 3.165032e-07, 3.23167e-07, 3.033651e-07, 3.089617e-07, 
    2.844443e-07, 3.008028e-07, 2.722163e-07, 2.883019e-07, 2.857479e-07, 
    3.013515e-07, 4.042574e-07, 3.835413e-07, 4.055042e-07, 4.025062e-07, 
    4.038503e-07, 4.203826e-07, 4.288571e-07, 4.469269e-07, 4.436152e-07, 
    4.303595e-07, 4.011624e-07, 4.109427e-07, 3.865585e-07, 3.870997e-07, 
    3.609445e-07, 3.726051e-07, 3.302402e-07, 3.419755e-07, 3.087269e-07, 
    3.168981e-07, 3.091076e-07, 3.114579e-07, 3.09077e-07, 3.211128e-07, 
    3.159224e-07, 3.266374e-07, 3.704043e-07, 3.572042e-07, 3.974027e-07, 
    4.227747e-07, 4.40133e-07, 4.526912e-07, 4.509036e-07, 4.475065e-07, 
    4.302826e-07, 4.144426e-07, 4.025995e-07, 3.947877e-07, 3.871776e-07, 
    3.646602e-07, 3.530651e-07, 3.278958e-07, 3.323584e-07, 3.248208e-07, 
    3.17718e-07, 3.06001e-07, 3.079118e-07, 3.028136e-07, 3.250196e-07, 
    3.101563e-07, 3.349159e-07, 3.280312e-07, 3.851161e-07, 4.082911e-07, 
    4.183725e-07, 4.273189e-07, 4.495318e-07, 4.341229e-07, 4.401604e-07, 
    4.258766e-07, 4.169393e-07, 4.213462e-07, 3.945754e-07, 4.048624e-07, 
    3.523847e-07, 3.744683e-07, 3.185417e-07, 3.314397e-07, 3.154956e-07, 
    3.235734e-07, 3.098064e-07, 3.221805e-07, 3.009297e-07, 2.964164e-07, 
    2.99496e-07, 2.877723e-07, 3.228748e-07, 3.09107e-07, 4.214698e-07, 
    4.20749e-07, 4.174015e-07, 4.322308e-07, 4.331481e-07, 4.470176e-07, 
    4.34665e-07, 4.294641e-07, 4.164252e-07, 4.088199e-07, 4.016656e-07, 
    3.86192e-07, 3.693258e-07, 3.464789e-07, 3.305943e-07, 3.201929e-07, 
    3.265478e-07, 3.209334e-07, 3.272133e-07, 3.301819e-07, 2.981023e-07, 
    3.158738e-07, 2.894412e-07, 2.908679e-07, 3.026927e-07, 2.907069e-07, 
    4.202435e-07, 4.243976e-07, 4.389998e-07, 4.275482e-07, 4.485431e-07, 
    4.367194e-07, 4.300018e-07, 4.046442e-07, 3.991935e-07, 3.94175e-07, 
    3.843732e-07, 3.720029e-07, 3.508715e-07, 3.330755e-07, 3.17308e-07, 
    3.184479e-07, 3.180463e-07, 3.145805e-07, 3.23206e-07, 3.131778e-07, 
    3.115126e-07, 3.158767e-07, 2.910592e-07, 2.980253e-07, 2.908982e-07, 
    2.954213e-07, 4.230449e-07, 4.160817e-07, 4.19836e-07, 4.12792e-07, 
    4.177468e-07, 3.959733e-07, 3.895763e-07, 3.604471e-07, 3.722438e-07, 
    3.535758e-07, 3.703223e-07, 3.673214e-07, 3.529734e-07, 3.694062e-07, 
    3.340412e-07, 3.577862e-07, 3.144463e-07, 3.373325e-07, 3.130438e-07, 
    3.173752e-07, 3.102237e-07, 3.039005e-07, 2.960575e-07, 2.819067e-07, 
    2.851466e-07, 2.735531e-07, 4.058251e-07, 3.970202e-07, 3.977923e-07, 
    3.886881e-07, 3.820332e-07, 3.678403e-07, 3.457293e-07, 3.5395e-07, 
    3.389469e-07, 3.359807e-07, 3.588092e-07, 3.446868e-07, 3.911908e-07, 
    3.834427e-07, 3.880461e-07, 4.051257e-07, 3.520437e-07, 3.78742e-07, 
    3.303352e-07, 3.441338e-07, 3.047972e-07, 3.240037e-07, 2.869394e-07, 
    2.719121e-07, 2.582201e-07, 2.427576e-07, 3.922633e-07, 3.981924e-07, 
    3.876139e-07, 3.732478e-07, 3.602045e-07, 3.432823e-07, 3.415786e-07, 
    3.384705e-07, 3.304992e-07, 3.238835e-07, 3.3749e-07, 3.222376e-07, 
    3.816558e-07, 3.497808e-07, 4.004461e-07, 3.847669e-07, 3.740865e-07, 
    3.787515e-07, 3.548971e-07, 3.494066e-07, 3.276127e-07, 3.387759e-07, 
    2.755746e-07, 3.025732e-07, 2.313786e-07, 2.50107e-07, 4.002758e-07, 
    3.922843e-07, 3.651966e-07, 3.779443e-07, 3.421704e-07, 3.336839e-07, 
    3.26879e-07, 3.182994e-07, 3.173821e-07, 3.123716e-07, 3.20607e-07, 
    3.126949e-07, 3.432468e-07, 3.293848e-07, 3.682373e-07, 3.585449e-07, 
    3.629854e-07, 3.67892e-07, 3.528726e-07, 3.372729e-07, 3.369462e-07, 
    3.320347e-07, 3.184205e-07, 3.420298e-07, 2.721973e-07, 3.141927e-07, 
    3.836763e-07, 3.687393e-07, 3.666366e-07, 3.723622e-07, 3.34529e-07, 
    3.479616e-07, 3.124934e-07, 3.218566e-07, 3.066018e-07, 3.141267e-07, 
    3.152429e-07, 3.25089e-07, 3.313096e-07, 3.473385e-07, 3.607117e-07, 
    3.715288e-07, 3.689971e-07, 3.571726e-07, 3.363327e-07, 3.172982e-07, 
    3.214112e-07, 3.077457e-07, 3.446941e-07, 3.288966e-07, 3.349497e-07, 
    3.193041e-07, 3.541695e-07, 3.243384e-07, 3.620432e-07, 3.586398e-07, 
    3.482315e-07, 3.278396e-07, 3.234295e-07, 3.187561e-07, 3.216355e-07, 
    3.358136e-07, 3.38172e-07, 3.484828e-07, 3.513608e-07, 3.593793e-07, 
    3.660974e-07, 3.599559e-07, 3.535714e-07, 3.358084e-07, 3.20262e-07, 
    3.038108e-07, 2.998645e-07, 2.81441e-07, 2.963826e-07, 2.719731e-07, 
    2.92641e-07, 2.57443e-07, 3.226603e-07, 2.932665e-07, 3.477629e-07, 
    3.416261e-07, 3.306878e-07, 3.063991e-07, 3.193767e-07, 3.042322e-07, 
    3.382648e-07, 3.567676e-07, 3.616522e-07, 3.708655e-07, 3.614432e-07, 
    3.622043e-07, 3.533099e-07, 3.561541e-07, 3.35228e-07, 3.463757e-07, 
    3.152705e-07, 3.043506e-07, 2.747538e-07, 2.575082e-07, 2.406522e-07, 
    2.334317e-07, 2.31261e-07, 2.303572e-07,
  4.058013e-08, 3.816184e-08, 3.862414e-08, 3.673085e-08, 3.777318e-08, 
    3.654495e-08, 4.008179e-08, 3.806781e-08, 3.934541e-08, 4.035844e-08, 
    3.3239e-08, 3.664792e-08, 2.993632e-08, 3.193628e-08, 2.707956e-08, 
    3.024157e-08, 2.647108e-08, 2.716762e-08, 2.510943e-08, 2.568756e-08, 
    2.317632e-08, 2.484569e-08, 2.194502e-08, 2.356772e-08, 2.330843e-08, 
    2.490212e-08, 3.594376e-08, 3.365097e-08, 3.608281e-08, 3.574865e-08, 
    3.589838e-08, 3.775136e-08, 3.870921e-08, 4.07693e-08, 4.038995e-08, 
    3.887958e-08, 3.559909e-08, 3.669077e-08, 3.398281e-08, 3.40424e-08, 
    3.118892e-08, 3.245425e-08, 2.791124e-08, 2.915455e-08, 2.566325e-08, 
    2.651224e-08, 2.570266e-08, 2.594633e-08, 2.56995e-08, 2.695248e-08, 
    2.641054e-08, 2.753192e-08, 3.221459e-08, 3.078541e-08, 3.518139e-08, 
    3.802119e-08, 3.999193e-08, 4.143149e-08, 4.122587e-08, 4.083578e-08, 
    3.887085e-08, 3.70832e-08, 3.575904e-08, 3.489152e-08, 3.405098e-08, 
    3.159092e-08, 3.034022e-08, 2.766428e-08, 2.813477e-08, 2.734109e-08, 
    2.659776e-08, 2.538136e-08, 2.557888e-08, 2.505261e-08, 2.736196e-08, 
    2.581132e-08, 2.840519e-08, 2.767853e-08, 3.382408e-08, 3.639408e-08, 
    3.752496e-08, 3.853495e-08, 4.106824e-08, 3.930707e-08, 3.999507e-08, 
    3.837172e-08, 3.736372e-08, 3.786001e-08, 3.486801e-08, 3.601123e-08, 
    3.026718e-08, 3.265745e-08, 2.668373e-08, 2.803777e-08, 2.636609e-08, 
    2.721022e-08, 2.577506e-08, 2.706425e-08, 2.485874e-08, 2.439561e-08, 
    2.471143e-08, 2.35139e-08, 2.713699e-08, 2.57026e-08, 3.787394e-08, 
    3.779267e-08, 3.741571e-08, 3.909201e-08, 3.919624e-08, 4.07797e-08, 
    3.936873e-08, 3.877802e-08, 3.730592e-08, 3.64532e-08, 3.565508e-08, 
    3.394245e-08, 3.209729e-08, 2.963479e-08, 2.794857e-08, 2.685625e-08, 
    2.752251e-08, 2.693371e-08, 2.759247e-08, 2.790509e-08, 2.456839e-08, 
    2.640549e-08, 2.368358e-08, 2.382885e-08, 2.504016e-08, 2.381245e-08, 
    3.773569e-08, 3.820449e-08, 3.98626e-08, 3.856092e-08, 4.095472e-08, 
    3.960262e-08, 3.8839e-08, 3.598689e-08, 3.538021e-08, 3.482368e-08, 
    3.374238e-08, 3.238863e-08, 3.010487e-08, 2.821054e-08, 2.655498e-08, 
    2.667394e-08, 2.663202e-08, 2.627083e-08, 2.71717e-08, 2.612495e-08, 
    2.595201e-08, 2.640579e-08, 2.384835e-08, 2.456049e-08, 2.383194e-08, 
    2.429375e-08, 3.80517e-08, 3.726732e-08, 3.768977e-08, 3.689801e-08, 
    3.745455e-08, 3.502289e-08, 3.431543e-08, 3.113519e-08, 3.241487e-08, 
    3.039507e-08, 3.220567e-08, 3.187952e-08, 3.033038e-08, 3.210602e-08, 
    2.831264e-08, 3.084811e-08, 2.625686e-08, 2.866122e-08, 2.611102e-08, 
    2.656199e-08, 2.581831e-08, 2.516461e-08, 2.435887e-08, 2.291961e-08, 
    2.324747e-08, 2.207893e-08, 3.611864e-08, 3.513896e-08, 3.522463e-08, 
    3.421745e-08, 3.348537e-08, 3.193587e-08, 2.955474e-08, 3.043527e-08, 
    2.883255e-08, 2.851794e-08, 3.095841e-08, 2.944347e-08, 3.449368e-08, 
    3.364013e-08, 3.414668e-08, 3.604059e-08, 3.023058e-08, 3.312461e-08, 
    2.792125e-08, 2.938449e-08, 2.525709e-08, 2.725536e-08, 2.342931e-08, 
    2.191458e-08, 2.055365e-08, 1.903953e-08, 3.46122e-08, 3.526904e-08, 
    3.409905e-08, 3.252431e-08, 3.110899e-08, 2.929373e-08, 2.911231e-08, 
    2.878197e-08, 2.793855e-08, 2.724274e-08, 2.867793e-08, 2.707024e-08, 
    3.344396e-08, 2.998799e-08, 3.551943e-08, 3.378567e-08, 3.261579e-08, 
    3.312565e-08, 3.053708e-08, 2.994792e-08, 2.763449e-08, 2.881439e-08, 
    2.228175e-08, 2.502786e-08, 1.794123e-08, 1.975614e-08, 3.55005e-08, 
    3.461452e-08, 3.164904e-08, 3.30373e-08, 2.91753e-08, 2.827486e-08, 
    2.755732e-08, 2.665843e-08, 2.656271e-08, 2.604119e-08, 2.689956e-08, 
    2.607477e-08, 2.928994e-08, 2.782108e-08, 3.197898e-08, 3.092991e-08, 
    3.140958e-08, 3.194148e-08, 3.031955e-08, 2.86549e-08, 2.862026e-08, 
    2.810058e-08, 2.667107e-08, 2.916032e-08, 2.194312e-08, 2.623048e-08, 
    3.36658e-08, 3.203353e-08, 3.18052e-08, 3.242778e-08, 2.836424e-08, 
    2.979329e-08, 2.605384e-08, 2.703033e-08, 2.544343e-08, 2.622362e-08, 
    2.633978e-08, 2.736925e-08, 2.802405e-08, 2.972665e-08, 3.116377e-08, 
    3.2337e-08, 3.206155e-08, 3.0782e-08, 2.855523e-08, 2.655396e-08, 
    2.69837e-08, 2.55617e-08, 2.944425e-08, 2.776965e-08, 2.840877e-08, 
    2.676336e-08, 3.045886e-08, 2.729047e-08, 3.130766e-08, 3.094014e-08, 
    2.982215e-08, 2.765837e-08, 2.719513e-08, 2.670612e-08, 2.700718e-08, 
    2.850024e-08, 2.875029e-08, 2.984904e-08, 3.015733e-08, 3.101992e-08, 
    3.17467e-08, 3.108216e-08, 3.03946e-08, 2.849969e-08, 2.686348e-08, 
    2.515536e-08, 2.474926e-08, 2.287256e-08, 2.439215e-08, 2.192069e-08, 
    2.400965e-08, 2.047698e-08, 2.711452e-08, 2.407351e-08, 2.977202e-08, 
    2.911736e-08, 2.795844e-08, 2.542248e-08, 2.677094e-08, 2.519882e-08, 
    2.876013e-08, 3.073838e-08, 3.12654e-08, 3.226477e-08, 3.12428e-08, 
    3.132509e-08, 3.036651e-08, 3.067233e-08, 2.843822e-08, 2.962376e-08, 
    2.634265e-08, 2.521102e-08, 2.219935e-08, 2.048341e-08, 1.883528e-08, 
    1.813838e-08, 1.792996e-08, 1.784333e-08,
  1.171668e-09, 1.083894e-09, 1.100559e-09, 1.032659e-09, 1.069926e-09, 
    1.026042e-09, 1.15346e-09, 1.080511e-09, 1.126669e-09, 1.16356e-09, 
    9.099356e-10, 1.029706e-09, 7.97034e-10, 8.650212e-10, 7.02047e-10, 
    8.073335e-10, 6.821527e-10, 7.049359e-10, 6.38082e-10, 6.56717e-10, 
    5.76618e-10, 6.29619e-10, 5.381735e-10, 5.889554e-10, 5.80776e-10, 
    6.314279e-10, 1.004707e-09, 9.242397e-10, 1.009633e-09, 9.978038e-10, 
    1.003101e-09, 1.069143e-09, 1.103632e-09, 1.178595e-09, 1.164712e-09, 
    1.109791e-09, 9.925191e-10, 1.031231e-09, 9.35796e-10, 9.378748e-10, 
    8.394763e-10, 8.828209e-10, 7.294336e-10, 7.707858e-10, 6.55931e-10, 
    6.834946e-10, 6.572054e-10, 6.650947e-10, 6.571031e-10, 6.978821e-10, 
    6.801804e-10, 7.169152e-10, 8.745755e-10, 8.257526e-10, 9.777917e-10, 
    1.078835e-09, 1.150184e-09, 1.202914e-09, 1.195351e-09, 1.181032e-09, 
    1.109475e-09, 1.045224e-09, 9.981712e-10, 9.675991e-10, 9.381739e-10, 
    8.531963e-10, 8.106679e-10, 7.212781e-10, 7.368322e-10, 7.106348e-10, 
    6.862846e-10, 6.468331e-10, 6.532052e-10, 6.362566e-10, 7.11321e-10, 
    6.60721e-10, 7.458041e-10, 7.217482e-10, 9.302646e-10, 1.020679e-09, 
    1.061025e-09, 1.09734e-09, 1.18956e-09, 1.125277e-09, 1.150298e-09, 
    1.091453e-09, 1.055252e-09, 1.073043e-09, 9.667732e-10, 1.007096e-09, 
    8.081987e-10, 8.898252e-10, 6.890915e-10, 7.336196e-10, 6.787327e-10, 
    7.063347e-10, 6.595475e-10, 7.01545e-10, 6.300371e-10, 6.152323e-10, 
    6.253198e-10, 5.872556e-10, 7.039308e-10, 6.572035e-10, 1.073543e-09, 
    1.070625e-09, 1.057113e-09, 1.117481e-09, 1.121258e-09, 1.178976e-09, 
    1.127515e-09, 1.106118e-09, 1.053184e-09, 1.02278e-09, 9.944967e-10, 
    9.34389e-10, 8.705459e-10, 7.868877e-10, 7.306682e-10, 6.947318e-10, 
    7.166051e-10, 6.972671e-10, 7.189105e-10, 7.292301e-10, 6.207467e-10, 
    6.800157e-10, 5.926182e-10, 5.972171e-10, 6.358569e-10, 5.966976e-10, 
    1.06858e-09, 1.085429e-09, 1.145471e-09, 1.098277e-09, 1.185394e-09, 
    1.136011e-09, 1.108323e-09, 1.006235e-09, 9.847958e-10, 9.65217e-10, 
    9.274201e-10, 8.805619e-10, 8.027174e-10, 7.393437e-10, 6.848888e-10, 
    6.887718e-10, 6.874027e-10, 6.756325e-10, 7.050701e-10, 6.70891e-10, 
    6.652789e-10, 6.800255e-10, 5.978351e-10, 6.204945e-10, 5.973152e-10, 
    6.119863e-10, 1.079931e-09, 1.051804e-09, 1.066933e-09, 1.038616e-09, 
    1.058503e-09, 9.722153e-10, 9.474106e-10, 8.37646e-10, 8.814652e-10, 
    8.125233e-10, 8.742689e-10, 8.630756e-10, 8.103351e-10, 8.708458e-10, 
    7.427309e-10, 8.278822e-10, 6.751782e-10, 7.543199e-10, 6.704386e-10, 
    6.851174e-10, 6.609473e-10, 6.398558e-10, 6.140608e-10, 5.685566e-10, 
    5.788566e-10, 5.42327e-10, 1.010903e-09, 9.762982e-10, 9.793139e-10, 
    9.439863e-10, 9.184842e-10, 8.65007e-10, 7.841989e-10, 8.138836e-10, 
    7.600295e-10, 7.495516e-10, 8.316305e-10, 7.804646e-10, 9.536475e-10, 
    9.238625e-10, 9.415142e-10, 1.008137e-09, 8.069622e-10, 9.059724e-10, 
    7.297647e-10, 7.784867e-10, 6.428306e-10, 7.078172e-10, 5.845864e-10, 
    5.372302e-10, 4.954228e-10, 4.497741e-10, 9.577993e-10, 9.808782e-10, 
    9.398516e-10, 8.852347e-10, 8.367541e-10, 7.754451e-10, 7.693731e-10, 
    7.583429e-10, 7.303366e-10, 7.074028e-10, 7.548762e-10, 7.017412e-10, 
    9.170462e-10, 7.987753e-10, 9.897069e-10, 9.28927e-10, 8.883881e-10, 
    9.060082e-10, 8.173311e-10, 7.974247e-10, 7.202957e-10, 7.594241e-10, 
    5.486309e-10, 6.354619e-10, 4.172595e-10, 4.712625e-10, 9.890385e-10, 
    9.578807e-10, 8.551839e-10, 9.029497e-10, 7.7148e-10, 7.41477e-10, 
    7.177521e-10, 6.882652e-10, 6.85141e-10, 6.681715e-10, 6.961493e-10, 
    6.692616e-10, 7.753184e-10, 7.26454e-10, 8.664856e-10, 8.306616e-10, 
    8.470013e-10, 8.651996e-10, 8.09969e-10, 7.541094e-10, 7.529561e-10, 
    7.356997e-10, 6.886782e-10, 7.709791e-10, 5.381144e-10, 6.743203e-10, 
    9.247553e-10, 8.683572e-10, 8.605292e-10, 8.819094e-10, 7.44444e-10, 
    7.922175e-10, 6.685821e-10, 7.004329e-10, 6.488341e-10, 6.740972e-10, 
    6.778761e-10, 7.115608e-10, 7.331654e-10, 7.899759e-10, 8.386195e-10, 
    8.787849e-10, 8.693187e-10, 8.25637e-10, 7.50792e-10, 6.848555e-10, 
    6.989049e-10, 6.526504e-10, 7.804907e-10, 7.247553e-10, 7.459229e-10, 
    6.916936e-10, 8.146822e-10, 7.08971e-10, 8.435239e-10, 8.310094e-10, 
    7.931888e-10, 7.210832e-10, 7.058393e-10, 6.898229e-10, 6.996742e-10, 
    7.489631e-10, 7.57287e-10, 7.940941e-10, 8.044881e-10, 8.337225e-10, 
    8.58526e-10, 8.358404e-10, 8.125073e-10, 7.489447e-10, 6.949683e-10, 
    6.395584e-10, 6.265308e-10, 5.670818e-10, 6.151219e-10, 5.374193e-10, 
    6.029519e-10, 4.930888e-10, 7.031936e-10, 6.0498e-10, 7.915021e-10, 
    7.695419e-10, 7.309947e-10, 6.481586e-10, 6.919414e-10, 6.409557e-10, 
    7.57615e-10, 8.241564e-10, 8.420827e-10, 8.763007e-10, 8.413125e-10, 
    8.441183e-10, 8.115572e-10, 8.219153e-10, 7.469015e-10, 7.865174e-10, 
    6.779695e-10, 6.413484e-10, 5.46068e-10, 4.932844e-10, 4.436887e-10, 
    4.230579e-10, 4.169285e-10, 4.143864e-10,
  9.441462e-12, 8.513e-12, 8.687612e-12, 7.981235e-12, 8.367261e-12, 
    7.913131e-12, 9.247104e-12, 8.477653e-12, 8.962772e-12, 9.354805e-12, 
    6.740193e-12, 7.950826e-12, 5.642604e-12, 6.298231e-12, 4.755479e-12, 
    5.740857e-12, 4.574221e-12, 4.781935e-12, 4.178641e-12, 4.34489e-12, 
    3.64136e-12, 4.103644e-12, 3.314397e-12, 3.747804e-12, 3.677154e-12, 
    4.119646e-12, 7.694435e-12, 6.882366e-12, 7.744806e-12, 7.62397e-12, 
    7.678023e-12, 8.359109e-12, 8.719895e-12, 9.51565e-12, 9.367105e-12, 
    8.784683e-12, 7.570124e-12, 7.966532e-12, 6.997717e-12, 7.018513e-12, 
    6.04996e-12, 6.472562e-12, 5.007637e-12, 5.393987e-12, 4.337848e-12, 
    4.586395e-12, 4.349268e-12, 4.420121e-12, 4.348351e-12, 4.717396e-12, 
    4.55634e-12, 4.892001e-12, 6.391671e-12, 5.917531e-12, 7.420529e-12, 
    8.460148e-12, 9.212223e-12, 9.7771e-12, 9.695625e-12, 9.541773e-12, 
    8.78136e-12, 8.110937e-12, 7.627715e-12, 7.317394e-12, 7.021506e-12, 
    6.183022e-12, 5.772749e-12, 4.932232e-12, 5.076273e-12, 4.834225e-12, 
    4.611732e-12, 4.256525e-12, 4.313445e-12, 4.162438e-12, 4.840529e-12, 
    4.380809e-12, 5.159791e-12, 4.93657e-12, 6.942451e-12, 7.858023e-12, 
    8.274695e-12, 8.653818e-12, 9.633341e-12, 8.948062e-12, 9.213441e-12, 
    8.592099e-12, 8.214778e-12, 8.399735e-12, 7.309052e-12, 7.718858e-12, 
    5.749128e-12, 6.541459e-12, 4.637254e-12, 5.046443e-12, 4.543226e-12, 
    4.794757e-12, 4.370274e-12, 4.750885e-12, 4.107341e-12, 3.976885e-12, 
    4.065667e-12, 3.733096e-12, 4.772726e-12, 4.349251e-12, 8.404949e-12, 
    8.374545e-12, 8.234076e-12, 8.865727e-12, 8.905592e-12, 9.519731e-12, 
    8.971724e-12, 8.746038e-12, 8.193339e-12, 7.879601e-12, 7.590263e-12, 
    6.983649e-12, 6.352223e-12, 5.546195e-12, 5.019075e-12, 4.68864e-12, 
    4.889145e-12, 4.71178e-12, 4.91039e-12, 5.005752e-12, 4.025361e-12, 
    4.554847e-12, 3.779544e-12, 3.819485e-12, 4.158892e-12, 3.814968e-12, 
    8.353252e-12, 8.52905e-12, 9.162111e-12, 8.663651e-12, 9.588583e-12, 
    9.061695e-12, 8.769234e-12, 7.710045e-12, 7.49159e-12, 7.293339e-12, 
    6.914067e-12, 6.450378e-12, 5.696773e-12, 5.09962e-12, 4.599051e-12, 
    4.634346e-12, 4.621894e-12, 4.515173e-12, 4.783164e-12, 4.472346e-12, 
    4.421778e-12, 4.554937e-12, 3.824859e-12, 4.023141e-12, 3.820338e-12, 
    3.948415e-12, 8.471597e-12, 8.179034e-12, 8.336109e-12, 8.042666e-12, 
    8.248507e-12, 7.364064e-12, 7.114089e-12, 6.032261e-12, 6.459246e-12, 
    5.790513e-12, 6.388667e-12, 6.279241e-12, 5.769565e-12, 6.355157e-12, 
    5.131148e-12, 5.938037e-12, 4.511065e-12, 5.239355e-12, 4.468264e-12, 
    4.601129e-12, 4.38284e-12, 4.1944e-12, 3.966605e-12, 3.572202e-12, 
    3.66062e-12, 3.34937e-12, 7.757803e-12, 7.405397e-12, 7.435959e-12, 
    7.079734e-12, 6.825077e-12, 6.298091e-12, 5.52071e-12, 5.803544e-12, 
    5.292856e-12, 5.19477e-12, 5.974169e-12, 5.485362e-12, 7.176757e-12, 
    6.878608e-12, 7.054956e-12, 7.729498e-12, 5.737308e-12, 6.70092e-12, 
    5.010704e-12, 5.46666e-12, 4.220862e-12, 4.808355e-12, 3.710027e-12, 
    3.306468e-12, 2.95961e-12, 2.591697e-12, 7.218544e-12, 7.451824e-12, 
    7.038302e-12, 6.496287e-12, 6.023639e-12, 5.43793e-12, 5.380679e-12, 
    5.27704e-12, 5.016003e-12, 4.804553e-12, 5.244562e-12, 4.75268e-12, 
    6.810783e-12, 5.659188e-12, 7.541507e-12, 6.929101e-12, 6.52731e-12, 
    6.701274e-12, 5.8366e-12, 5.646324e-12, 4.923166e-12, 5.287178e-12, 
    3.402613e-12, 4.155389e-12, 2.337007e-12, 2.763428e-12, 7.534709e-12, 
    7.219363e-12, 6.202353e-12, 6.671003e-12, 5.400529e-12, 5.119472e-12, 
    4.899712e-12, 4.629738e-12, 4.601342e-12, 4.447824e-12, 4.701574e-12, 
    4.45765e-12, 5.436734e-12, 4.980056e-12, 6.312532e-12, 5.964825e-12, 
    6.122858e-12, 6.299972e-12, 5.76606e-12, 5.237385e-12, 5.226593e-12, 
    5.065752e-12, 4.633495e-12, 5.395807e-12, 3.313901e-12, 4.503312e-12, 
    6.887502e-12, 6.330821e-12, 6.254408e-12, 6.463609e-12, 5.14711e-12, 
    5.59679e-12, 4.451525e-12, 4.740712e-12, 4.27438e-12, 4.501295e-12, 
    4.535471e-12, 4.842732e-12, 5.042229e-12, 5.575498e-12, 6.041672e-12, 
    6.432938e-12, 6.340221e-12, 5.916419e-12, 5.20636e-12, 4.598749e-12, 
    4.726742e-12, 4.308482e-12, 5.485609e-12, 4.964349e-12, 5.160899e-12, 
    4.660944e-12, 5.811197e-12, 4.818945e-12, 6.089146e-12, 5.968178e-12, 
    5.606023e-12, 4.930433e-12, 4.790215e-12, 4.64391e-12, 4.733774e-12, 
    5.189273e-12, 5.267142e-12, 5.614629e-12, 5.713674e-12, 5.994357e-12, 
    6.234888e-12, 6.01481e-12, 5.79036e-12, 5.189102e-12, 4.690797e-12, 
    4.191757e-12, 4.076356e-12, 3.559582e-12, 3.975916e-12, 3.308057e-12, 
    3.869429e-12, 2.940518e-12, 4.765975e-12, 3.887127e-12, 5.589992e-12, 
    5.382269e-12, 5.022101e-12, 4.268351e-12, 4.663202e-12, 4.20418e-12, 
    5.270216e-12, 5.902172e-12, 6.075187e-12, 6.408577e-12, 6.06773e-12, 
    6.094905e-12, 5.78126e-12, 5.880623e-12, 5.170028e-12, 5.542683e-12, 
    4.536317e-12, 4.207672e-12, 3.380943e-12, 2.942117e-12, 2.543549e-12, 
    2.381957e-12, 2.334447e-12, 2.314811e-12,
  1.192371e-14, 9.864111e-15, 1.024209e-14, 8.741158e-15, 9.55208e-15, 
    8.600494e-15, 1.148261e-14, 9.788142e-15, 1.084667e-14, 1.172641e-14, 
    6.29845e-15, 8.67826e-15, 4.373449e-15, 5.494627e-15, 3.006864e-15, 
    4.53577e-15, 2.751131e-15, 3.044892e-15, 2.223329e-15, 2.439943e-15, 
    1.578357e-15, 2.128161e-15, 1.230292e-15, 1.699161e-15, 1.61858e-15, 
    2.148332e-15, 8.153779e-15, 6.564767e-15, 8.255987e-15, 8.011492e-15, 
    8.120568e-15, 9.53472e-15, 1.031246e-14, 1.209342e-14, 1.175435e-14, 
    1.045414e-14, 7.903312e-15, 8.710728e-15, 6.783517e-15, 6.823207e-15, 
    5.059703e-15, 5.807258e-15, 3.376392e-15, 3.972129e-15, 2.430612e-15, 
    2.768041e-15, 2.44575e-15, 2.540469e-15, 2.444533e-15, 2.952435e-15, 
    2.726364e-15, 3.204984e-15, 5.661465e-15, 4.832804e-15, 7.605282e-15, 
    9.750592e-15, 1.1404e-14, 1.269732e-14, 1.250817e-14, 1.215335e-14, 
    1.044686e-14, 9.011063e-15, 8.019033e-15, 7.401998e-15, 6.828926e-15, 
    5.291278e-15, 4.588902e-15, 3.264248e-15, 3.479663e-15, 3.120571e-15, 
    2.803358e-15, 2.323848e-15, 2.398383e-15, 2.202632e-15, 3.129742e-15, 
    2.487747e-15, 3.606841e-15, 3.270662e-15, 6.678419e-15, 8.487207e-15, 
    9.355553e-15, 1.016859e-14, 1.236415e-14, 1.081408e-14, 1.140674e-14, 
    1.003478e-14, 9.229029e-15, 9.621331e-15, 7.385633e-15, 8.203282e-15, 
    4.549529e-15, 5.932421e-15, 2.839102e-15, 3.434642e-15, 2.708254e-15, 
    3.063386e-15, 2.47369e-15, 3.000279e-15, 2.132815e-15, 1.971009e-15, 
    2.080587e-15, 1.682256e-15, 3.031636e-15, 2.445727e-15, 9.632467e-15, 
    9.5676e-15, 9.269718e-15, 1.063221e-14, 1.072015e-14, 1.210278e-14, 
    1.086652e-14, 1.036955e-14, 9.183892e-15, 8.531506e-15, 7.943715e-15, 
    6.756712e-15, 5.590825e-15, 4.216205e-15, 3.393524e-15, 2.911579e-15, 
    3.20079e-15, 2.944439e-15, 3.232023e-15, 3.373573e-15, 2.030554e-15, 
    2.724301e-15, 1.735869e-15, 1.782505e-15, 2.198113e-15, 1.777207e-15, 
    9.522255e-15, 9.898665e-15, 1.129134e-14, 1.018996e-14, 1.226097e-14, 
    1.106665e-14, 1.04203e-14, 8.185411e-15, 7.746385e-15, 7.354843e-15, 
    6.624644e-15, 5.76715e-15, 4.462683e-15, 3.515049e-15, 2.785662e-15, 
    2.835021e-15, 2.81757e-15, 2.669665e-15, 3.046664e-15, 2.611155e-15, 
    2.542702e-15, 2.724424e-15, 1.788818e-15, 2.027811e-15, 1.783506e-15, 
    1.936362e-15, 9.775141e-15, 9.153814e-15, 9.485795e-15, 8.868668e-15, 
    9.300185e-15, 7.493766e-15, 7.006604e-15, 5.029171e-15, 5.783173e-15, 
    4.618589e-15, 5.656076e-15, 5.460928e-15, 4.583588e-15, 5.596067e-15, 
    3.563039e-15, 4.867703e-15, 2.664031e-15, 3.729522e-15, 2.605604e-15, 
    2.788557e-15, 2.490461e-15, 2.243531e-15, 1.958471e-15, 1.5018e-15, 
    1.59995e-15, 1.265811e-15, 8.282425e-15, 7.575343e-15, 7.635848e-15, 
    6.940495e-15, 6.457008e-15, 5.494379e-15, 4.174979e-15, 4.640409e-15, 
    3.812842e-15, 3.660593e-15, 4.929404e-15, 4.118036e-15, 7.127722e-15, 
    6.557677e-15, 6.892946e-15, 8.224881e-15, 4.52987e-15, 6.225532e-15, 
    3.380983e-15, 4.088021e-15, 2.277608e-15, 3.083045e-15, 1.655879e-15, 
    1.222297e-15, 8.94437e-16, 5.963338e-16, 7.20886e-15, 7.667319e-15, 
    6.861047e-15, 5.850257e-15, 5.014319e-15, 4.042063e-15, 3.951036e-15, 
    3.788141e-15, 3.388919e-15, 3.077543e-15, 3.737602e-15, 3.002851e-15, 
    6.430217e-15, 4.4007e-15, 7.846011e-15, 6.653107e-15, 5.906644e-15, 
    6.226187e-15, 4.695924e-15, 4.379555e-15, 3.250859e-15, 3.803967e-15, 
    1.320688e-15, 2.193651e-15, 4.22506e-16, 7.288196e-16, 7.832418e-15, 
    7.210453e-15, 5.325213e-15, 6.170178e-15, 3.982513e-15, 3.545238e-15, 
    3.216312e-15, 2.828558e-15, 2.788856e-15, 2.577875e-15, 2.92993e-15, 
    2.59119e-15, 4.040153e-15, 3.335213e-15, 5.520051e-15, 4.913421e-15, 
    5.186129e-15, 5.497719e-15, 4.577739e-15, 3.726466e-15, 3.709745e-15, 
    3.46376e-15, 2.833828e-15, 3.975017e-15, 1.229791e-15, 2.653412e-15, 
    6.574451e-15, 5.552626e-15, 5.416968e-15, 5.79106e-15, 3.587425e-15, 
    4.298472e-15, 2.582887e-15, 2.985715e-15, 2.347131e-15, 2.650651e-15, 
    2.697566e-15, 3.132949e-15, 3.428299e-15, 4.263783e-15, 5.045399e-15, 
    5.735684e-15, 5.569391e-15, 4.830913e-15, 3.678467e-15, 2.785241e-15, 
    2.965758e-15, 2.391848e-15, 4.118432e-15, 3.311845e-15, 3.60854e-15, 
    2.872432e-15, 4.653242e-15, 3.098387e-15, 5.127529e-15, 4.919155e-15, 
    4.313544e-15, 3.26159e-15, 3.05683e-15, 2.848453e-15, 2.975797e-15, 
    3.652128e-15, 3.772713e-15, 4.327612e-15, 4.490654e-15, 4.963996e-15, 
    5.382497e-15, 4.999127e-15, 4.618333e-15, 3.651864e-15, 2.914637e-15, 
    2.240137e-15, 2.093934e-15, 1.487998e-15, 1.969826e-15, 1.223898e-15, 
    1.841508e-15, 8.776711e-16, 3.02193e-15, 1.862599e-15, 4.287386e-15, 
    3.953554e-15, 3.398062e-15, 2.339259e-15, 2.875616e-15, 2.256102e-15, 
    3.777503e-15, 4.806722e-15, 5.103332e-15, 5.691831e-15, 5.090422e-15, 
    5.137524e-15, 4.603117e-15, 4.77021e-15, 3.622543e-15, 4.210514e-15, 
    2.69873e-15, 2.260598e-15, 1.298237e-15, 8.790702e-16, 5.613584e-16, 
    4.511528e-16, 4.209018e-16, 4.086898e-16,
  4.033582e-20, 3.344133e-20, 3.470789e-20, 2.967473e-20, 3.239529e-20, 
    2.920249e-20, 3.886064e-20, 3.31867e-20, 3.673254e-20, 3.967606e-20, 
    2.145906e-20, 2.946358e-20, 1.495704e-20, 1.874748e-20, 1.032122e-20, 
    1.550648e-20, 9.451181e-21, 1.045052e-20, 7.652363e-21, 8.391163e-21, 
    5.447169e-21, 7.32751e-21, 4.252981e-21, 5.860896e-21, 5.584964e-21, 
    7.396378e-21, 2.770215e-20, 2.235647e-20, 2.804551e-20, 2.722404e-20, 
    2.759056e-20, 3.233708e-20, 3.494364e-20, 4.09032e-20, 3.976951e-20, 
    3.541817e-20, 2.686047e-20, 2.957258e-20, 2.309326e-20, 2.322691e-20, 
    1.727834e-20, 1.980264e-20, 1.157684e-20, 1.359766e-20, 8.359356e-21, 
    9.50874e-21, 8.410961e-21, 8.733759e-21, 8.406812e-21, 1.013612e-20, 
    9.366871e-21, 1.099463e-20, 1.931066e-20, 1.651129e-20, 2.585853e-20, 
    3.306083e-20, 3.859764e-20, 4.292137e-20, 4.228937e-20, 4.110355e-20, 
    3.539378e-20, 3.058057e-20, 2.724938e-20, 2.517484e-20, 2.324616e-20, 
    1.806077e-20, 1.568627e-20, 1.119597e-20, 1.192744e-20, 1.070777e-20, 
    9.628939e-21, 7.995301e-21, 8.249479e-21, 7.581729e-21, 1.073894e-20, 
    8.554101e-21, 1.235903e-20, 1.121776e-20, 2.27393e-20, 2.88221e-20, 
    3.173624e-20, 3.446165e-20, 4.180811e-20, 3.662342e-20, 3.860681e-20, 
    3.40133e-20, 3.131185e-20, 3.262749e-20, 2.511979e-20, 2.786846e-20, 
    1.555304e-20, 2.022487e-20, 9.750575e-21, 1.177461e-20, 9.305216e-21, 
    1.051339e-20, 8.506191e-21, 1.029882e-20, 7.3434e-21, 6.790702e-21, 
    7.165054e-21, 5.803022e-21, 1.040544e-20, 8.410882e-21, 3.266482e-20, 
    3.244733e-20, 3.144834e-20, 3.601451e-20, 3.630895e-20, 4.093448e-20, 
    3.679898e-20, 3.513487e-20, 3.116043e-20, 2.897085e-20, 2.699627e-20, 
    2.300299e-20, 1.907223e-20, 1.442456e-20, 1.163501e-20, 9.997154e-21, 
    1.098038e-20, 1.010892e-20, 1.108649e-20, 1.156727e-20, 6.994155e-21, 
    9.359847e-21, 5.986544e-21, 6.146132e-21, 7.566304e-21, 6.128003e-21, 
    3.229528e-20, 3.355714e-20, 3.822074e-20, 3.453324e-20, 4.146327e-20, 
    3.746884e-20, 3.530483e-20, 2.780842e-20, 2.633297e-20, 2.501621e-20, 
    2.255817e-20, 1.966731e-20, 1.525912e-20, 1.204755e-20, 9.568713e-21, 
    9.736687e-21, 9.677306e-21, 9.173823e-21, 1.045654e-20, 8.97456e-21, 
    8.741366e-21, 9.360266e-21, 6.167728e-21, 6.984786e-21, 6.149557e-21, 
    6.672284e-21, 3.314312e-20, 3.105953e-20, 3.217303e-20, 3.010271e-20, 
    3.155053e-20, 2.54835e-20, 2.384435e-20, 1.717515e-20, 1.972137e-20, 
    1.578672e-20, 1.929247e-20, 1.86337e-20, 1.566829e-20, 1.908993e-20, 
    1.22104e-20, 1.662929e-20, 9.15464e-21, 1.277519e-20, 8.955653e-21, 
    9.578568e-21, 8.56335e-21, 7.721299e-21, 6.74785e-21, 5.184794e-21, 
    5.521147e-21, 4.375006e-21, 2.813432e-20, 2.575785e-20, 2.596132e-20, 
    2.36218e-20, 2.199341e-20, 1.874664e-20, 1.428491e-20, 1.586054e-20, 
    1.305772e-20, 1.254139e-20, 1.68379e-20, 1.409201e-20, 2.4252e-20, 
    2.233258e-20, 2.346172e-20, 2.794102e-20, 1.548651e-20, 2.121326e-20, 
    1.159243e-20, 1.399033e-20, 7.837567e-21, 1.058022e-20, 5.712705e-21, 
    4.22551e-21, 3.097023e-21, 2.067004e-21, 2.452505e-20, 2.606713e-20, 
    2.335432e-20, 1.99477e-20, 1.712495e-20, 1.383463e-20, 1.352618e-20, 
    1.297397e-20, 1.161938e-20, 1.056152e-20, 1.280259e-20, 1.030757e-20, 
    2.190313e-20, 1.50493e-20, 2.666787e-20, 2.265405e-20, 2.013792e-20, 
    2.121547e-20, 1.604834e-20, 1.497771e-20, 1.115049e-20, 1.302763e-20, 
    4.563458e-21, 7.551076e-21, 1.463983e-21, 2.52531e-21, 2.662218e-20, 
    2.453041e-20, 1.817538e-20, 2.102665e-20, 1.363285e-20, 1.215e-20, 
    1.103312e-20, 9.714696e-21, 9.579584e-21, 8.861197e-21, 1.005957e-20, 
    8.906556e-21, 1.382816e-20, 1.1437e-20, 1.883331e-20, 1.678387e-20, 
    1.770555e-20, 1.875792e-20, 1.56485e-20, 1.276482e-20, 1.270811e-20, 
    1.187346e-20, 9.732629e-21, 1.360745e-20, 4.25126e-21, 9.118478e-21, 
    2.238909e-20, 1.894328e-20, 1.848526e-20, 1.974798e-20, 1.229315e-20, 
    1.470317e-20, 8.878271e-21, 1.02493e-20, 8.074713e-21, 9.109075e-21, 
    9.268825e-21, 1.074984e-20, 1.175308e-20, 1.45857e-20, 1.722999e-20, 
    1.956113e-20, 1.899988e-20, 1.650489e-20, 1.260202e-20, 9.567281e-21, 
    1.018143e-20, 8.227196e-21, 1.409335e-20, 1.135764e-20, 1.236479e-20, 
    9.863978e-21, 1.590396e-20, 1.063237e-20, 1.750755e-20, 1.680325e-20, 
    1.475421e-20, 1.118694e-20, 1.04911e-20, 9.782391e-21, 1.021557e-20, 
    1.251267e-20, 1.292165e-20, 1.480184e-20, 1.535379e-20, 1.695485e-20, 
    1.836885e-20, 1.70736e-20, 1.578585e-20, 1.251177e-20, 1.000755e-20, 
    7.709719e-21, 7.210638e-21, 5.137474e-21, 6.786658e-21, 4.23101e-21, 
    6.347969e-21, 3.039203e-21, 1.037245e-20, 6.420096e-21, 1.466563e-20, 
    1.353471e-20, 1.165042e-20, 8.047866e-21, 9.874809e-21, 7.764194e-21, 
    1.29379e-20, 1.642309e-20, 1.742578e-20, 1.941314e-20, 1.738215e-20, 
    1.754132e-20, 1.573437e-20, 1.629961e-20, 1.24123e-20, 1.440528e-20, 
    9.272789e-21, 7.779534e-21, 4.486368e-21, 3.044028e-21, 1.945841e-21, 
    1.563516e-21, 1.458407e-21, 1.415954e-21,
  2.961579e-26, 2.457414e-26, 2.55006e-26, 2.181813e-26, 2.380889e-26, 
    2.147251e-26, 2.853735e-26, 2.438787e-26, 2.698131e-26, 2.913349e-26, 
    1.580156e-26, 2.16636e-26, 1.103304e-26, 1.381382e-26, 7.627164e-27, 
    1.14363e-26, 6.987229e-27, 7.722245e-27, 5.663203e-27, 6.207167e-27, 
    4.037843e-27, 5.423938e-27, 3.156261e-27, 4.343012e-27, 4.139496e-27, 
    5.474667e-27, 2.037426e-26, 1.645917e-26, 2.062562e-26, 2.002424e-26, 
    2.029257e-26, 2.37663e-26, 2.567303e-26, 3.003054e-26, 2.920181e-26, 
    2.602009e-26, 1.975806e-26, 2.174337e-26, 1.699899e-26, 1.709691e-26, 
    1.273635e-26, 1.458745e-26, 8.550265e-27, 1.003496e-26, 6.183754e-27, 
    7.029573e-27, 6.22174e-27, 6.459332e-27, 6.218686e-27, 7.491043e-27, 
    6.925202e-27, 8.122301e-27, 1.422676e-26, 1.217363e-26, 1.902441e-26, 
    2.429578e-26, 2.834507e-26, 3.150563e-26, 3.104373e-26, 3.017699e-26, 
    2.600226e-26, 2.248106e-26, 2.004279e-26, 1.852373e-26, 1.711102e-26, 
    1.331023e-26, 1.156825e-26, 8.27031e-27, 8.807931e-27, 7.911404e-27, 
    7.117997e-27, 5.915733e-27, 6.102866e-27, 5.611183e-27, 7.934319e-27, 
    6.327102e-27, 9.125071e-27, 8.286327e-27, 1.673967e-26, 2.119408e-26, 
    2.33267e-26, 2.532049e-26, 3.069197e-26, 2.690152e-26, 2.835177e-26, 
    2.499254e-26, 2.301617e-26, 2.397876e-26, 1.848341e-26, 2.049601e-26, 
    1.147048e-26, 1.489698e-26, 7.207472e-27, 8.695618e-27, 6.87984e-27, 
    7.768477e-27, 6.291838e-27, 7.610698e-27, 5.435643e-27, 5.028442e-27, 
    5.304264e-27, 4.300331e-27, 7.689102e-27, 6.221682e-27, 2.400608e-26, 
    2.384696e-26, 2.311604e-26, 2.645622e-26, 2.667155e-26, 3.005341e-26, 
    2.70299e-26, 2.58129e-26, 2.290537e-26, 2.130296e-26, 1.985748e-26, 
    1.693286e-26, 1.405195e-26, 1.064216e-26, 8.593019e-27, 7.388839e-27, 
    8.111825e-27, 7.471041e-27, 8.189835e-27, 8.543229e-27, 5.178355e-27, 
    6.920034e-27, 4.435668e-27, 4.553338e-27, 5.599823e-27, 4.539971e-27, 
    2.373572e-26, 2.465886e-26, 2.80695e-26, 2.537286e-26, 3.043993e-26, 
    2.751973e-26, 2.59372e-26, 2.045206e-26, 1.937182e-26, 1.840755e-26, 
    1.660696e-26, 1.448824e-26, 1.125476e-26, 8.896192e-27, 7.073693e-27, 
    7.197256e-27, 7.153576e-27, 6.783166e-27, 7.726674e-27, 6.636542e-27, 
    6.464931e-27, 6.920342e-27, 4.56926e-27, 5.171452e-27, 4.555862e-27, 
    4.941176e-27, 2.435599e-26, 2.283154e-26, 2.364627e-26, 2.213135e-26, 
    2.319081e-26, 1.874978e-26, 1.754922e-26, 1.266065e-26, 1.452788e-26, 
    1.164196e-26, 1.421343e-26, 1.373039e-26, 1.155505e-26, 1.406492e-26, 
    9.015864e-27, 1.226021e-26, 6.769051e-27, 9.430821e-27, 6.622629e-27, 
    7.080943e-27, 6.33391e-27, 5.71397e-27, 4.996864e-27, 3.84425e-27, 
    4.092419e-27, 3.246399e-27, 2.069063e-26, 1.895069e-26, 1.909968e-26, 
    1.73862e-26, 1.619314e-26, 1.381321e-26, 1.053963e-26, 1.169614e-26, 
    9.638376e-27, 9.259056e-27, 1.241325e-26, 1.0398e-26, 1.784783e-26, 
    1.644167e-26, 1.726893e-26, 2.054913e-26, 1.142165e-26, 1.562143e-26, 
    8.561722e-27, 1.032334e-26, 5.799589e-27, 7.817617e-27, 4.233719e-27, 
    3.135966e-27, 2.30157e-27, 1.538392e-27, 1.804782e-26, 1.917716e-26, 
    1.719025e-26, 1.46938e-26, 1.262383e-26, 1.0209e-26, 9.982461e-27, 
    9.576853e-27, 8.581527e-27, 7.803865e-27, 9.450953e-27, 7.61713e-27, 
    1.612699e-26, 1.110076e-26, 1.961704e-26, 1.667721e-26, 1.483324e-26, 
    1.562305e-26, 1.183395e-26, 1.104821e-26, 8.236876e-27, 9.616272e-27, 
    3.38558e-27, 5.588608e-27, 1.090552e-27, 1.878207e-27, 1.958358e-26, 
    1.805175e-26, 1.339429e-26, 1.548466e-26, 1.006081e-26, 8.971479e-27, 
    8.150595e-27, 7.18108e-27, 7.08169e-27, 6.553118e-27, 7.434747e-27, 
    6.586499e-27, 1.020425e-26, 8.447485e-27, 1.387676e-26, 1.237361e-26, 
    1.30497e-26, 1.382148e-26, 1.154053e-26, 9.423206e-27, 9.381542e-27, 
    8.768262e-27, 7.194271e-27, 1.004215e-26, 3.154989e-27, 6.742443e-27, 
    1.648307e-26, 1.39574e-26, 1.362154e-26, 1.454738e-26, 9.076667e-27, 
    1.084669e-26, 6.565683e-27, 7.574277e-27, 5.974202e-27, 6.735524e-27, 
    6.853066e-27, 7.942333e-27, 8.679791e-27, 1.076045e-26, 1.270088e-26, 
    1.44104e-26, 1.399889e-26, 1.216894e-26, 9.303601e-27, 7.07264e-27, 
    7.524366e-27, 6.086463e-27, 1.039899e-26, 8.38915e-27, 9.129306e-27, 
    7.290886e-27, 1.1728e-26, 7.855963e-27, 1.290447e-26, 1.238783e-26, 
    1.088416e-26, 8.263674e-27, 7.752088e-27, 7.230875e-27, 7.549474e-27, 
    9.237956e-27, 9.538422e-27, 1.091912e-26, 1.132425e-26, 1.249904e-26, 
    1.353617e-26, 1.258616e-26, 1.164133e-26, 9.237299e-27, 7.396488e-27, 
    5.705443e-27, 5.337845e-27, 3.80933e-27, 5.025462e-27, 3.140029e-27, 
    4.702136e-27, 2.258776e-27, 7.664837e-27, 4.755303e-27, 1.081913e-26, 
    9.988729e-27, 8.604343e-27, 5.954435e-27, 7.298853e-27, 5.745559e-27, 
    9.550354e-27, 1.210891e-26, 1.28445e-26, 1.43019e-26, 1.28125e-26, 
    1.292925e-26, 1.160355e-26, 1.201831e-26, 9.164215e-27, 1.062801e-26, 
    6.855982e-27, 5.756855e-27, 3.32865e-27, 2.262348e-27, 1.448482e-27, 
    1.164538e-27, 1.086406e-27, 1.054839e-27,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_SAT =
  0.004421118, 0.004418409, 0.004418937, 0.00441675, 0.004417965, 
    0.004416532, 0.004420571, 0.0044183, 0.004419751, 0.004420877, 
    0.004412503, 0.004416653, 0.004408218, 0.004410858, 0.004404236, 
    0.004408626, 0.004403352, 0.004404367, 0.004401325, 0.004402197, 
    0.004398296, 0.004400922, 0.004396284, 0.004398926, 0.004398511, 
    0.004401008, 0.004415823, 0.004413018, 0.004415988, 0.004415588, 
    0.004415769, 0.004417938, 0.004419029, 0.004421329, 0.004420912, 
    0.004419225, 0.004415409, 0.004416707, 0.004413445, 0.004413519, 
    0.004409887, 0.004411524, 0.004405428, 0.004407161, 0.00440216, 
    0.004403417, 0.004402218, 0.004402582, 0.004402214, 0.004404056, 
    0.004403267, 0.00440489, 0.004411216, 0.004409355, 0.004414907, 
    0.004418242, 0.00442047, 0.004422049, 0.004421826, 0.004421399, 
    0.004419215, 0.004417166, 0.004415604, 0.004414558, 0.004413529, 
    0.004410403, 0.00440876, 0.004405076, 0.004405744, 0.004404615, 
    0.004403542, 0.004401735, 0.004402033, 0.004401236, 0.004404648, 
    0.004402379, 0.004406125, 0.004405099, 0.004413233, 0.004416357, 
    0.004417671, 0.004418835, 0.004421654, 0.004419706, 0.004420473, 
    0.004418652, 0.004417492, 0.004418066, 0.00441453, 0.004415904, 
    0.004408663, 0.00441178, 0.004403667, 0.004405607, 0.004403202, 
    0.00440443, 0.004402325, 0.00440422, 0.004400941, 0.004400226, 
    0.004400714, 0.004398843, 0.004404325, 0.004402217, 0.004418082, 
    0.004417988, 0.004417553, 0.004419464, 0.004419582, 0.004421339, 
    0.004419777, 0.004419111, 0.004417426, 0.004416427, 0.004415478, 
    0.004413394, 0.004411064, 0.004407813, 0.004405482, 0.004403919, 
    0.004404878, 0.004404031, 0.004404977, 0.004405422, 0.004400493, 
    0.004403258, 0.004399112, 0.004399342, 0.004401217, 0.004399316, 
    0.004417922, 0.004418461, 0.004420327, 0.004418867, 0.004421531, 
    0.004420037, 0.004419178, 0.004415872, 0.004415149, 0.004414475, 
    0.004413147, 0.00441144, 0.004408448, 0.004405849, 0.00440348, 
    0.004403654, 0.004403593, 0.004403062, 0.004404374, 0.004402847, 
    0.004402589, 0.004403261, 0.004399373, 0.004400483, 0.004399347, 
    0.004400071, 0.004418286, 0.00441738, 0.00441787, 0.004416949, 
    0.004417596, 0.004414713, 0.004413849, 0.004409813, 0.004411473, 
    0.004408835, 0.004411206, 0.004410785, 0.004408742, 0.004411079, 
    0.004405989, 0.004409433, 0.004403041, 0.004406471, 0.004402826, 
    0.00440349, 0.004402392, 0.004401407, 0.004400171, 0.004397887, 
    0.004398416, 0.00439651, 0.004416032, 0.004414856, 0.004414962, 
    0.004413734, 0.004412825, 0.00441086, 0.004407706, 0.004408893, 
    0.004406718, 0.00440628, 0.004409587, 0.004407553, 0.004414071, 
    0.004413014, 0.004413646, 0.004415937, 0.004408615, 0.004412369, 
    0.004405443, 0.004407475, 0.004401547, 0.004404491, 0.004398707, 
    0.004396229, 0.004393912, 0.004391189, 0.004414217, 0.004415016, 
    0.004413589, 0.004411609, 0.004409783, 0.00440735, 0.004407103, 
    0.004406647, 0.004405469, 0.004404477, 0.004406499, 0.004404229, 
    0.004412762, 0.004408291, 0.004415315, 0.004413194, 0.004411728, 
    0.004412374, 0.004409029, 0.00440824, 0.004405034, 0.004406693, 
    0.004396838, 0.004401194, 0.004389127, 0.004392494, 0.004415294, 
    0.004414221, 0.004410486, 0.004412263, 0.00440719, 0.00440594, 
    0.004404928, 0.004403629, 0.004403491, 0.004402722, 0.004403982, 
    0.004402773, 0.004407345, 0.004405302, 0.004410916, 0.004409547, 
    0.004410178, 0.004410868, 0.004408739, 0.004406467, 0.004406423, 
    0.004405694, 0.004403631, 0.004407169, 0.004396266, 0.004402987, 
    0.004413052, 0.00441098, 0.00441069, 0.004411492, 0.004406066, 
    0.00440803, 0.004402741, 0.004404171, 0.00440183, 0.004402993, 
    0.004403163, 0.004404658, 0.004405588, 0.004407939, 0.004409854, 
    0.004411376, 0.004411023, 0.004409351, 0.004406329, 0.004403476, 
    0.0044041, 0.004402008, 0.004407557, 0.004405227, 0.004406125, 
    0.004403783, 0.004408923, 0.00440453, 0.004410045, 0.004409562, 
    0.004408069, 0.004405065, 0.004404408, 0.004403698, 0.004404137, 
    0.004406253, 0.004406603, 0.004408107, 0.00440852, 0.004409668, 
    0.004410616, 0.004409749, 0.004408836, 0.004406255, 0.004403927, 
    0.004401392, 0.004400774, 0.004397803, 0.004400214, 0.004396228, 
    0.004399606, 0.004393764, 0.004404283, 0.004399716, 0.004408003, 
    0.004407111, 0.004405492, 0.004401792, 0.004403794, 0.004401455, 
    0.004406617, 0.004409291, 0.004409989, 0.004411282, 0.00440996, 
    0.004410068, 0.004408802, 0.004409209, 0.004406169, 0.004407802, 
    0.004403166, 0.004401475, 0.004396708, 0.004393784, 0.004390818, 
    0.004389506, 0.004389108, 0.004388941,
  8.305721e-06, 8.305594e-06, 8.305626e-06, 8.305499e-06, 8.30558e-06, 
    8.305487e-06, 8.305708e-06, 8.305578e-06, 8.305669e-06, 8.305726e-06, 
    8.305187e-06, 8.305496e-06, 8.304923e-06, 8.305136e-06, 8.304598e-06, 
    8.304943e-06, 8.304526e-06, 8.304633e-06, 8.304365e-06, 8.304445e-06, 
    8.304025e-06, 8.304327e-06, 8.303832e-06, 8.304112e-06, 8.30406e-06, 
    8.304332e-06, 8.30546e-06, 8.30522e-06, 8.305468e-06, 8.305436e-06, 
    8.305457e-06, 8.305569e-06, 8.305607e-06, 8.305748e-06, 8.305728e-06, 
    8.305632e-06, 8.305423e-06, 8.305515e-06, 8.305324e-06, 8.305329e-06, 
    8.30507e-06, 8.30519e-06, 8.304723e-06, 8.304871e-06, 8.304442e-06, 
    8.304552e-06, 8.304443e-06, 8.304481e-06, 8.304443e-06, 8.304604e-06, 
    8.304535e-06, 8.304681e-06, 8.305164e-06, 8.305024e-06, 8.3054e-06, 
    8.305552e-06, 8.305698e-06, 8.305776e-06, 8.305765e-06, 8.305739e-06, 
    8.305631e-06, 8.305539e-06, 8.305455e-06, 8.305391e-06, 8.305329e-06, 
    8.305062e-06, 8.304964e-06, 8.30468e-06, 8.304754e-06, 8.304643e-06, 
    8.304564e-06, 8.304397e-06, 8.304428e-06, 8.304347e-06, 8.304662e-06, 
    8.304448e-06, 8.304792e-06, 8.304699e-06, 8.305229e-06, 8.305494e-06, 
    8.305527e-06, 8.305617e-06, 8.305755e-06, 8.305658e-06, 8.305695e-06, 
    8.30562e-06, 8.305556e-06, 8.305591e-06, 8.30539e-06, 8.305468e-06, 
    8.304958e-06, 8.305195e-06, 8.304574e-06, 8.304741e-06, 8.304535e-06, 
    8.304646e-06, 8.304447e-06, 8.304627e-06, 8.304323e-06, 8.304243e-06, 
    8.304296e-06, 8.304119e-06, 8.304634e-06, 8.304436e-06, 8.305588e-06, 
    8.305582e-06, 8.305563e-06, 8.305644e-06, 8.305653e-06, 8.305744e-06, 
    8.305671e-06, 8.305631e-06, 8.305558e-06, 8.305497e-06, 8.305441e-06, 
    8.305313e-06, 8.305142e-06, 8.304904e-06, 8.30473e-06, 8.304602e-06, 
    8.304686e-06, 8.304611e-06, 8.304692e-06, 8.304733e-06, 8.304268e-06, 
    8.304529e-06, 8.304145e-06, 8.30417e-06, 8.304341e-06, 8.304168e-06, 
    8.305579e-06, 8.305612e-06, 8.305695e-06, 8.305631e-06, 8.305754e-06, 
    8.305677e-06, 8.305624e-06, 8.305449e-06, 8.305426e-06, 8.305379e-06, 
    8.305301e-06, 8.305184e-06, 8.304955e-06, 8.304752e-06, 8.304563e-06, 
    8.304579e-06, 8.304572e-06, 8.30452e-06, 8.304638e-06, 8.304502e-06, 
    8.30447e-06, 8.304539e-06, 8.304173e-06, 8.304282e-06, 8.30417e-06, 
    8.304244e-06, 8.305604e-06, 8.305551e-06, 8.305578e-06, 8.305522e-06, 
    8.305556e-06, 8.305376e-06, 8.305317e-06, 8.305044e-06, 8.305182e-06, 
    8.304982e-06, 8.305169e-06, 8.305132e-06, 8.30494e-06, 8.305165e-06, 
    8.304748e-06, 8.305006e-06, 8.304518e-06, 8.304768e-06, 8.3045e-06, 
    8.304564e-06, 8.304465e-06, 8.304365e-06, 8.304251e-06, 8.304006e-06, 
    8.304068e-06, 8.303869e-06, 8.305477e-06, 8.305395e-06, 8.305417e-06, 
    8.305338e-06, 8.305275e-06, 8.305147e-06, 8.304905e-06, 8.305004e-06, 
    8.304837e-06, 8.304796e-06, 8.305059e-06, 8.304886e-06, 8.305349e-06, 
    8.305266e-06, 8.305327e-06, 8.305461e-06, 8.30496e-06, 8.305225e-06, 
    8.304723e-06, 8.304891e-06, 8.304377e-06, 8.304628e-06, 8.304097e-06, 
    8.303804e-06, 8.304232e-06, 8.304897e-06, 8.305365e-06, 8.305421e-06, 
    8.305334e-06, 8.305175e-06, 8.305064e-06, 8.304878e-06, 8.304867e-06, 
    8.304825e-06, 8.304735e-06, 8.304649e-06, 8.304797e-06, 8.304629e-06, 
    8.305214e-06, 8.304943e-06, 8.305427e-06, 8.305274e-06, 8.305192e-06, 
    8.305244e-06, 8.305019e-06, 8.304957e-06, 8.304681e-06, 8.304835e-06, 
    8.303864e-06, 8.304321e-06, 8.305442e-06, 8.304572e-06, 8.305436e-06, 
    8.305373e-06, 8.305105e-06, 8.305239e-06, 8.304874e-06, 8.304767e-06, 
    8.304691e-06, 8.304563e-06, 8.304562e-06, 8.304486e-06, 8.304607e-06, 
    8.304497e-06, 8.304878e-06, 8.304716e-06, 8.305155e-06, 8.305047e-06, 
    8.305103e-06, 8.305152e-06, 8.304995e-06, 8.304791e-06, 8.304812e-06, 
    8.304739e-06, 8.304482e-06, 8.304873e-06, 8.303755e-06, 8.304436e-06, 
    8.305297e-06, 8.305126e-06, 8.305131e-06, 8.305195e-06, 8.304777e-06, 
    8.304934e-06, 8.304492e-06, 8.304623e-06, 8.304411e-06, 8.304516e-06, 
    8.30453e-06, 8.304665e-06, 8.304739e-06, 8.304922e-06, 8.305067e-06, 
    8.305188e-06, 8.305163e-06, 8.305028e-06, 8.304783e-06, 8.30455e-06, 
    8.3046e-06, 8.304429e-06, 8.304901e-06, 8.304699e-06, 8.304771e-06, 
    8.304585e-06, 8.305001e-06, 8.304574e-06, 8.305094e-06, 8.305056e-06, 
    8.304936e-06, 8.304668e-06, 8.304643e-06, 8.30457e-06, 8.304621e-06, 
    8.304782e-06, 8.304819e-06, 8.304945e-06, 8.304967e-06, 8.305066e-06, 
    8.305135e-06, 8.305066e-06, 8.304987e-06, 8.304793e-06, 8.304589e-06, 
    8.30436e-06, 8.304311e-06, 8.303955e-06, 8.304211e-06, 8.303745e-06, 
    8.304091e-06, 8.304194e-06, 8.304585e-06, 8.304153e-06, 8.304939e-06, 
    8.304869e-06, 8.30471e-06, 8.304374e-06, 8.304586e-06, 8.30435e-06, 
    8.304823e-06, 8.305011e-06, 8.305087e-06, 8.305176e-06, 8.305085e-06, 
    8.305095e-06, 8.305002e-06, 8.305034e-06, 8.304786e-06, 8.304923e-06, 
    8.304523e-06, 8.304358e-06, 8.30388e-06, 8.304236e-06, 8.305031e-06, 
    8.305358e-06, 8.305459e-06, 8.3055e-06,
  1.677104e-10, 1.677883e-10, 1.677733e-10, 1.67836e-10, 1.678015e-10, 
    1.678424e-10, 1.677265e-10, 1.677911e-10, 1.6775e-10, 1.677179e-10, 
    1.679575e-10, 1.678389e-10, 1.68085e-10, 1.68008e-10, 1.682031e-10, 
    1.680725e-10, 1.682297e-10, 1.682001e-10, 1.682913e-10, 1.682652e-10, 
    1.683808e-10, 1.683034e-10, 1.684423e-10, 1.683627e-10, 1.683749e-10, 
    1.683007e-10, 1.678634e-10, 1.679424e-10, 1.678585e-10, 1.678698e-10, 
    1.678649e-10, 1.678019e-10, 1.677698e-10, 1.67705e-10, 1.677169e-10, 
    1.677647e-10, 1.678749e-10, 1.678379e-10, 1.679328e-10, 1.679307e-10, 
    1.680366e-10, 1.679888e-10, 1.681685e-10, 1.681174e-10, 1.682663e-10, 
    1.682286e-10, 1.682644e-10, 1.682536e-10, 1.682645e-10, 1.682093e-10, 
    1.682329e-10, 1.681847e-10, 1.679976e-10, 1.680521e-10, 1.678897e-10, 
    1.677919e-10, 1.677292e-10, 1.676843e-10, 1.676907e-10, 1.677026e-10, 
    1.67765e-10, 1.678246e-10, 1.6787e-10, 1.679003e-10, 1.679304e-10, 
    1.680198e-10, 1.68069e-10, 1.681785e-10, 1.681593e-10, 1.681923e-10, 
    1.682249e-10, 1.682788e-10, 1.6827e-10, 1.682936e-10, 1.681919e-10, 
    1.682592e-10, 1.681483e-10, 1.681785e-10, 1.67936e-10, 1.67848e-10, 
    1.678086e-10, 1.677761e-10, 1.676955e-10, 1.67751e-10, 1.67729e-10, 
    1.677818e-10, 1.678152e-10, 1.677988e-10, 1.679012e-10, 1.678612e-10, 
    1.680719e-10, 1.679808e-10, 1.682211e-10, 1.681633e-10, 1.682351e-10, 
    1.681985e-10, 1.682609e-10, 1.682048e-10, 1.683026e-10, 1.683237e-10, 
    1.683092e-10, 1.683658e-10, 1.682016e-10, 1.682641e-10, 1.677982e-10, 
    1.678009e-10, 1.678135e-10, 1.677578e-10, 1.677546e-10, 1.677045e-10, 
    1.677493e-10, 1.677682e-10, 1.678173e-10, 1.678459e-10, 1.678734e-10, 
    1.67934e-10, 1.680016e-10, 1.680974e-10, 1.68167e-10, 1.682138e-10, 
    1.681853e-10, 1.682104e-10, 1.681822e-10, 1.681691e-10, 1.683156e-10, 
    1.68233e-10, 1.683576e-10, 1.683508e-10, 1.682941e-10, 1.683516e-10, 
    1.678028e-10, 1.677874e-10, 1.677334e-10, 1.677757e-10, 1.676991e-10, 
    1.677416e-10, 1.677659e-10, 1.678614e-10, 1.678832e-10, 1.679025e-10, 
    1.679414e-10, 1.679912e-10, 1.680788e-10, 1.681558e-10, 1.682269e-10, 
    1.682217e-10, 1.682235e-10, 1.682392e-10, 1.682001e-10, 1.682456e-10, 
    1.68253e-10, 1.682333e-10, 1.683499e-10, 1.683165e-10, 1.683507e-10, 
    1.68329e-10, 1.677925e-10, 1.678184e-10, 1.678044e-10, 1.678307e-10, 
    1.678119e-10, 1.678949e-10, 1.679199e-10, 1.68038e-10, 1.679901e-10, 
    1.680672e-10, 1.679981e-10, 1.680102e-10, 1.680687e-10, 1.68002e-10, 
    1.681511e-10, 1.680489e-10, 1.682398e-10, 1.681361e-10, 1.682462e-10, 
    1.682266e-10, 1.682594e-10, 1.682886e-10, 1.683258e-10, 1.683941e-10, 
    1.683783e-10, 1.68436e-10, 1.678575e-10, 1.678911e-10, 1.678886e-10, 
    1.679243e-10, 1.679506e-10, 1.680084e-10, 1.681009e-10, 1.680662e-10, 
    1.681306e-10, 1.681434e-10, 1.680459e-10, 1.681052e-10, 1.679141e-10, 
    1.679443e-10, 1.679266e-10, 1.678599e-10, 1.680736e-10, 1.679632e-10, 
    1.681681e-10, 1.681079e-10, 1.682843e-10, 1.681958e-10, 1.683696e-10, 
    1.684432e-10, 1.685323e-10, 1.686413e-10, 1.679101e-10, 1.678871e-10, 
    1.679287e-10, 1.679855e-10, 1.680398e-10, 1.681115e-10, 1.681191e-10, 
    1.681325e-10, 1.681677e-10, 1.681971e-10, 1.681362e-10, 1.682045e-10, 
    1.679503e-10, 1.680834e-10, 1.67878e-10, 1.679389e-10, 1.679823e-10, 
    1.679637e-10, 1.680624e-10, 1.680855e-10, 1.681799e-10, 1.681313e-10, 
    1.684246e-10, 1.682941e-10, 1.687262e-10, 1.685887e-10, 1.67879e-10, 
    1.679102e-10, 1.680187e-10, 1.679671e-10, 1.681166e-10, 1.681534e-10, 
    1.681838e-10, 1.68222e-10, 1.682265e-10, 1.682492e-10, 1.682119e-10, 
    1.682479e-10, 1.681116e-10, 1.681725e-10, 1.680069e-10, 1.680467e-10, 
    1.680285e-10, 1.680083e-10, 1.680708e-10, 1.681371e-10, 1.681393e-10, 
    1.681604e-10, 1.682188e-10, 1.681172e-10, 1.6844e-10, 1.682385e-10, 
    1.679443e-10, 1.680037e-10, 1.680132e-10, 1.679899e-10, 1.681496e-10, 
    1.680915e-10, 1.682487e-10, 1.682062e-10, 1.682762e-10, 1.682413e-10, 
    1.682361e-10, 1.681917e-10, 1.681639e-10, 1.68094e-10, 1.680376e-10, 
    1.679934e-10, 1.680037e-10, 1.680523e-10, 1.681413e-10, 1.682265e-10, 
    1.682077e-10, 1.682708e-10, 1.681056e-10, 1.681743e-10, 1.681475e-10, 
    1.682176e-10, 1.680651e-10, 1.681926e-10, 1.680325e-10, 1.680466e-10, 
    1.680903e-10, 1.681784e-10, 1.681991e-10, 1.682199e-10, 1.682073e-10, 
    1.681437e-10, 1.681337e-10, 1.680895e-10, 1.680769e-10, 1.680436e-10, 
    1.680157e-10, 1.68041e-10, 1.680674e-10, 1.681441e-10, 1.68213e-10, 
    1.682889e-10, 1.683078e-10, 1.68395e-10, 1.683229e-10, 1.68441e-10, 
    1.683389e-10, 1.685354e-10, 1.682011e-10, 1.683375e-10, 1.680926e-10, 
    1.68119e-10, 1.68166e-10, 1.68276e-10, 1.682173e-10, 1.682864e-10, 
    1.681333e-10, 1.680536e-10, 1.68034e-10, 1.67996e-10, 1.680349e-10, 
    1.680318e-10, 1.680691e-10, 1.680571e-10, 1.681466e-10, 1.680985e-10, 
    1.682358e-10, 1.68286e-10, 1.684296e-10, 1.685364e-10, 1.686578e-10, 
    1.687111e-10, 1.687274e-10, 1.687342e-10,
  4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 4.159382e-13, 
    4.159382e-13, 4.159382e-13, 4.159382e-13,
  4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 4.031953e-13, 
    4.031953e-13, 4.031953e-13, 4.031953e-13,
  3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 3.980121e-13, 
    3.980121e-13, 3.980121e-13, 3.980121e-13,
  3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 3.96582e-13, 
    3.96582e-13, 3.96582e-13, 3.96582e-13,
  3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 3.973374e-13, 
    3.973374e-13, 3.973374e-13, 3.973374e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CONC_O2_UNSAT =
  1.068899, 1.049683, 1.05342, 1.037911, 1.046516, 1.036359, 1.065005, 
    1.04892, 1.05919, 1.067171, 1.007782, 1.037219, 0.9771675, 0.9959709, 
    0.948707, 0.9800941, 0.9423731, 0.9496139, 0.9278157, 0.9340627, 
    0.9061567, 0.924932, 0.8916788, 0.9106424, 0.9076765, 0.9255509, 
    1.031299, 1.011449, 1.032475, 1.029645, 1.030915, 1.046338, 1.054106, 
    1.070368, 1.067417, 1.055473, 1.028373, 1.037576, 1.014376, 1.0149, 
    0.9890433, 1.000705, 0.9572017, 0.9695749, 0.9338021, 0.9428037, 
    0.9342248, 0.9368266, 0.9341909, 0.9473915, 0.9417366, 0.9533492, 
    0.9985214, 0.9852548, 1.024799, 1.048542, 1.0643, 1.075475, 1.073895, 
    1.070884, 1.055403, 1.040838, 1.029733, 1.022301, 1.014976, 0.9927861, 
    0.9810347, 0.9546984, 0.9594543, 0.9513975, 0.9436991, 0.9307671, 
    0.9328963, 0.9271967, 0.9516107, 0.9353878, 0.9621627, 0.9548425, 
    1.012981, 1.035094, 1.044484, 1.052702, 1.072681, 1.058885, 1.064325, 
    1.051383, 1.043156, 1.047225, 1.022097, 1.03187, 0.980338, 1.002549, 
    0.9445971, 0.9584783, 0.9412688, 0.9500522, 0.9350001, 0.9485474, 
    0.9250754, 0.9199609, 0.9234561, 0.9100279, 0.949298, 0.9342245, 
    1.047339, 1.046675, 1.043583, 1.057172, 1.058003, 1.070449, 1.059375, 
    1.054658, 1.042679, 1.03559, 1.028849, 1.014021, 0.9974489, 0.9742557, 
    0.9575787, 0.9463928, 0.9532527, 0.9471965, 0.9539664, 0.957139, 
    0.9218772, 0.9416837, 0.9119598, 0.9136056, 0.9270611, 0.9134202, 
    1.046209, 1.050028, 1.063282, 1.052911, 1.071804, 1.06123, 1.055148, 
    1.031665, 1.026503, 1.021714, 1.012255, 1.000108, 0.9787849, 0.9602156, 
    0.9432513, 0.9444947, 0.9440569, 0.9402653, 0.9496558, 0.9387233, 
    0.9368877, 0.9416864, 0.913826, 0.9217891, 0.9136406, 0.9188259, 
    1.048787, 1.042361, 1.045833, 1.039302, 1.043903, 1.023436, 1.017295, 
    0.9885418, 1.000347, 0.9815565, 0.9984396, 0.9954488, 0.9809421, 
    0.9975278, 0.9612393, 0.9858471, 0.9401179, 0.9647131, 0.9385757, 
    0.9433246, 0.9354616, 0.9284168, 0.9195514, 0.9031835, 0.9069749, 
    0.8932803, 1.032777, 1.024434, 1.025169, 1.016436, 1.009976, 0.9959666, 
    0.9734789, 0.981938, 0.9664065, 0.9632871, 0.9868825, 0.9723977, 1.01885, 
    1.011351, 1.015816, 1.032118, 0.9799882, 1.006756, 0.9573029, 0.9718226, 
    0.9294213, 0.9505177, 0.9090616, 0.8913147, 0.8746023, 0.8550528, 
    1.019881, 1.02555, 1.015398, 1.001343, 0.9882954, 0.9709371, 0.9691607, 
    0.9659069, 0.9574772, 0.9503868, 0.9648774, 0.9486091, 1.00961, 
    0.9776635, 1.027693, 1.012639, 1.002172, 1.006765, 0.9829047, 0.9772773, 
    0.9543952, 0.9662271, 0.8956956, 0.9269277, 0.8401586, 0.8644397, 
    1.027531, 1.0199, 0.9933223, 1.005972, 0.9697782, 0.96086, 0.953608, 
    0.9443334, 0.9433323, 0.9378352, 0.9468424, 0.9381913, 0.9709002, 
    0.9562892, 0.9963625, 0.9866151, 0.9911, 0.996018, 0.980836, 0.9646493, 
    0.9643041, 0.9591112, 0.9444696, 0.9696315, 0.8916597, 0.9398432, 
    1.011577, 0.9968649, 0.9947639, 1.000464, 0.9617542, 0.9757878, 
    0.9379693, 0.9481968, 0.9314371, 0.9397668, 0.9409919, 0.9516853, 
    0.95834, 0.9751444, 0.9888082, 0.9996377, 0.9971201, 0.9852225, 0.963659, 
    0.9432412, 0.9477153, 0.9327113, 0.9724045, 0.9557683, 0.9621994, 
    0.9454271, 0.9821625, 0.9508812, 0.990151, 0.9867109, 0.9760663, 
    0.9546389, 0.949897, 0.944831, 0.9479573, 0.9631115, 0.9655936, 
    0.9763253, 0.979287, 0.98746, 0.9942238, 0.9880438, 0.9815518, 0.9631054, 
    0.9464686, 0.9283164, 0.9238723, 0.9026382, 0.9199239, 0.8913909, 
    0.9156496, 0.8736408, 0.9490686, 0.9163645, 0.9755821, 0.9692101, 
    0.9576795, 0.9312127, 0.945506, 0.9287896, 0.9656909, 0.9848114, 
    0.9897569, 0.9989793, 0.9895461, 0.9903135, 0.9812834, 0.9841857, 
    0.9624927, 0.9741479, 0.9410225, 0.9289219, 0.8947155, 0.8737198, 
    0.8523293, 0.8428789, 0.8400019, 0.838799,
  0.4486648, 0.4327411, 0.4358204, 0.4230985, 0.4301388, 0.4218332, 
    0.4454201, 0.4321127, 0.440591, 0.4472236, 0.3988173, 0.4225344, 
    0.3747537, 0.3894614, 0.352949, 0.3770268, 0.3481727, 0.353636, 
    0.3373024, 0.3419491, 0.3214065, 0.3351667, 0.3109722, 0.3246713, 
    0.3225111, 0.3356245, 0.4177211, 0.4017409, 0.4186749, 0.4163797, 
    0.4174094, 0.4299924, 0.4363853, 0.4498917, 0.4474287, 0.4375146, 
    0.4153493, 0.4228259, 0.4040835, 0.4045032, 0.3840156, 0.3932016, 
    0.3593996, 0.3688836, 0.3417547, 0.3484972, 0.3420699, 0.3440138, 
    0.3420446, 0.3519554, 0.3476948, 0.3564684, 0.3914745, 0.3810507, 
    0.4124607, 0.4318009, 0.444833, 0.4541656, 0.4528419, 0.4503222, 
    0.4374568, 0.4254885, 0.4164512, 0.4104469, 0.4045636, 0.3869524, 
    0.3777591, 0.3574933, 0.3611186, 0.3549869, 0.349171, 0.339494, 
    0.3410792, 0.3368431, 0.3551491, 0.3429379, 0.3631898, 0.3576035, 
    0.4029645, 0.4208041, 0.4284706, 0.4352277, 0.4518251, 0.4403385, 
    0.4448535, 0.4341411, 0.427384, 0.4307212, 0.4102831, 0.418184, 
    0.3772169, 0.3946616, 0.3498473, 0.3603734, 0.3473435, 0.3539681, 
    0.3426484, 0.3528293, 0.3352726, 0.3314985, 0.3340755, 0.3242237, 
    0.3533971, 0.3420695, 0.4308146, 0.4302696, 0.4277344, 0.4389197, 
    0.4396077, 0.449959, 0.4407446, 0.4368416, 0.4269939, 0.4212076, 
    0.4157352, 0.4037992, 0.390627, 0.3724979, 0.3596871, 0.3512016, 
    0.3563954, 0.3518083, 0.3569375, 0.3593522, 0.3329102, 0.3476548, 
    0.325633, 0.326836, 0.3367425, 0.3267003, 0.4298871, 0.4330258, 0.443987, 
    0.4354002, 0.4510916, 0.4422825, 0.4372458, 0.4180171, 0.4138375, 
    0.4099745, 0.402387, 0.3927293, 0.37601, 0.3616999, 0.3488341, 0.3497703, 
    0.3494406, 0.34659, 0.3536679, 0.3454337, 0.3440591, 0.3476572, 
    0.3269972, 0.3328457, 0.3268616, 0.3306641, 0.4320047, 0.4267333, 
    0.4295787, 0.4242336, 0.4279962, 0.4113605, 0.4064218, 0.3836219, 
    0.3929183, 0.3781658, 0.39141, 0.3890499, 0.3776862, 0.3906901, 
    0.3624821, 0.3815128, 0.3464794, 0.365143, 0.3453231, 0.3488893, 
    0.3429935, 0.337748, 0.3311976, 0.3192517, 0.3220016, 0.3121193, 
    0.4189204, 0.4121664, 0.4127603, 0.4057341, 0.4005674, 0.3894583, 
    0.3718972, 0.3784636, 0.3664452, 0.3640509, 0.382324, 0.3710612, 
    0.4076705, 0.4016639, 0.4052368, 0.4183855, 0.376945, 0.3980023, 
    0.3594767, 0.3706174, 0.3384937, 0.3543198, 0.3235195, 0.3107112, 
    0.2988642, 0.28527, 0.4084991, 0.4130681, 0.4049019, 0.3937056, 
    0.3834297, 0.3699338, 0.3685644, 0.3660611, 0.3596099, 0.3542215, 
    0.36527, 0.352876, 0.4002738, 0.3751391, 0.4147996, 0.402693, 0.3943626, 
    0.3980096, 0.3792172, 0.3748401, 0.3572629, 0.3663073, 0.3138511, 
    0.3366431, 0.2751098, 0.291761, 0.4146688, 0.4085153, 0.3873753, 
    0.3973795, 0.3690403, 0.3621927, 0.3566652, 0.3496484, 0.348895, 
    0.3447684, 0.351541, 0.3450352, 0.3699053, 0.3587045, 0.3897707, 
    0.3821145, 0.3856295, 0.389499, 0.3776056, 0.3650948, 0.3648309, 
    0.3608561, 0.3497483, 0.3689272, 0.3109563, 0.3462709, 0.4018454, 
    0.3901658, 0.3885105, 0.3930111, 0.3628768, 0.3736848, 0.3448689, 
    0.3525642, 0.3399927, 0.3462161, 0.3471355, 0.3552057, 0.3602678, 
    0.3731861, 0.3838313, 0.3923573, 0.3903684, 0.3810256, 0.3643354, 
    0.3488261, 0.3521997, 0.3409415, 0.371067, 0.3583076, 0.3632173, 
    0.3504729, 0.3786383, 0.3545935, 0.3848847, 0.3821896, 0.3739006, 
    0.3574477, 0.3538505, 0.3500234, 0.3523832, 0.3639159, 0.3658203, 
    0.3741016, 0.3764004, 0.3827759, 0.3880855, 0.3832328, 0.3781623, 
    0.3639116, 0.3512583, 0.3376733, 0.3343833, 0.3188559, 0.3314704, 
    0.3107639, 0.3283293, 0.298187, 0.353222, 0.328855, 0.3735257, 0.3686026, 
    0.3597632, 0.3398246, 0.3505324, 0.3380241, 0.3658951, 0.3807041, 
    0.3845755, 0.3918366, 0.3844101, 0.3850121, 0.3779539, 0.3802165, 
    0.3634423, 0.3724151, 0.3471583, 0.3381225, 0.3131483, 0.2982436, 
    0.2834002, 0.2769531, 0.2750041, 0.2741911,
  0.2043858, 0.1962332, 0.1978064, 0.1913176, 0.1949051, 0.1906739, 0.202721, 
    0.1959123, 0.2002468, 0.2036462, 0.1790125, 0.1910306, 0.1669241, 
    0.1742999, 0.1560656, 0.1680614, 0.1536995, 0.1564063, 0.1483316, 
    0.1506233, 0.1405254, 0.1472797, 0.1354304, 0.1421244, 0.1410662, 
    0.1475051, 0.1885835, 0.1804885, 0.1890681, 0.1879023, 0.1884252, 
    0.1948303, 0.1980951, 0.2050157, 0.2037514, 0.1986726, 0.1873791, 
    0.1911789, 0.1816725, 0.1818846, 0.1715642, 0.176182, 0.1592683, 
    0.1639919, 0.1505273, 0.1538601, 0.1506829, 0.151643, 0.1506704, 
    0.155573, 0.153463, 0.157812, 0.1753125, 0.1700771, 0.1859138, 0.1957532, 
    0.20242, 0.2072121, 0.2065315, 0.2052368, 0.198643, 0.1925345, 0.1879386, 
    0.184893, 0.1819152, 0.1730387, 0.168428, 0.158321, 0.1601232, 0.1570765, 
    0.1541937, 0.1494119, 0.1501939, 0.1481053, 0.157157, 0.1511115, 
    0.161154, 0.1583757, 0.1811067, 0.1901505, 0.1940542, 0.1975034, 
    0.2060089, 0.2001175, 0.2024305, 0.1969482, 0.1935003, 0.1952022, 
    0.1848101, 0.1888187, 0.1681566, 0.1769173, 0.1545286, 0.1597525, 
    0.1532892, 0.1565711, 0.1509685, 0.1560063, 0.1473319, 0.1454753, 
    0.1467427, 0.1419051, 0.1562878, 0.1506827, 0.1952499, 0.1949718, 
    0.1936789, 0.1993914, 0.1997434, 0.2050503, 0.2003254, 0.1983284, 
    0.1933015, 0.1903557, 0.187575, 0.1815287, 0.1748861, 0.1657965, 
    0.1594113, 0.1551995, 0.1577757, 0.1555002, 0.1580449, 0.1592448, 
    0.1461694, 0.1534432, 0.1425959, 0.1431859, 0.1480557, 0.1431193, 
    0.1947767, 0.1963786, 0.2019864, 0.1975916, 0.2056321, 0.201113, 
    0.1985351, 0.1887339, 0.186612, 0.1846537, 0.1808151, 0.1759442, 
    0.1675526, 0.1604124, 0.1540269, 0.1544905, 0.1543272, 0.1529165, 
    0.1564221, 0.1523447, 0.1516653, 0.1534444, 0.143265, 0.1461377, 
    0.1431984, 0.1450653, 0.1958573, 0.1931687, 0.1946193, 0.1918955, 
    0.1938124, 0.185356, 0.182855, 0.1713666, 0.1760393, 0.1686317, 
    0.1752801, 0.1740929, 0.1683915, 0.1749179, 0.1608016, 0.1703087, 
    0.1528618, 0.1621267, 0.15229, 0.1540542, 0.151139, 0.1485511, 0.1453275, 
    0.1394714, 0.1408168, 0.1359893, 0.1891928, 0.1857645, 0.1860657, 
    0.1825071, 0.179896, 0.1742983, 0.1654965, 0.1687808, 0.1627757, 
    0.1615827, 0.1707155, 0.1650789, 0.1834869, 0.1804497, 0.1822556, 
    0.188921, 0.1680205, 0.1786015, 0.1593067, 0.1648573, 0.1489187, 
    0.1567455, 0.1415601, 0.1353031, 0.1295474, 0.122981, 0.1839065, 
    0.1862218, 0.1820862, 0.1764357, 0.1712702, 0.164516, 0.1638326, 
    0.1625843, 0.1593729, 0.1566968, 0.16219, 0.1560294, 0.1797477, 
    0.1671169, 0.1871002, 0.1809696, 0.1767667, 0.1786052, 0.1691583, 
    0.1669674, 0.1582065, 0.162707, 0.1368338, 0.1480067, 0.1181009, 
    0.1261111, 0.1870338, 0.1839147, 0.1732513, 0.1782874, 0.1640701, 
    0.1606576, 0.1579097, 0.1544301, 0.154057, 0.1520158, 0.1553677, 
    0.1521477, 0.1645018, 0.1589228, 0.1744554, 0.1706104, 0.1723744, 
    0.1743188, 0.1683512, 0.1621027, 0.1619713, 0.1599926, 0.1544794, 
    0.1640136, 0.1354225, 0.1527585, 0.1805415, 0.1746541, 0.1738218, 
    0.1760861, 0.1609982, 0.1663897, 0.1520655, 0.1558748, 0.1496579, 
    0.1527315, 0.1531863, 0.1571851, 0.1597001, 0.1661405, 0.1714717, 
    0.1757569, 0.1747561, 0.1700645, 0.1617244, 0.1540229, 0.1556941, 
    0.150126, 0.1650818, 0.1587256, 0.1611676, 0.1548384, 0.1688683, 
    0.1568812, 0.1720004, 0.1706481, 0.1664976, 0.1582983, 0.1565127, 
    0.1546157, 0.1557851, 0.1615155, 0.1624643, 0.1665981, 0.1677479, 
    0.1709422, 0.1736082, 0.1711714, 0.1686299, 0.1615134, 0.1552276, 
    0.1485143, 0.1468942, 0.1392778, 0.1454615, 0.1353287, 0.1439185, 
    0.1292192, 0.1562009, 0.1441766, 0.1663102, 0.1638517, 0.1594491, 
    0.1495749, 0.1548679, 0.1486872, 0.1625016, 0.1699033, 0.1718452, 
    0.1754948, 0.1717622, 0.1720644, 0.1685256, 0.169659, 0.1612797, 
    0.1657552, 0.1531975, 0.1487357, 0.136491, 0.1292467, 0.1220811, 
    0.1189845, 0.1180503, 0.1176608,
  0.04993047, 0.04752967, 0.0479911, 0.04609365, 0.04714081, 0.04590623, 
    0.04943832, 0.04743567, 0.04870865, 0.04971169, 0.04253784, 0.04601007, 
    0.03910066, 0.04119113, 0.03606242, 0.0394216, 0.03540676, 0.03615704, 
    0.03392795, 0.03455782, 0.03179934, 0.03363961, 0.03042435, 0.03223322, 
    0.03194596, 0.03370136, 0.0452987, 0.04296136, 0.04543941, 0.04510107, 
    0.04525276, 0.04711895, 0.04807588, 0.05011695, 0.04974281, 0.04824555, 
    0.04494942, 0.04605326, 0.04330169, 0.04336274, 0.04041328, 0.04172795, 
    0.03695359, 0.03827553, 0.03453139, 0.03545121, 0.03457424, 0.03483878, 
    0.0345708, 0.03592574, 0.03534136, 0.03654784, 0.0414798, 0.03999167, 
    0.04452515, 0.04738905, 0.04934943, 0.05076825, 0.05056626, 0.05018244, 
    0.04823686, 0.04644834, 0.0451116, 0.04423009, 0.04337152, 0.04083217, 
    0.03952516, 0.03668956, 0.03719216, 0.03634327, 0.03554352, 0.0342246, 
    0.03443964, 0.03386588, 0.03636565, 0.03469227, 0.03748024, 0.0367048, 
    0.043139, 0.04575396, 0.04689201, 0.04790217, 0.05041126, 0.04867058, 
    0.04935254, 0.04773929, 0.0467302, 0.04722775, 0.04420613, 0.04536698, 
    0.03944848, 0.04193806, 0.03563625, 0.03708868, 0.03529331, 0.0362028, 
    0.0346529, 0.03604596, 0.03365389, 0.03314606, 0.03349257, 0.03217364, 
    0.03612413, 0.03457417, 0.0472417, 0.04716032, 0.04678238, 0.04845688, 
    0.04856048, 0.05012719, 0.0487318, 0.04814442, 0.04667216, 0.04581365, 
    0.0450062, 0.04326034, 0.0413582, 0.03878295, 0.03699347, 0.03582216, 
    0.03653776, 0.03590553, 0.03661269, 0.03694702, 0.03333575, 0.03533589, 
    0.03236136, 0.03252184, 0.03385228, 0.03250374, 0.04710324, 0.04757228, 
    0.04922143, 0.04792806, 0.05029955, 0.04896384, 0.04820515, 0.04534236, 
    0.04472722, 0.04416096, 0.04305518, 0.04166005, 0.03927795, 0.03727294, 
    0.03549735, 0.0356257, 0.03558047, 0.0351903, 0.03616143, 0.03503239, 
    0.03484495, 0.03533622, 0.03254337, 0.03332708, 0.03252526, 0.0330341, 
    0.04741955, 0.04663339, 0.04705723, 0.04626201, 0.04682136, 0.04436387, 
    0.04364213, 0.04035721, 0.04168721, 0.03958272, 0.04147055, 0.04113219, 
    0.03951483, 0.04136725, 0.03738172, 0.04005728, 0.03517519, 0.03775247, 
    0.0350173, 0.03550492, 0.03469986, 0.0339882, 0.03310568, 0.03151395, 
    0.03187832, 0.03057464, 0.04547564, 0.04448199, 0.04456912, 0.04354192, 
    0.04279124, 0.0411907, 0.03869849, 0.03962488, 0.03793433, 0.03760019, 
    0.04017258, 0.03858102, 0.04382428, 0.04295022, 0.0434695, 0.0453967, 
    0.03941005, 0.04242004, 0.03696429, 0.03851871, 0.03408911, 0.03625127, 
    0.03207996, 0.03039017, 0.02885124, 0.02711422, 0.04394528, 0.04461427, 
    0.04342075, 0.04180043, 0.04032987, 0.03842277, 0.03823083, 0.03788066, 
    0.03698276, 0.03623772, 0.03777021, 0.03605239, 0.04274869, 0.03915503, 
    0.04486859, 0.04309959, 0.041895, 0.0424211, 0.03973163, 0.03911286, 
    0.03665768, 0.03791507, 0.03080193, 0.03383884, 0.02583653, 0.02793973, 
    0.04484937, 0.04394764, 0.04089263, 0.04233006, 0.03829749, 0.03734147, 
    0.03657505, 0.03560897, 0.0355057, 0.03494163, 0.03586879, 0.03497803, 
    0.03841877, 0.03685726, 0.04123545, 0.04014279, 0.04064335, 0.04119653, 
    0.03950346, 0.03774575, 0.03770895, 0.0371557, 0.03562262, 0.03828165, 
    0.03042223, 0.03514665, 0.04297657, 0.04129206, 0.04105499, 0.04170056, 
    0.03743666, 0.03895003, 0.03495535, 0.03600948, 0.03429221, 0.03513921, 
    0.03526487, 0.03637347, 0.03707404, 0.03887981, 0.04038704, 0.04160659, 
    0.04132112, 0.03998811, 0.03763983, 0.03549625, 0.03595933, 0.03442095, 
    0.03858184, 0.03680227, 0.03748405, 0.03572209, 0.03964962, 0.03628897, 
    0.04053713, 0.04015348, 0.03898044, 0.03668324, 0.03618659, 0.03566039, 
    0.03598459, 0.03758137, 0.03784703, 0.03900876, 0.03933309, 0.04023684, 
    0.04099419, 0.04030184, 0.03958222, 0.03758078, 0.03582994, 0.0339781, 
    0.03353402, 0.03146158, 0.03314226, 0.03039704, 0.03272133, 0.02876394, 
    0.03609999, 0.03279169, 0.03892763, 0.03823617, 0.03700401, 0.0342694, 
    0.03573026, 0.03402554, 0.03785748, 0.03994247, 0.04049306, 0.04153179, 
    0.04046949, 0.0405553, 0.03955275, 0.03987331, 0.03751539, 0.03877132, 
    0.03526797, 0.03403886, 0.03070964, 0.02877126, 0.02687777, 0.02606703, 
    0.02582333, 0.02572187,
  0.004358431, 0.0040972, 0.004147128, 0.003942681, 0.004055228, 0.003922612, 
    0.004304588, 0.004087045, 0.004225036, 0.004334477, 0.003565839, 
    0.003933729, 0.003209692, 0.003425325, 0.002901867, 0.003242597, 
    0.00283633, 0.002911351, 0.002689714, 0.002751958, 0.002481662, 
    0.002661322, 0.002349204, 0.002523777, 0.002495877, 0.002667397, 
    0.003857713, 0.003610284, 0.003872723, 0.003836653, 0.003852815, 
    0.004052872, 0.004156317, 0.004378871, 0.004337882, 0.004174718, 
    0.003820509, 0.003938355, 0.003646086, 0.003652516, 0.003344733, 
    0.003481188, 0.002991459, 0.00312543, 0.00274934, 0.002840763, 
    0.002753584, 0.002779821, 0.002753243, 0.002888179, 0.002829811, 
    0.002950595, 0.00345534, 0.003301226, 0.003775427, 0.004082011, 
    0.00429488, 0.004450427, 0.004428207, 0.004386054, 0.004173776, 
    0.003980724, 0.003837774, 0.003744143, 0.003653441, 0.003388082, 
    0.003253231, 0.002964854, 0.003015542, 0.002930038, 0.002849974, 
    0.00271899, 0.002740256, 0.002683597, 0.002932285, 0.002765284, 
    0.003044679, 0.002966389, 0.003628961, 0.003906324, 0.004028424, 
    0.004137495, 0.004411174, 0.004220894, 0.004295219, 0.004119865, 
    0.004011013, 0.004064604, 0.003741605, 0.003864995, 0.003245357, 
    0.003503106, 0.002859232, 0.003005091, 0.002825024, 0.002915941, 
    0.00276138, 0.002900218, 0.002662727, 0.002612876, 0.002646869, 
    0.002517985, 0.002908052, 0.002753578, 0.004066108, 0.004057332, 
    0.004016626, 0.004197664, 0.004208922, 0.004379994, 0.004227555, 
    0.004163748, 0.004004772, 0.003912707, 0.003826552, 0.003641732, 
    0.003442689, 0.00317719, 0.002995481, 0.002877814, 0.00294958, 
    0.002886156, 0.002957118, 0.002990796, 0.002631473, 0.002829267, 
    0.002536245, 0.002551878, 0.002682257, 0.002550113, 0.004051179, 
    0.004101805, 0.004280907, 0.0041403, 0.004398907, 0.004252821, 
    0.004170335, 0.003862369, 0.003796885, 0.003736822, 0.003620146, 
    0.003474112, 0.00322786, 0.003023706, 0.002845366, 0.002858178, 
    0.002853663, 0.002814765, 0.002911792, 0.002799056, 0.002780433, 
    0.002829299, 0.002553976, 0.002630623, 0.002552211, 0.002601912, 
    0.004085304, 0.004000604, 0.00404622, 0.003960729, 0.00402082, 
    0.00375832, 0.003681976, 0.00333894, 0.003476942, 0.003259145, 
    0.003454378, 0.003419204, 0.003252171, 0.003443631, 0.003034707, 
    0.003307988, 0.002813261, 0.003072269, 0.002797556, 0.002846121, 
    0.002766036, 0.002695655, 0.00260892, 0.002454042, 0.002489317, 
    0.002363607, 0.00387659, 0.003770847, 0.003780093, 0.003671404, 
    0.003592418, 0.00342528, 0.003168562, 0.003263478, 0.003090729, 
    0.003056828, 0.003319879, 0.00315657, 0.00370121, 0.003609114, 
    0.003663767, 0.003868165, 0.003241412, 0.003553499, 0.002992538, 
    0.003150213, 0.002705611, 0.002920803, 0.002508884, 0.002345931, 
    0.002199586, 0.002036844, 0.003714, 0.003784886, 0.003658628, 
    0.003488746, 0.003336115, 0.00314043, 0.003120878, 0.003085279, 
    0.002994401, 0.002919444, 0.003074068, 0.002900862, 0.003587951, 
    0.003215262, 0.003811912, 0.003624816, 0.003498612, 0.003553611, 
    0.003274454, 0.003210942, 0.002961644, 0.003088773, 0.002385423, 
    0.002680933, 0.001918846, 0.002113857, 0.003809867, 0.003714251, 
    0.003394349, 0.00354408, 0.003127666, 0.003030636, 0.002953331, 
    0.002856508, 0.002846199, 0.002790035, 0.002882479, 0.002793652, 
    0.003140023, 0.002981746, 0.00342993, 0.003316806, 0.003368526, 
    0.003425886, 0.003251003, 0.003071587, 0.003067854, 0.003011859, 
    0.002857871, 0.003126053, 0.002349001, 0.002810421, 0.003611882, 
    0.003435813, 0.003411189, 0.003478333, 0.003040267, 0.003194274, 
    0.002791398, 0.002896564, 0.002725673, 0.002809681, 0.002822191, 
    0.002933071, 0.003003613, 0.003187092, 0.003342021, 0.003468542, 
    0.003438834, 0.003300859, 0.003060847, 0.002845257, 0.002891542, 
    0.002738406, 0.003156653, 0.002976205, 0.003045065, 0.002867809, 
    0.003266021, 0.002924586, 0.003357536, 0.003317909, 0.003197385, 
    0.002964217, 0.002914315, 0.002861644, 0.00289407, 0.003054921, 
    0.003081865, 0.003200283, 0.003233515, 0.003326511, 0.00340488, 
    0.003333221, 0.003259094, 0.003054862, 0.002878593, 0.002694659, 
    0.002650942, 0.002448981, 0.002612503, 0.002346588, 0.002571337, 
    0.002191344, 0.002905632, 0.002578209, 0.003191982, 0.003121423, 
    0.002996545, 0.002723418, 0.002868625, 0.002699337, 0.003082926, 
    0.003296156, 0.003352979, 0.003460752, 0.003350543, 0.003359416, 
    0.003256065, 0.003289034, 0.003048238, 0.003176002, 0.002822499, 
    0.002700652, 0.00237656, 0.002192034, 0.002014897, 0.001940024, 
    0.001917635, 0.00190833,
  0.0001201083, 0.0001110804, 0.0001127942, 0.0001058123, 0.0001096441, 
    0.0001051321, 0.0001182353, 0.0001107326, 0.0001154795, 0.0001192743, 
    9.319912e-05, 0.0001055088, 8.160235e-05, 8.858483e-05, 7.18514e-05, 
    8.265997e-05, 6.980984e-05, 7.214787e-05, 6.528819e-05, 6.719997e-05, 
    5.898418e-05, 6.442003e-05, 5.504247e-05, 6.024935e-05, 5.941056e-05, 
    6.460559e-05, 0.0001029389, 9.466886e-05, 0.0001034452, 0.0001022292, 
    0.0001027737, 0.0001095636, 0.0001131102, 0.000120821, 0.0001193928, 
    0.0001137437, 0.000101686, 0.0001056656, 9.585632e-05, 9.606993e-05, 
    8.596098e-05, 9.041333e-05, 7.466222e-05, 7.890727e-05, 6.711934e-05, 
    6.994753e-05, 6.725009e-05, 6.805953e-05, 6.723959e-05, 7.142396e-05, 
    6.960744e-05, 7.337733e-05, 8.956629e-05, 8.45515e-05, 0.0001001723, 
    0.0001105602, 0.0001178983, 0.000123323, 0.0001225449, 0.0001210717, 
    0.0001137112, 0.0001071042, 0.000102267, 9.912467e-05, 9.610067e-05, 
    8.737022e-05, 8.300238e-05, 7.382513e-05, 7.542165e-05, 7.273276e-05, 
    7.023383e-05, 6.618595e-05, 6.683968e-05, 6.510093e-05, 7.280317e-05, 
    6.76108e-05, 7.634262e-05, 7.387337e-05, 9.528796e-05, 0.0001045807, 
    0.0001087289, 0.0001124631, 0.0001219491, 0.0001153364, 0.00011791, 
    0.0001118577, 0.0001081353, 0.0001099646, 9.903979e-05, 0.0001031845, 
    8.274881e-05, 9.113292e-05, 7.052186e-05, 7.509189e-05, 6.94589e-05, 
    7.229143e-05, 6.749039e-05, 7.179988e-05, 6.446292e-05, 6.294432e-05, 
    6.397903e-05, 6.007502e-05, 7.204472e-05, 6.724989e-05, 0.000110016, 
    0.000109716, 0.0001083266, 0.0001145346, 0.000114923, 0.0001208602, 
    0.0001155666, 0.000113366, 0.0001079227, 0.0001047967, 0.0001018893, 
    9.571174e-05, 8.915235e-05, 8.056051e-05, 7.478894e-05, 7.110067e-05, 
    7.33455e-05, 7.136085e-05, 7.358212e-05, 7.464133e-05, 6.350994e-05, 
    6.959055e-05, 6.062496e-05, 6.109662e-05, 6.505993e-05, 6.104333e-05, 
    0.0001095057, 0.0001112383, 0.0001174135, 0.0001125595, 0.0001215204, 
    0.0001164405, 0.0001135927, 0.0001030959, 0.0001008922, 9.887985e-05, 
    9.499563e-05, 9.018127e-05, 8.218594e-05, 7.567946e-05, 7.009059e-05, 
    7.048906e-05, 7.034856e-05, 6.914078e-05, 7.216165e-05, 6.865427e-05, 
    6.807844e-05, 6.959155e-05, 6.115999e-05, 6.348407e-05, 6.110667e-05, 
    6.261138e-05, 0.0001106729, 0.0001077807, 0.0001093363, 0.0001064248, 
    0.0001084696, 9.959913e-05, 9.704989e-05, 8.577301e-05, 9.027406e-05, 
    8.319291e-05, 8.953479e-05, 8.838497e-05, 8.296821e-05, 8.918315e-05, 
    7.602716e-05, 8.477022e-05, 6.909417e-05, 7.721684e-05, 6.860784e-05, 
    7.011405e-05, 6.763401e-05, 6.547016e-05, 6.282416e-05, 5.815756e-05, 
    5.921373e-05, 5.546827e-05, 0.0001035758, 0.0001000188, 0.0001003287, 
    9.669797e-05, 9.407743e-05, 8.858337e-05, 8.028442e-05, 8.33326e-05, 
    7.780297e-05, 7.672733e-05, 8.515517e-05, 7.990101e-05, 9.769083e-05, 
    9.463009e-05, 9.644393e-05, 0.0001032914, 8.262183e-05, 9.279189e-05, 
    7.46962e-05, 7.969792e-05, 6.577534e-05, 7.244359e-05, 5.98013e-05, 
    5.494579e-05, 5.066054e-05, 4.598314e-05, 9.81175e-05, 0.0001004895, 
    9.627308e-05, 9.066132e-05, 8.568139e-05, 7.938564e-05, 7.876223e-05, 
    7.762983e-05, 7.475491e-05, 7.240105e-05, 7.727394e-05, 7.182001e-05, 
    9.39297e-05, 8.178115e-05, 0.000101397, 9.515049e-05, 9.098528e-05, 
    9.279556e-05, 8.368663e-05, 8.164245e-05, 7.37243e-05, 7.774082e-05, 
    5.611457e-05, 6.501942e-05, 4.265254e-05, 4.818475e-05, 0.0001013283, 
    9.812586e-05, 8.757436e-05, 9.248132e-05, 7.897854e-05, 7.589845e-05, 
    7.346323e-05, 7.043708e-05, 7.011648e-05, 6.837522e-05, 7.124614e-05, 
    6.848708e-05, 7.937263e-05, 7.435637e-05, 8.873525e-05, 8.505567e-05, 
    8.673387e-05, 8.860315e-05, 8.293059e-05, 7.719522e-05, 7.707681e-05, 
    7.53054e-05, 7.047949e-05, 7.892711e-05, 5.503645e-05, 6.900617e-05, 
    9.472181e-05, 8.892753e-05, 8.812341e-05, 9.03197e-05, 7.620301e-05, 
    8.110776e-05, 6.841736e-05, 7.168575e-05, 6.639124e-05, 6.898325e-05, 
    6.9371e-05, 7.282778e-05, 7.504526e-05, 8.087759e-05, 8.587298e-05, 
    8.999871e-05, 8.902628e-05, 8.453964e-05, 7.685467e-05, 7.008718e-05, 
    7.152894e-05, 6.678276e-05, 7.990369e-05, 7.418203e-05, 7.635482e-05, 
    7.07889e-05, 8.34146e-05, 7.256202e-05, 8.63767e-05, 8.509138e-05, 
    8.12075e-05, 7.380514e-05, 7.224058e-05, 7.059692e-05, 7.160788e-05, 
    7.666692e-05, 7.752142e-05, 8.130045e-05, 8.236777e-05, 8.537003e-05, 
    8.791764e-05, 8.558755e-05, 8.319127e-05, 7.666503e-05, 7.112494e-05, 
    6.543965e-05, 6.410325e-05, 5.800634e-05, 6.293301e-05, 5.496519e-05, 
    6.168481e-05, 5.042137e-05, 7.196907e-05, 6.18928e-05, 8.10343e-05, 
    7.877957e-05, 7.482246e-05, 6.632195e-05, 7.081433e-05, 6.558301e-05, 
    7.75551e-05, 8.438758e-05, 8.622868e-05, 8.974352e-05, 8.614957e-05, 
    8.643775e-05, 8.309368e-05, 8.415741e-05, 7.645528e-05, 8.052247e-05, 
    6.938059e-05, 6.562329e-05, 5.58518e-05, 5.044141e-05, 4.535971e-05, 
    4.324642e-05, 4.261864e-05, 4.235828e-05,
  9.233383e-07, 8.324391e-07, 8.495325e-07, 7.803872e-07, 8.181727e-07, 
    7.737215e-07, 9.043083e-07, 8.289789e-07, 8.764705e-07, 9.148534e-07, 
    6.589369e-07, 7.774109e-07, 5.5156e-07, 6.156955e-07, 4.647986e-07, 
    5.611706e-07, 4.470745e-07, 4.673857e-07, 4.083967e-07, 4.246511e-07, 
    3.558722e-07, 4.010644e-07, 3.23913e-07, 3.662774e-07, 3.593711e-07, 
    4.026289e-07, 7.523169e-07, 6.72848e-07, 7.572467e-07, 7.454205e-07, 
    7.507106e-07, 8.173747e-07, 8.52693e-07, 9.306024e-07, 9.160577e-07, 
    8.590354e-07, 7.401507e-07, 7.789482e-07, 6.841349e-07, 6.861698e-07, 
    5.914073e-07, 6.327512e-07, 4.894573e-07, 5.272426e-07, 4.239625e-07, 
    4.482649e-07, 4.250791e-07, 4.320067e-07, 4.249895e-07, 4.610747e-07, 
    4.453261e-07, 4.78149e-07, 6.248371e-07, 5.784527e-07, 7.255105e-07, 
    8.272655e-07, 9.008932e-07, 9.562033e-07, 9.482252e-07, 9.331602e-07, 
    8.587102e-07, 7.930824e-07, 7.45787e-07, 7.154174e-07, 6.864627e-07, 
    6.044247e-07, 5.642901e-07, 4.820832e-07, 4.961696e-07, 4.72499e-07, 
    4.507423e-07, 4.160114e-07, 4.215766e-07, 4.068125e-07, 4.731155e-07, 
    4.28163e-07, 5.043375e-07, 4.825075e-07, 6.787274e-07, 7.683277e-07, 
    8.091118e-07, 8.462242e-07, 9.421263e-07, 8.750303e-07, 9.010124e-07, 
    8.401822e-07, 8.032467e-07, 8.213514e-07, 7.14601e-07, 7.547071e-07, 
    5.619796e-07, 6.39492e-07, 4.53238e-07, 4.932524e-07, 4.440438e-07, 
    4.686395e-07, 4.27133e-07, 4.643494e-07, 4.014259e-07, 3.88672e-07, 
    3.973516e-07, 3.648396e-07, 4.664852e-07, 4.250774e-07, 8.218619e-07, 
    8.188856e-07, 8.051356e-07, 8.669696e-07, 8.708724e-07, 9.31002e-07, 
    8.773468e-07, 8.552522e-07, 8.011481e-07, 7.704396e-07, 7.421216e-07, 
    6.827584e-07, 6.209778e-07, 5.4213e-07, 4.905759e-07, 4.582627e-07, 
    4.778696e-07, 4.605254e-07, 4.799472e-07, 4.89273e-07, 3.934111e-07, 
    4.451801e-07, 3.693801e-07, 3.732846e-07, 4.064659e-07, 3.72843e-07, 
    8.168014e-07, 8.340102e-07, 8.959867e-07, 8.471868e-07, 9.377437e-07, 
    8.861554e-07, 8.57523e-07, 7.538447e-07, 7.324647e-07, 7.130633e-07, 
    6.759497e-07, 6.305807e-07, 5.568584e-07, 4.984529e-07, 4.495024e-07, 
    4.529536e-07, 4.517361e-07, 4.413008e-07, 4.675059e-07, 4.371132e-07, 
    4.321689e-07, 4.451888e-07, 3.738099e-07, 3.931941e-07, 3.733679e-07, 
    3.858886e-07, 8.28386e-07, 7.997479e-07, 8.151232e-07, 7.864001e-07, 
    8.065483e-07, 7.199847e-07, 6.955224e-07, 5.896759e-07, 6.314484e-07, 
    5.660277e-07, 6.245432e-07, 6.138376e-07, 5.639787e-07, 6.212647e-07, 
    5.015363e-07, 5.804587e-07, 4.408991e-07, 5.121191e-07, 4.367141e-07, 
    4.497055e-07, 4.283616e-07, 4.099375e-07, 3.876669e-07, 3.49112e-07, 
    3.577549e-07, 3.273312e-07, 7.585187e-07, 7.240296e-07, 7.270204e-07, 
    6.921605e-07, 6.672422e-07, 6.156818e-07, 5.396372e-07, 5.673024e-07, 
    5.173515e-07, 5.077585e-07, 5.839931e-07, 5.361798e-07, 7.016549e-07, 
    6.724802e-07, 6.897359e-07, 7.557485e-07, 5.608234e-07, 6.55094e-07, 
    4.897573e-07, 5.343506e-07, 4.125245e-07, 4.699693e-07, 3.625845e-07, 
    3.23138e-07, 2.89238e-07, 2.532848e-07, 7.05744e-07, 7.28573e-07, 
    6.881062e-07, 6.350724e-07, 5.888324e-07, 5.315405e-07, 5.25941e-07, 
    5.158046e-07, 4.902755e-07, 4.695974e-07, 5.126283e-07, 4.645249e-07, 
    6.658437e-07, 5.53182e-07, 7.3735e-07, 6.774209e-07, 6.381077e-07, 
    6.551286e-07, 5.705359e-07, 5.519237e-07, 4.811967e-07, 5.167961e-07, 
    3.325354e-07, 4.061234e-07, 2.283984e-07, 2.700662e-07, 7.366846e-07, 
    7.058241e-07, 6.063156e-07, 6.521668e-07, 5.278824e-07, 5.003944e-07, 
    4.78903e-07, 4.52503e-07, 4.497264e-07, 4.347156e-07, 4.595275e-07, 
    4.356762e-07, 5.314235e-07, 4.867601e-07, 6.170945e-07, 5.83079e-07, 
    5.985386e-07, 6.158658e-07, 5.636358e-07, 5.119263e-07, 5.108708e-07, 
    4.951407e-07, 4.528706e-07, 5.274206e-07, 3.238647e-07, 4.401412e-07, 
    6.733503e-07, 6.18884e-07, 6.114082e-07, 6.318752e-07, 5.030974e-07, 
    5.470786e-07, 4.350774e-07, 4.633546e-07, 4.177571e-07, 4.399438e-07, 
    4.432855e-07, 4.733309e-07, 4.928402e-07, 5.449961e-07, 5.905966e-07, 
    6.288744e-07, 6.198035e-07, 5.783438e-07, 5.08892e-07, 4.494729e-07, 
    4.619886e-07, 4.210913e-07, 5.362039e-07, 4.852241e-07, 5.044459e-07, 
    4.555545e-07, 5.680511e-07, 4.71005e-07, 5.952407e-07, 5.83407e-07, 
    5.479817e-07, 4.819074e-07, 4.681953e-07, 4.538889e-07, 4.626762e-07, 
    5.072209e-07, 5.148365e-07, 5.488236e-07, 5.585116e-07, 5.859679e-07, 
    6.094984e-07, 5.879687e-07, 5.660127e-07, 5.072042e-07, 4.584736e-07, 
    4.09679e-07, 3.983965e-07, 3.478785e-07, 3.885773e-07, 3.232935e-07, 
    3.781672e-07, 2.873724e-07, 4.658251e-07, 3.798972e-07, 5.464137e-07, 
    5.260965e-07, 4.908719e-07, 4.171677e-07, 4.557753e-07, 4.108937e-07, 
    5.151372e-07, 5.769502e-07, 5.938751e-07, 6.26491e-07, 5.931456e-07, 
    5.958041e-07, 5.651226e-07, 5.748421e-07, 5.053388e-07, 5.417863e-07, 
    4.433682e-07, 4.112351e-07, 3.304172e-07, 2.875286e-07, 2.485799e-07, 
    2.327904e-07, 2.281483e-07, 2.262296e-07,
  1.115461e-09, 9.230383e-10, 9.583536e-10, 8.181131e-10, 8.93884e-10, 
    8.049692e-10, 1.074252e-09, 9.159404e-10, 1.014839e-09, 1.097028e-09, 
    5.898345e-10, 8.122358e-10, 4.098776e-10, 5.14698e-10, 2.820693e-10, 
    4.250549e-10, 2.581446e-10, 2.856267e-10, 2.087564e-10, 2.290275e-10, 
    1.483791e-10, 1.998494e-10, 1.157796e-10, 1.596904e-10, 1.521455e-10, 
    2.017374e-10, 7.632262e-10, 6.14726e-10, 7.727771e-10, 7.499299e-10, 
    7.601227e-10, 8.92262e-10, 9.649287e-10, 1.131315e-09, 1.099639e-09, 
    9.78165e-10, 7.398208e-10, 8.152696e-10, 6.351707e-10, 6.388801e-10, 
    4.740395e-10, 5.43922e-10, 3.166351e-10, 3.723505e-10, 2.281544e-10, 
    2.597266e-10, 2.29571e-10, 2.384341e-10, 2.294571e-10, 2.769775e-10, 
    2.558274e-10, 3.006022e-10, 5.302938e-10, 4.528265e-10, 7.119698e-10, 
    9.12432e-10, 1.066907e-09, 1.187732e-09, 1.170061e-09, 1.136914e-09, 
    9.774848e-10, 8.43333e-10, 7.506346e-10, 6.929723e-10, 6.394147e-10, 
    4.956887e-10, 4.300227e-10, 3.061456e-10, 3.262942e-10, 2.927061e-10, 
    2.630308e-10, 2.181635e-10, 2.251385e-10, 2.068194e-10, 2.935639e-10, 
    2.335007e-10, 3.381888e-10, 3.067456e-10, 6.253483e-10, 7.943832e-10, 
    8.755215e-10, 9.514863e-10, 1.156607e-09, 1.011794e-09, 1.067163e-09, 
    9.389843e-10, 8.636993e-10, 9.003545e-10, 6.91443e-10, 7.678521e-10, 
    4.263414e-10, 5.556215e-10, 2.663749e-10, 3.220834e-10, 2.54133e-10, 
    2.873567e-10, 2.321854e-10, 2.814532e-10, 2.00285e-10, 1.8514e-10, 
    1.953967e-10, 1.581076e-10, 2.843866e-10, 2.295688e-10, 9.013949e-10, 
    8.95334e-10, 8.675012e-10, 9.948022e-10, 1.003018e-09, 1.132189e-09, 
    1.016693e-09, 9.702625e-10, 8.594818e-10, 7.985226e-10, 7.435963e-10, 
    6.326655e-10, 5.236906e-10, 3.951744e-10, 3.182375e-10, 2.731554e-10, 
    3.002099e-10, 2.762294e-10, 3.031313e-10, 3.163714e-10, 1.907136e-10, 
    2.556343e-10, 1.631273e-10, 1.674935e-10, 2.063964e-10, 1.669975e-10, 
    8.910972e-10, 9.262667e-10, 1.056383e-09, 9.534827e-10, 1.146968e-09, 
    1.035391e-09, 9.750035e-10, 7.661821e-10, 7.251559e-10, 6.885655e-10, 
    6.203221e-10, 5.401729e-10, 4.182212e-10, 3.296039e-10, 2.613752e-10, 
    2.659931e-10, 2.643605e-10, 2.505224e-10, 2.857924e-10, 2.45048e-10, 
    2.38643e-10, 2.556458e-10, 1.680845e-10, 1.904569e-10, 1.675872e-10, 
    1.818967e-10, 9.147255e-10, 8.566714e-10, 8.876906e-10, 8.300277e-10, 
    8.703479e-10, 7.015483e-10, 6.560204e-10, 4.711851e-10, 5.416707e-10, 
    4.327984e-10, 5.2979e-10, 5.115478e-10, 4.295259e-10, 5.241805e-10, 
    3.340922e-10, 4.560894e-10, 2.499954e-10, 3.496625e-10, 2.445286e-10, 
    2.616461e-10, 2.337547e-10, 2.10647e-10, 1.839663e-10, 1.4121e-10, 
    1.50401e-10, 1.191069e-10, 7.752475e-10, 7.091719e-10, 7.148261e-10, 
    6.498419e-10, 6.046542e-10, 5.146748e-10, 3.913193e-10, 4.348385e-10, 
    3.574545e-10, 3.432161e-10, 4.618578e-10, 3.859947e-10, 6.673397e-10, 
    6.140632e-10, 6.45398e-10, 7.698704e-10, 4.245033e-10, 5.830189e-10, 
    3.170645e-10, 3.831879e-10, 2.138362e-10, 2.891958e-10, 1.556379e-10, 
    1.150306e-10, 8.430732e-11, 5.635257e-11, 6.749226e-10, 7.177671e-10, 
    6.424167e-10, 5.479414e-10, 4.697965e-10, 3.788903e-10, 3.70378e-10, 
    3.551445e-10, 3.178068e-10, 2.886811e-10, 3.504181e-10, 2.816939e-10, 
    6.021503e-10, 4.124256e-10, 7.34466e-10, 6.229824e-10, 5.53212e-10, 
    5.8308e-10, 4.400289e-10, 4.104484e-10, 3.048933e-10, 3.566246e-10, 
    1.242474e-10, 2.059789e-10, 4.003784e-11, 6.877948e-11, 7.331957e-10, 
    6.750714e-10, 4.988609e-10, 5.77845e-10, 3.733215e-10, 3.324274e-10, 
    3.016618e-10, 2.653884e-10, 2.61674e-10, 2.419341e-10, 2.748721e-10, 
    2.431799e-10, 3.787117e-10, 3.127835e-10, 5.170746e-10, 4.603636e-10, 
    4.858586e-10, 5.149871e-10, 4.289789e-10, 3.493767e-10, 3.478128e-10, 
    3.248068e-10, 2.658816e-10, 3.726206e-10, 1.157327e-10, 2.490019e-10, 
    6.156308e-10, 5.201198e-10, 5.074383e-10, 5.424078e-10, 3.36373e-10, 
    4.028669e-10, 2.42403e-10, 2.800908e-10, 2.203424e-10, 2.487434e-10, 
    2.531329e-10, 2.938639e-10, 3.214901e-10, 3.996232e-10, 4.727022e-10, 
    5.372316e-10, 5.216869e-10, 4.526497e-10, 3.448877e-10, 2.613358e-10, 
    2.782239e-10, 2.245269e-10, 3.860317e-10, 3.105977e-10, 3.383477e-10, 
    2.69493e-10, 4.360384e-10, 2.90631e-10, 4.803803e-10, 4.608996e-10, 
    4.042762e-10, 3.058971e-10, 2.867434e-10, 2.672497e-10, 2.79163e-10, 
    3.424243e-10, 3.537017e-10, 4.055916e-10, 4.208365e-10, 4.650918e-10, 
    5.042159e-10, 4.683763e-10, 4.327744e-10, 3.423996e-10, 2.734414e-10, 
    2.103294e-10, 1.96646e-10, 1.399175e-10, 1.850293e-10, 1.151806e-10, 
    1.730174e-10, 8.273571e-11, 2.834787e-10, 1.749917e-10, 4.018302e-10, 
    3.706135e-10, 3.18662e-10, 2.196058e-10, 2.697909e-10, 2.118236e-10, 
    3.541497e-10, 4.50388e-10, 4.781183e-10, 5.331323e-10, 4.769113e-10, 
    4.813147e-10, 4.313517e-10, 4.469743e-10, 3.396574e-10, 3.946422e-10, 
    2.532419e-10, 2.122443e-10, 1.221444e-10, 8.286685e-11, 5.307095e-11, 
    4.272747e-11, 3.98872e-11, 3.874047e-11,
  4.052103e-13, 4.044533e-13, 4.045923e-13, 4.040399e-13, 4.043385e-13, 
    4.039881e-13, 4.050483e-13, 4.044253e-13, 4.048146e-13, 4.051378e-13, 
    4.031391e-13, 4.040168e-13, 4.024272e-13, 4.028421e-13, 4.019204e-13, 
    4.024873e-13, 4.018254e-13, 4.019345e-13, 4.016291e-13, 4.017097e-13, 
    4.013887e-13, 4.015936e-13, 4.012588e-13, 4.014338e-13, 4.014037e-13, 
    4.016011e-13, 4.038236e-13, 4.032375e-13, 4.038612e-13, 4.037711e-13, 
    4.038113e-13, 4.043321e-13, 4.046182e-13, 4.052726e-13, 4.051481e-13, 
    4.046703e-13, 4.037312e-13, 4.040287e-13, 4.033182e-13, 4.033329e-13, 
    4.026813e-13, 4.029577e-13, 4.020576e-13, 4.022785e-13, 4.017062e-13, 
    4.018317e-13, 4.017118e-13, 4.01747e-13, 4.017114e-13, 4.019002e-13, 
    4.018162e-13, 4.019939e-13, 4.029038e-13, 4.025973e-13, 4.036214e-13, 
    4.044115e-13, 4.050194e-13, 4.054943e-13, 4.054249e-13, 4.052946e-13, 
    4.046676e-13, 4.041393e-13, 4.037739e-13, 4.035464e-13, 4.03335e-13, 
    4.027669e-13, 4.02507e-13, 4.02016e-13, 4.020959e-13, 4.019626e-13, 
    4.018448e-13, 4.016665e-13, 4.016942e-13, 4.016214e-13, 4.01966e-13, 
    4.017275e-13, 4.021431e-13, 4.020183e-13, 4.032794e-13, 4.039464e-13, 
    4.042661e-13, 4.045653e-13, 4.05372e-13, 4.048026e-13, 4.050204e-13, 
    4.04516e-13, 4.042196e-13, 4.04364e-13, 4.035404e-13, 4.038418e-13, 
    4.024924e-13, 4.030039e-13, 4.018581e-13, 4.020792e-13, 4.018094e-13, 
    4.019414e-13, 4.017222e-13, 4.019179e-13, 4.015954e-13, 4.015351e-13, 
    4.015759e-13, 4.014275e-13, 4.019296e-13, 4.017118e-13, 4.043681e-13, 
    4.043442e-13, 4.042346e-13, 4.047358e-13, 4.047681e-13, 4.05276e-13, 
    4.048219e-13, 4.046392e-13, 4.04203e-13, 4.039627e-13, 4.037462e-13, 
    4.033083e-13, 4.028777e-13, 4.023689e-13, 4.020639e-13, 4.01885e-13, 
    4.019924e-13, 4.018972e-13, 4.02004e-13, 4.020565e-13, 4.015573e-13, 
    4.018154e-13, 4.014475e-13, 4.014649e-13, 4.016197e-13, 4.014629e-13, 
    4.043275e-13, 4.04466e-13, 4.04978e-13, 4.045731e-13, 4.053341e-13, 
    4.048954e-13, 4.046578e-13, 4.038352e-13, 4.036734e-13, 4.03529e-13, 
    4.032596e-13, 4.029428e-13, 4.024602e-13, 4.02109e-13, 4.018382e-13, 
    4.018566e-13, 4.018501e-13, 4.017951e-13, 4.019352e-13, 4.017733e-13, 
    4.017479e-13, 4.018154e-13, 4.014672e-13, 4.015563e-13, 4.014652e-13, 
    4.015222e-13, 4.044206e-13, 4.041919e-13, 4.043141e-13, 4.040869e-13, 
    4.042458e-13, 4.035802e-13, 4.034006e-13, 4.026699e-13, 4.029488e-13, 
    4.02518e-13, 4.029018e-13, 4.028297e-13, 4.02505e-13, 4.028796e-13, 
    4.021268e-13, 4.026102e-13, 4.01793e-13, 4.021886e-13, 4.017713e-13, 
    4.018393e-13, 4.017285e-13, 4.016366e-13, 4.015304e-13, 4.013602e-13, 
    4.013968e-13, 4.01272e-13, 4.03871e-13, 4.036103e-13, 4.036326e-13, 
    4.033762e-13, 4.031977e-13, 4.02842e-13, 4.023537e-13, 4.02526e-13, 
    4.022195e-13, 4.02163e-13, 4.02633e-13, 4.023326e-13, 4.034452e-13, 
    4.032349e-13, 4.033586e-13, 4.038498e-13, 4.024851e-13, 4.031122e-13, 
    4.020593e-13, 4.023214e-13, 4.016493e-13, 4.019487e-13, 4.014176e-13, 
    4.012558e-13, 4.011332e-13, 4.010215e-13, 4.034752e-13, 4.036442e-13, 
    4.033468e-13, 4.029736e-13, 4.026644e-13, 4.023044e-13, 4.022707e-13, 
    4.022103e-13, 4.020622e-13, 4.019466e-13, 4.021916e-13, 4.019189e-13, 
    4.031878e-13, 4.024373e-13, 4.037101e-13, 4.032701e-13, 4.029944e-13, 
    4.031124e-13, 4.025466e-13, 4.024294e-13, 4.02011e-13, 4.022162e-13, 
    4.012925e-13, 4.01618e-13, 4.009562e-13, 4.010711e-13, 4.037051e-13, 
    4.034758e-13, 4.027795e-13, 4.030918e-13, 4.022823e-13, 4.021202e-13, 
    4.019982e-13, 4.018541e-13, 4.018394e-13, 4.01761e-13, 4.018918e-13, 
    4.017659e-13, 4.023037e-13, 4.020423e-13, 4.028515e-13, 4.026271e-13, 
    4.02728e-13, 4.028433e-13, 4.025028e-13, 4.021874e-13, 4.021812e-13, 
    4.0209e-13, 4.018561e-13, 4.022796e-13, 4.012586e-13, 4.017891e-13, 
    4.032411e-13, 4.028636e-13, 4.028134e-13, 4.029517e-13, 4.021359e-13, 
    4.023994e-13, 4.017628e-13, 4.019125e-13, 4.016751e-13, 4.01788e-13, 
    4.018055e-13, 4.019672e-13, 4.020768e-13, 4.023866e-13, 4.026759e-13, 
    4.029312e-13, 4.028697e-13, 4.025966e-13, 4.021696e-13, 4.01838e-13, 
    4.019051e-13, 4.016918e-13, 4.023327e-13, 4.020336e-13, 4.021437e-13, 
    4.018705e-13, 4.025308e-13, 4.019544e-13, 4.027064e-13, 4.026292e-13, 
    4.02405e-13, 4.02015e-13, 4.01939e-13, 4.018615e-13, 4.019088e-13, 
    4.021599e-13, 4.022046e-13, 4.024102e-13, 4.024706e-13, 4.026458e-13, 
    4.028006e-13, 4.026588e-13, 4.025179e-13, 4.021598e-13, 4.018861e-13, 
    4.016353e-13, 4.015809e-13, 4.01355e-13, 4.015347e-13, 4.012564e-13, 
    4.014868e-13, 4.011269e-13, 4.01926e-13, 4.014947e-13, 4.023953e-13, 
    4.022716e-13, 4.020656e-13, 4.016722e-13, 4.018716e-13, 4.016413e-13, 
    4.022063e-13, 4.025876e-13, 4.026974e-13, 4.02915e-13, 4.026926e-13, 
    4.0271e-13, 4.025123e-13, 4.025741e-13, 4.021489e-13, 4.023668e-13, 
    4.018059e-13, 4.016429e-13, 4.012841e-13, 4.011274e-13, 4.010084e-13, 
    4.00967e-13, 4.009556e-13, 4.00951e-13,
  4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 4.008e-13, 
    4.008e-13, 4.008e-13,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC =
  8.949659e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 
    8.949658e-07, 8.949659e-07, 8.949658e-07, 8.949658e-07, 8.949659e-07, 
    8.949657e-07, 8.949658e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 
    8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949654e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949655e-07, 8.949658e-07, 8.949657e-07, 8.949658e-07, 8.949658e-07, 
    8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949659e-07, 8.949659e-07, 
    8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949657e-07, 8.949657e-07, 
    8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949656e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949656e-07, 8.949656e-07, 8.949658e-07, 
    8.949658e-07, 8.949659e-07, 8.949659e-07, 8.949659e-07, 8.949659e-07, 
    8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949657e-07, 8.949657e-07, 
    8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949657e-07, 8.949658e-07, 
    8.949658e-07, 8.949658e-07, 8.949659e-07, 8.949658e-07, 8.949659e-07, 
    8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949657e-07, 8.949658e-07, 
    8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949655e-07, 8.949655e-07, 8.949658e-07, 
    8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949659e-07, 
    8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 
    8.949657e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949655e-07, 8.949654e-07, 
    8.949658e-07, 8.949658e-07, 8.949659e-07, 8.949658e-07, 8.949659e-07, 
    8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949657e-07, 
    8.949657e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 
    8.949658e-07, 8.949658e-07, 8.949657e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949655e-07, 8.949656e-07, 8.949655e-07, 8.949656e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949654e-07, 8.949658e-07, 8.949658e-07, 8.949658e-07, 
    8.949657e-07, 8.949657e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949655e-07, 8.949656e-07, 8.949656e-07, 8.949657e-07, 
    8.949657e-07, 8.949657e-07, 8.949658e-07, 8.949656e-07, 8.949657e-07, 
    8.949655e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949652e-07, 8.949657e-07, 8.949658e-07, 
    8.949657e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949656e-07, 8.949655e-07, 
    8.949657e-07, 8.949656e-07, 8.949658e-07, 8.949657e-07, 8.949656e-07, 
    8.949657e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949656e-07, 
    8.949654e-07, 8.949655e-07, 8.949652e-07, 8.949652e-07, 8.949658e-07, 
    8.949657e-07, 8.949656e-07, 8.949657e-07, 8.949656e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949656e-07, 8.949655e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949655e-07, 8.949655e-07, 8.949656e-07, 8.949654e-07, 8.949655e-07, 
    8.949657e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 
    8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949655e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949656e-07, 8.949655e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949655e-07, 
    8.949655e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 8.949654e-07, 
    8.949654e-07, 8.949653e-07, 8.949655e-07, 8.949654e-07, 8.949656e-07, 
    8.949656e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 8.949655e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949656e-07, 
    8.949656e-07, 8.949656e-07, 8.949656e-07, 8.949655e-07, 8.949656e-07, 
    8.949655e-07, 8.949655e-07, 8.949654e-07, 8.949653e-07, 8.949652e-07, 
    8.949652e-07, 8.949652e-07, 8.949652e-07 ;

 CWDC_HR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDC_LOSS =
  6.710401e-16, 6.728806e-16, 6.72523e-16, 6.740064e-16, 6.731839e-16, 
    6.741548e-16, 6.714136e-16, 6.729534e-16, 6.719707e-16, 6.712063e-16, 
    6.768815e-16, 6.740726e-16, 6.797985e-16, 6.780092e-16, 6.82502e-16, 
    6.795197e-16, 6.83103e-16, 6.824168e-16, 6.844832e-16, 6.838915e-16, 
    6.865311e-16, 6.847564e-16, 6.878991e-16, 6.861078e-16, 6.863878e-16, 
    6.846977e-16, 6.746388e-16, 6.765318e-16, 6.745264e-16, 6.747965e-16, 
    6.746755e-16, 6.732007e-16, 6.724567e-16, 6.708999e-16, 6.711827e-16, 
    6.723264e-16, 6.74918e-16, 6.74039e-16, 6.762549e-16, 6.762049e-16, 
    6.786691e-16, 6.775583e-16, 6.816966e-16, 6.805213e-16, 6.839162e-16, 
    6.830628e-16, 6.83876e-16, 6.836295e-16, 6.838792e-16, 6.826276e-16, 
    6.831639e-16, 6.820624e-16, 6.777663e-16, 6.790295e-16, 6.752595e-16, 
    6.729889e-16, 6.714811e-16, 6.704101e-16, 6.705616e-16, 6.708501e-16, 
    6.72333e-16, 6.73727e-16, 6.747887e-16, 6.754985e-16, 6.761977e-16, 
    6.783112e-16, 6.794306e-16, 6.819338e-16, 6.814828e-16, 6.822472e-16, 
    6.82978e-16, 6.842035e-16, 6.840019e-16, 6.845416e-16, 6.822274e-16, 
    6.837655e-16, 6.812258e-16, 6.819206e-16, 6.763855e-16, 6.742762e-16, 
    6.733772e-16, 6.725917e-16, 6.706779e-16, 6.719996e-16, 6.714786e-16, 
    6.727183e-16, 6.735054e-16, 6.731163e-16, 6.755179e-16, 6.745844e-16, 
    6.794969e-16, 6.773822e-16, 6.828927e-16, 6.815754e-16, 6.832084e-16, 
    6.823754e-16, 6.838023e-16, 6.825182e-16, 6.847426e-16, 6.852264e-16, 
    6.848957e-16, 6.861663e-16, 6.824469e-16, 6.838758e-16, 6.731053e-16, 
    6.731687e-16, 6.734646e-16, 6.721636e-16, 6.720842e-16, 6.70892e-16, 
    6.71953e-16, 6.724045e-16, 6.735512e-16, 6.742288e-16, 6.748729e-16, 
    6.762885e-16, 6.778681e-16, 6.800758e-16, 6.816608e-16, 6.827226e-16, 
    6.820717e-16, 6.826463e-16, 6.820039e-16, 6.817028e-16, 6.850449e-16, 
    6.831688e-16, 6.859836e-16, 6.85828e-16, 6.845543e-16, 6.858456e-16, 
    6.732133e-16, 6.72848e-16, 6.715787e-16, 6.725721e-16, 6.707622e-16, 
    6.717752e-16, 6.723573e-16, 6.746034e-16, 6.750972e-16, 6.755542e-16, 
    6.764572e-16, 6.776152e-16, 6.796451e-16, 6.814102e-16, 6.830205e-16, 
    6.829026e-16, 6.829441e-16, 6.833035e-16, 6.824129e-16, 6.834497e-16, 
    6.836234e-16, 6.831688e-16, 6.858072e-16, 6.850538e-16, 6.858247e-16, 
    6.853343e-16, 6.729668e-16, 6.735815e-16, 6.732493e-16, 6.738738e-16, 
    6.734337e-16, 6.753893e-16, 6.759753e-16, 6.787162e-16, 6.775923e-16, 
    6.793813e-16, 6.777742e-16, 6.78059e-16, 6.794387e-16, 6.778613e-16, 
    6.813124e-16, 6.789724e-16, 6.833175e-16, 6.809819e-16, 6.834637e-16, 
    6.830136e-16, 6.83759e-16, 6.844261e-16, 6.852655e-16, 6.868128e-16, 
    6.864547e-16, 6.877483e-16, 6.744977e-16, 6.752943e-16, 6.752246e-16, 
    6.760582e-16, 6.766744e-16, 6.7801e-16, 6.801499e-16, 6.793456e-16, 
    6.808225e-16, 6.811187e-16, 6.788751e-16, 6.802525e-16, 6.758275e-16, 
    6.765426e-16, 6.761172e-16, 6.745604e-16, 6.795304e-16, 6.769808e-16, 
    6.816869e-16, 6.803075e-16, 6.843309e-16, 6.823305e-16, 6.862574e-16, 
    6.879328e-16, 6.895103e-16, 6.913499e-16, 6.757293e-16, 6.751882e-16, 
    6.761574e-16, 6.774969e-16, 6.787403e-16, 6.803916e-16, 6.805607e-16, 
    6.808698e-16, 6.816707e-16, 6.823436e-16, 6.809671e-16, 6.825123e-16, 
    6.767075e-16, 6.797517e-16, 6.749832e-16, 6.764195e-16, 6.774182e-16, 
    6.769806e-16, 6.792537e-16, 6.79789e-16, 6.819627e-16, 6.808395e-16, 
    6.875191e-16, 6.845664e-16, 6.927509e-16, 6.904667e-16, 6.74999e-16, 
    6.757277e-16, 6.782613e-16, 6.770563e-16, 6.80502e-16, 6.813492e-16, 
    6.82038e-16, 6.829175e-16, 6.830127e-16, 6.835337e-16, 6.826799e-16, 
    6.835002e-16, 6.803951e-16, 6.817833e-16, 6.779724e-16, 6.789002e-16, 
    6.784736e-16, 6.780051e-16, 6.794505e-16, 6.809887e-16, 6.810222e-16, 
    6.81515e-16, 6.82902e-16, 6.80516e-16, 6.878985e-16, 6.833411e-16, 
    6.765219e-16, 6.779235e-16, 6.781244e-16, 6.775815e-16, 6.812643e-16, 
    6.799304e-16, 6.835211e-16, 6.825514e-16, 6.841403e-16, 6.833508e-16, 
    6.832346e-16, 6.822204e-16, 6.815886e-16, 6.799915e-16, 6.786914e-16, 
    6.776603e-16, 6.779002e-16, 6.790327e-16, 6.810828e-16, 6.830211e-16, 
    6.825966e-16, 6.840196e-16, 6.802523e-16, 6.818324e-16, 6.812216e-16, 
    6.82814e-16, 6.793241e-16, 6.822943e-16, 6.78564e-16, 6.788914e-16, 
    6.79904e-16, 6.819391e-16, 6.823901e-16, 6.828703e-16, 6.825741e-16, 
    6.81135e-16, 6.808995e-16, 6.798795e-16, 6.795975e-16, 6.788202e-16, 
    6.781761e-16, 6.787644e-16, 6.793819e-16, 6.811359e-16, 6.82715e-16, 
    6.844355e-16, 6.848566e-16, 6.86863e-16, 6.852289e-16, 6.879238e-16, 
    6.856315e-16, 6.895987e-16, 6.824673e-16, 6.855654e-16, 6.799502e-16, 
    6.80556e-16, 6.816506e-16, 6.841604e-16, 6.828065e-16, 6.843902e-16, 
    6.808903e-16, 6.790714e-16, 6.786015e-16, 6.777229e-16, 6.786215e-16, 
    6.785485e-16, 6.79408e-16, 6.791319e-16, 6.811941e-16, 6.800866e-16, 
    6.832315e-16, 6.843778e-16, 6.876126e-16, 6.895926e-16, 6.916072e-16, 
    6.924956e-16, 6.92766e-16, 6.928789e-16 ;

 CWDC_TO_LITR2C =
  5.099905e-16, 5.113893e-16, 5.111175e-16, 5.122449e-16, 5.116198e-16, 
    5.123577e-16, 5.102744e-16, 5.114445e-16, 5.106978e-16, 5.101168e-16, 
    5.144299e-16, 5.122952e-16, 5.166468e-16, 5.15287e-16, 5.187015e-16, 
    5.16435e-16, 5.191583e-16, 5.186367e-16, 5.202073e-16, 5.197575e-16, 
    5.217636e-16, 5.204148e-16, 5.228033e-16, 5.214419e-16, 5.216548e-16, 
    5.203702e-16, 5.127255e-16, 5.141641e-16, 5.126401e-16, 5.128454e-16, 
    5.127534e-16, 5.116325e-16, 5.110671e-16, 5.098839e-16, 5.100989e-16, 
    5.10968e-16, 5.129376e-16, 5.122696e-16, 5.139537e-16, 5.139157e-16, 
    5.157885e-16, 5.149443e-16, 5.180893e-16, 5.171962e-16, 5.197763e-16, 
    5.191278e-16, 5.197458e-16, 5.195585e-16, 5.197482e-16, 5.187969e-16, 
    5.192046e-16, 5.183674e-16, 5.151024e-16, 5.160624e-16, 5.131973e-16, 
    5.114715e-16, 5.103257e-16, 5.095117e-16, 5.096268e-16, 5.098461e-16, 
    5.109731e-16, 5.120326e-16, 5.128394e-16, 5.133788e-16, 5.139102e-16, 
    5.155165e-16, 5.163673e-16, 5.182697e-16, 5.179269e-16, 5.185078e-16, 
    5.190632e-16, 5.199947e-16, 5.198415e-16, 5.202516e-16, 5.184928e-16, 
    5.196618e-16, 5.177316e-16, 5.182596e-16, 5.14053e-16, 5.1245e-16, 
    5.117667e-16, 5.111697e-16, 5.097153e-16, 5.107197e-16, 5.103237e-16, 
    5.112659e-16, 5.118641e-16, 5.115684e-16, 5.133936e-16, 5.126842e-16, 
    5.164177e-16, 5.148105e-16, 5.189985e-16, 5.179973e-16, 5.192384e-16, 
    5.186053e-16, 5.196898e-16, 5.187138e-16, 5.204043e-16, 5.207721e-16, 
    5.205208e-16, 5.214864e-16, 5.186597e-16, 5.197456e-16, 5.1156e-16, 
    5.116082e-16, 5.118331e-16, 5.108444e-16, 5.107839e-16, 5.098779e-16, 
    5.106843e-16, 5.110274e-16, 5.118989e-16, 5.124139e-16, 5.129034e-16, 
    5.139793e-16, 5.151798e-16, 5.168576e-16, 5.180622e-16, 5.188691e-16, 
    5.183745e-16, 5.188112e-16, 5.18323e-16, 5.180942e-16, 5.206341e-16, 
    5.192083e-16, 5.213476e-16, 5.212293e-16, 5.202613e-16, 5.212426e-16, 
    5.116421e-16, 5.113645e-16, 5.103998e-16, 5.111548e-16, 5.097792e-16, 
    5.105491e-16, 5.109915e-16, 5.126986e-16, 5.130738e-16, 5.134212e-16, 
    5.141074e-16, 5.149876e-16, 5.165303e-16, 5.178717e-16, 5.190956e-16, 
    5.19006e-16, 5.190375e-16, 5.193107e-16, 5.186338e-16, 5.194218e-16, 
    5.195538e-16, 5.192083e-16, 5.212135e-16, 5.206409e-16, 5.212268e-16, 
    5.208541e-16, 5.114548e-16, 5.119219e-16, 5.116695e-16, 5.121441e-16, 
    5.118096e-16, 5.132959e-16, 5.137413e-16, 5.158243e-16, 5.149701e-16, 
    5.163298e-16, 5.151084e-16, 5.153248e-16, 5.163734e-16, 5.151745e-16, 
    5.177974e-16, 5.16019e-16, 5.193212e-16, 5.175462e-16, 5.194324e-16, 
    5.190903e-16, 5.196568e-16, 5.201638e-16, 5.208018e-16, 5.219777e-16, 
    5.217055e-16, 5.226887e-16, 5.126183e-16, 5.132237e-16, 5.131707e-16, 
    5.138042e-16, 5.142725e-16, 5.152876e-16, 5.169139e-16, 5.163026e-16, 
    5.174251e-16, 5.176502e-16, 5.159451e-16, 5.169919e-16, 5.136289e-16, 
    5.141723e-16, 5.13849e-16, 5.126659e-16, 5.164431e-16, 5.145054e-16, 
    5.18082e-16, 5.170337e-16, 5.200915e-16, 5.185712e-16, 5.215557e-16, 
    5.228289e-16, 5.240278e-16, 5.254259e-16, 5.135543e-16, 5.13143e-16, 
    5.138796e-16, 5.148977e-16, 5.158426e-16, 5.170976e-16, 5.172262e-16, 
    5.17461e-16, 5.180697e-16, 5.185812e-16, 5.17535e-16, 5.187094e-16, 
    5.142977e-16, 5.166113e-16, 5.129872e-16, 5.140789e-16, 5.148378e-16, 
    5.145052e-16, 5.162329e-16, 5.166396e-16, 5.182917e-16, 5.174381e-16, 
    5.225145e-16, 5.202705e-16, 5.264906e-16, 5.247548e-16, 5.129993e-16, 
    5.13553e-16, 5.154786e-16, 5.145627e-16, 5.171815e-16, 5.178254e-16, 
    5.183489e-16, 5.190173e-16, 5.190897e-16, 5.194856e-16, 5.188367e-16, 
    5.194602e-16, 5.171003e-16, 5.181553e-16, 5.15259e-16, 5.159642e-16, 
    5.156399e-16, 5.152839e-16, 5.163824e-16, 5.175514e-16, 5.175769e-16, 
    5.179514e-16, 5.190056e-16, 5.171921e-16, 5.228029e-16, 5.193392e-16, 
    5.141567e-16, 5.152218e-16, 5.153745e-16, 5.149619e-16, 5.177608e-16, 
    5.167472e-16, 5.19476e-16, 5.187391e-16, 5.199466e-16, 5.193466e-16, 
    5.192583e-16, 5.184875e-16, 5.180073e-16, 5.167935e-16, 5.158055e-16, 
    5.150219e-16, 5.152041e-16, 5.160648e-16, 5.17623e-16, 5.19096e-16, 
    5.187734e-16, 5.198548e-16, 5.169917e-16, 5.181926e-16, 5.177284e-16, 
    5.189387e-16, 5.162863e-16, 5.185436e-16, 5.157086e-16, 5.159575e-16, 
    5.16727e-16, 5.182737e-16, 5.186165e-16, 5.189814e-16, 5.187564e-16, 
    5.176626e-16, 5.174836e-16, 5.167085e-16, 5.164941e-16, 5.159034e-16, 
    5.154138e-16, 5.15861e-16, 5.163303e-16, 5.176633e-16, 5.188634e-16, 
    5.20171e-16, 5.20491e-16, 5.220159e-16, 5.20774e-16, 5.228221e-16, 
    5.210799e-16, 5.24095e-16, 5.186751e-16, 5.210297e-16, 5.167622e-16, 
    5.172226e-16, 5.180545e-16, 5.199619e-16, 5.18933e-16, 5.201365e-16, 
    5.174766e-16, 5.160943e-16, 5.157371e-16, 5.150694e-16, 5.157523e-16, 
    5.156968e-16, 5.163501e-16, 5.161402e-16, 5.177075e-16, 5.168659e-16, 
    5.19256e-16, 5.201271e-16, 5.225856e-16, 5.240904e-16, 5.256215e-16, 
    5.262966e-16, 5.265021e-16, 5.26588e-16 ;

 CWDC_TO_LITR3C =
  1.610496e-16, 1.614913e-16, 1.614055e-16, 1.617615e-16, 1.615641e-16, 
    1.617972e-16, 1.611393e-16, 1.615088e-16, 1.61273e-16, 1.610895e-16, 
    1.624516e-16, 1.617774e-16, 1.631516e-16, 1.627222e-16, 1.638005e-16, 
    1.630847e-16, 1.639447e-16, 1.6378e-16, 1.64276e-16, 1.64134e-16, 
    1.647675e-16, 1.643415e-16, 1.650958e-16, 1.646659e-16, 1.647331e-16, 
    1.643274e-16, 1.619133e-16, 1.623676e-16, 1.618863e-16, 1.619512e-16, 
    1.619221e-16, 1.615682e-16, 1.613896e-16, 1.61016e-16, 1.610838e-16, 
    1.613583e-16, 1.619803e-16, 1.617694e-16, 1.623012e-16, 1.622892e-16, 
    1.628806e-16, 1.62614e-16, 1.636072e-16, 1.633251e-16, 1.641399e-16, 
    1.639351e-16, 1.641302e-16, 1.640711e-16, 1.64131e-16, 1.638306e-16, 
    1.639593e-16, 1.63695e-16, 1.626639e-16, 1.629671e-16, 1.620623e-16, 
    1.615173e-16, 1.611555e-16, 1.608984e-16, 1.609348e-16, 1.61004e-16, 
    1.613599e-16, 1.616945e-16, 1.619493e-16, 1.621196e-16, 1.622874e-16, 
    1.627947e-16, 1.630633e-16, 1.636641e-16, 1.635559e-16, 1.637393e-16, 
    1.639147e-16, 1.642089e-16, 1.641605e-16, 1.6429e-16, 1.637346e-16, 
    1.641037e-16, 1.634942e-16, 1.63661e-16, 1.623325e-16, 1.618263e-16, 
    1.616105e-16, 1.61422e-16, 1.609627e-16, 1.612799e-16, 1.611549e-16, 
    1.614524e-16, 1.616413e-16, 1.615479e-16, 1.621243e-16, 1.619002e-16, 
    1.630793e-16, 1.625717e-16, 1.638943e-16, 1.635781e-16, 1.6397e-16, 
    1.637701e-16, 1.641126e-16, 1.638044e-16, 1.643382e-16, 1.644543e-16, 
    1.64375e-16, 1.646799e-16, 1.637873e-16, 1.641302e-16, 1.615453e-16, 
    1.615605e-16, 1.616315e-16, 1.613193e-16, 1.613002e-16, 1.610141e-16, 
    1.612687e-16, 1.613771e-16, 1.616523e-16, 1.618149e-16, 1.619695e-16, 
    1.623092e-16, 1.626883e-16, 1.632182e-16, 1.635986e-16, 1.638534e-16, 
    1.636972e-16, 1.638351e-16, 1.636809e-16, 1.636087e-16, 1.644108e-16, 
    1.639605e-16, 1.646361e-16, 1.645987e-16, 1.64293e-16, 1.646029e-16, 
    1.615712e-16, 1.614835e-16, 1.611789e-16, 1.614173e-16, 1.609829e-16, 
    1.61226e-16, 1.613657e-16, 1.619048e-16, 1.620233e-16, 1.62133e-16, 
    1.623497e-16, 1.626276e-16, 1.631148e-16, 1.635384e-16, 1.639249e-16, 
    1.638966e-16, 1.639066e-16, 1.639928e-16, 1.637791e-16, 1.640279e-16, 
    1.640696e-16, 1.639605e-16, 1.645937e-16, 1.644129e-16, 1.645979e-16, 
    1.644802e-16, 1.61512e-16, 1.616596e-16, 1.615798e-16, 1.617297e-16, 
    1.616241e-16, 1.620934e-16, 1.622341e-16, 1.628919e-16, 1.626221e-16, 
    1.630515e-16, 1.626658e-16, 1.627342e-16, 1.630653e-16, 1.626867e-16, 
    1.63515e-16, 1.629534e-16, 1.639962e-16, 1.634356e-16, 1.640313e-16, 
    1.639233e-16, 1.641022e-16, 1.642623e-16, 1.644637e-16, 1.648351e-16, 
    1.647491e-16, 1.650596e-16, 1.618795e-16, 1.620706e-16, 1.620539e-16, 
    1.62254e-16, 1.624019e-16, 1.627224e-16, 1.63236e-16, 1.630429e-16, 
    1.633974e-16, 1.634685e-16, 1.6293e-16, 1.632606e-16, 1.621986e-16, 
    1.623702e-16, 1.622681e-16, 1.618945e-16, 1.630873e-16, 1.624754e-16, 
    1.636049e-16, 1.632738e-16, 1.642394e-16, 1.637593e-16, 1.647018e-16, 
    1.651039e-16, 1.654825e-16, 1.65924e-16, 1.62175e-16, 1.620452e-16, 
    1.622778e-16, 1.625993e-16, 1.628977e-16, 1.63294e-16, 1.633346e-16, 
    1.634087e-16, 1.63601e-16, 1.637625e-16, 1.634321e-16, 1.63803e-16, 
    1.624098e-16, 1.631404e-16, 1.61996e-16, 1.623407e-16, 1.625804e-16, 
    1.624753e-16, 1.630209e-16, 1.631494e-16, 1.636711e-16, 1.634015e-16, 
    1.650046e-16, 1.642959e-16, 1.662602e-16, 1.65712e-16, 1.619998e-16, 
    1.621746e-16, 1.627827e-16, 1.624935e-16, 1.633205e-16, 1.635238e-16, 
    1.636891e-16, 1.639002e-16, 1.639231e-16, 1.640481e-16, 1.638432e-16, 
    1.6404e-16, 1.632948e-16, 1.63628e-16, 1.627134e-16, 1.629361e-16, 
    1.628337e-16, 1.627212e-16, 1.630681e-16, 1.634373e-16, 1.634453e-16, 
    1.635636e-16, 1.638965e-16, 1.633238e-16, 1.650957e-16, 1.640019e-16, 
    1.623653e-16, 1.627016e-16, 1.627499e-16, 1.626196e-16, 1.635034e-16, 
    1.631833e-16, 1.640451e-16, 1.638123e-16, 1.641937e-16, 1.640042e-16, 
    1.639763e-16, 1.637329e-16, 1.635813e-16, 1.63198e-16, 1.628859e-16, 
    1.626385e-16, 1.62696e-16, 1.629678e-16, 1.634599e-16, 1.639251e-16, 
    1.638232e-16, 1.641647e-16, 1.632606e-16, 1.636398e-16, 1.634932e-16, 
    1.638754e-16, 1.630378e-16, 1.637506e-16, 1.628554e-16, 1.629339e-16, 
    1.63177e-16, 1.636654e-16, 1.637736e-16, 1.638889e-16, 1.638178e-16, 
    1.634724e-16, 1.634159e-16, 1.631711e-16, 1.631034e-16, 1.629168e-16, 
    1.627623e-16, 1.629035e-16, 1.630517e-16, 1.634726e-16, 1.638516e-16, 
    1.642645e-16, 1.643656e-16, 1.648471e-16, 1.644549e-16, 1.651017e-16, 
    1.645515e-16, 1.655037e-16, 1.637921e-16, 1.645357e-16, 1.631881e-16, 
    1.633335e-16, 1.635961e-16, 1.641985e-16, 1.638736e-16, 1.642536e-16, 
    1.634137e-16, 1.629771e-16, 1.628643e-16, 1.626535e-16, 1.628692e-16, 
    1.628516e-16, 1.630579e-16, 1.629917e-16, 1.634866e-16, 1.632208e-16, 
    1.639756e-16, 1.642507e-16, 1.65027e-16, 1.655022e-16, 1.659857e-16, 
    1.661989e-16, 1.662638e-16, 1.66291e-16 ;

 CWDC_vr =
  5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 
    5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110348e-05, 5.110348e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110346e-05, 5.110346e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 
    5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 
    5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 
    5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 
    5.110346e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110345e-05, 5.110347e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110347e-05, 
    5.110347e-05, 5.110347e-05, 5.110347e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110347e-05, 5.110347e-05, 
    5.110347e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110347e-05, 5.110346e-05, 5.110347e-05, 5.110347e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 5.110347e-05, 
    5.110347e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 
    5.110345e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110347e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110345e-05, 
    5.110345e-05, 5.110344e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110345e-05, 5.110346e-05, 5.110345e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 5.110346e-05, 
    5.110345e-05, 5.110345e-05, 5.110345e-05, 5.110344e-05, 5.110344e-05, 
    5.110344e-05, 5.110344e-05, 5.110344e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 CWDN =
  1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 
    1.789931e-09, 1.789932e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789932e-09, 1.789931e-09, 1.789932e-09, 1.789932e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 
    1.789932e-09, 1.789931e-09, 1.789932e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789932e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789931e-09, 1.789932e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789932e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 
    1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 1.789932e-09, 
    1.789932e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789932e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789932e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.78993e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 
    1.789931e-09, 1.789931e-09, 1.789931e-09, 1.789931e-09, 1.78993e-09, 
    1.78993e-09, 1.78993e-09, 1.78993e-09 ;

 CWDN_TO_LITR2N =
  1.019981e-18, 1.022779e-18, 1.022235e-18, 1.02449e-18, 1.02324e-18, 
    1.024715e-18, 1.020549e-18, 1.022889e-18, 1.021395e-18, 1.020234e-18, 
    1.02886e-18, 1.02459e-18, 1.033294e-18, 1.030574e-18, 1.037403e-18, 
    1.03287e-18, 1.038317e-18, 1.037273e-18, 1.040415e-18, 1.039515e-18, 
    1.043527e-18, 1.04083e-18, 1.045607e-18, 1.042884e-18, 1.043309e-18, 
    1.04074e-18, 1.025451e-18, 1.028328e-18, 1.02528e-18, 1.025691e-18, 
    1.025507e-18, 1.023265e-18, 1.022134e-18, 1.019768e-18, 1.020198e-18, 
    1.021936e-18, 1.025875e-18, 1.024539e-18, 1.027907e-18, 1.027831e-18, 
    1.031577e-18, 1.029889e-18, 1.036179e-18, 1.034392e-18, 1.039553e-18, 
    1.038255e-18, 1.039492e-18, 1.039117e-18, 1.039496e-18, 1.037594e-18, 
    1.038409e-18, 1.036735e-18, 1.030205e-18, 1.032125e-18, 1.026395e-18, 
    1.022943e-18, 1.020651e-18, 1.019023e-18, 1.019254e-18, 1.019692e-18, 
    1.021946e-18, 1.024065e-18, 1.025679e-18, 1.026758e-18, 1.027821e-18, 
    1.031033e-18, 1.032734e-18, 1.036539e-18, 1.035854e-18, 1.037016e-18, 
    1.038126e-18, 1.039989e-18, 1.039683e-18, 1.040503e-18, 1.036986e-18, 
    1.039324e-18, 1.035463e-18, 1.036519e-18, 1.028106e-18, 1.0249e-18, 
    1.023533e-18, 1.022339e-18, 1.01943e-18, 1.021439e-18, 1.020648e-18, 
    1.022532e-18, 1.023728e-18, 1.023137e-18, 1.026787e-18, 1.025368e-18, 
    1.032835e-18, 1.029621e-18, 1.037997e-18, 1.035995e-18, 1.038477e-18, 
    1.037211e-18, 1.03938e-18, 1.037428e-18, 1.040809e-18, 1.041544e-18, 
    1.041042e-18, 1.042973e-18, 1.037319e-18, 1.039491e-18, 1.02312e-18, 
    1.023216e-18, 1.023666e-18, 1.021689e-18, 1.021568e-18, 1.019756e-18, 
    1.021369e-18, 1.022055e-18, 1.023798e-18, 1.024828e-18, 1.025807e-18, 
    1.027959e-18, 1.03036e-18, 1.033715e-18, 1.036124e-18, 1.037738e-18, 
    1.036749e-18, 1.037622e-18, 1.036646e-18, 1.036188e-18, 1.041268e-18, 
    1.038416e-18, 1.042695e-18, 1.042459e-18, 1.040523e-18, 1.042485e-18, 
    1.023284e-18, 1.022729e-18, 1.0208e-18, 1.02231e-18, 1.019558e-18, 
    1.021098e-18, 1.021983e-18, 1.025397e-18, 1.026148e-18, 1.026842e-18, 
    1.028215e-18, 1.029975e-18, 1.03306e-18, 1.035743e-18, 1.038191e-18, 
    1.038012e-18, 1.038075e-18, 1.038621e-18, 1.037268e-18, 1.038844e-18, 
    1.039108e-18, 1.038417e-18, 1.042427e-18, 1.041282e-18, 1.042454e-18, 
    1.041708e-18, 1.02291e-18, 1.023844e-18, 1.023339e-18, 1.024288e-18, 
    1.023619e-18, 1.026592e-18, 1.027483e-18, 1.031649e-18, 1.02994e-18, 
    1.03266e-18, 1.030217e-18, 1.03065e-18, 1.032747e-18, 1.030349e-18, 
    1.035595e-18, 1.032038e-18, 1.038643e-18, 1.035092e-18, 1.038865e-18, 
    1.038181e-18, 1.039314e-18, 1.040328e-18, 1.041604e-18, 1.043955e-18, 
    1.043411e-18, 1.045378e-18, 1.025237e-18, 1.026447e-18, 1.026341e-18, 
    1.027608e-18, 1.028545e-18, 1.030575e-18, 1.033828e-18, 1.032605e-18, 
    1.03485e-18, 1.0353e-18, 1.03189e-18, 1.033984e-18, 1.027258e-18, 
    1.028345e-18, 1.027698e-18, 1.025332e-18, 1.032886e-18, 1.029011e-18, 
    1.036164e-18, 1.034067e-18, 1.040183e-18, 1.037142e-18, 1.043111e-18, 
    1.045658e-18, 1.048056e-18, 1.050852e-18, 1.027109e-18, 1.026286e-18, 
    1.027759e-18, 1.029795e-18, 1.031685e-18, 1.034195e-18, 1.034452e-18, 
    1.034922e-18, 1.036139e-18, 1.037162e-18, 1.03507e-18, 1.037419e-18, 
    1.028595e-18, 1.033223e-18, 1.025974e-18, 1.028158e-18, 1.029676e-18, 
    1.029011e-18, 1.032466e-18, 1.033279e-18, 1.036583e-18, 1.034876e-18, 
    1.045029e-18, 1.040541e-18, 1.052981e-18, 1.049509e-18, 1.025998e-18, 
    1.027106e-18, 1.030957e-18, 1.029125e-18, 1.034363e-18, 1.035651e-18, 
    1.036698e-18, 1.038035e-18, 1.038179e-18, 1.038971e-18, 1.037673e-18, 
    1.03892e-18, 1.034201e-18, 1.036311e-18, 1.030518e-18, 1.031928e-18, 
    1.03128e-18, 1.030568e-18, 1.032765e-18, 1.035103e-18, 1.035154e-18, 
    1.035903e-18, 1.038011e-18, 1.034384e-18, 1.045606e-18, 1.038678e-18, 
    1.028313e-18, 1.030444e-18, 1.030749e-18, 1.029924e-18, 1.035522e-18, 
    1.033494e-18, 1.038952e-18, 1.037478e-18, 1.039893e-18, 1.038693e-18, 
    1.038517e-18, 1.036975e-18, 1.036015e-18, 1.033587e-18, 1.031611e-18, 
    1.030044e-18, 1.030408e-18, 1.03213e-18, 1.035246e-18, 1.038192e-18, 
    1.037547e-18, 1.03971e-18, 1.033984e-18, 1.036385e-18, 1.035457e-18, 
    1.037877e-18, 1.032573e-18, 1.037087e-18, 1.031417e-18, 1.031915e-18, 
    1.033454e-18, 1.036547e-18, 1.037233e-18, 1.037963e-18, 1.037513e-18, 
    1.035325e-18, 1.034967e-18, 1.033417e-18, 1.032988e-18, 1.031807e-18, 
    1.030828e-18, 1.031722e-18, 1.032661e-18, 1.035327e-18, 1.037727e-18, 
    1.040342e-18, 1.040982e-18, 1.044032e-18, 1.041548e-18, 1.045644e-18, 
    1.04216e-18, 1.04819e-18, 1.03735e-18, 1.042059e-18, 1.033524e-18, 
    1.034445e-18, 1.036109e-18, 1.039924e-18, 1.037866e-18, 1.040273e-18, 
    1.034953e-18, 1.032189e-18, 1.031474e-18, 1.030139e-18, 1.031505e-18, 
    1.031394e-18, 1.0327e-18, 1.03228e-18, 1.035415e-18, 1.033732e-18, 
    1.038512e-18, 1.040254e-18, 1.045171e-18, 1.048181e-18, 1.051243e-18, 
    1.052593e-18, 1.053004e-18, 1.053176e-18 ;

 CWDN_TO_LITR3N =
  3.220992e-19, 3.229827e-19, 3.228111e-19, 3.235231e-19, 3.231283e-19, 
    3.235943e-19, 3.222786e-19, 3.230176e-19, 3.225459e-19, 3.22179e-19, 
    3.249031e-19, 3.235549e-19, 3.263033e-19, 3.254444e-19, 3.27601e-19, 
    3.261695e-19, 3.278895e-19, 3.2756e-19, 3.28552e-19, 3.282679e-19, 
    3.295349e-19, 3.28683e-19, 3.301916e-19, 3.293317e-19, 3.294662e-19, 
    3.286549e-19, 3.238266e-19, 3.247352e-19, 3.237727e-19, 3.239023e-19, 
    3.238442e-19, 3.231363e-19, 3.227792e-19, 3.220319e-19, 3.221677e-19, 
    3.227167e-19, 3.239606e-19, 3.235387e-19, 3.246023e-19, 3.245784e-19, 
    3.257611e-19, 3.25228e-19, 3.272143e-19, 3.266502e-19, 3.282798e-19, 
    3.278701e-19, 3.282605e-19, 3.281422e-19, 3.28262e-19, 3.276612e-19, 
    3.279187e-19, 3.273899e-19, 3.253278e-19, 3.259342e-19, 3.241246e-19, 
    3.230346e-19, 3.223109e-19, 3.217969e-19, 3.218695e-19, 3.22008e-19, 
    3.227199e-19, 3.23389e-19, 3.238986e-19, 3.242393e-19, 3.245749e-19, 
    3.255894e-19, 3.261267e-19, 3.273282e-19, 3.271118e-19, 3.274786e-19, 
    3.278294e-19, 3.284177e-19, 3.283209e-19, 3.285799e-19, 3.274692e-19, 
    3.282074e-19, 3.269884e-19, 3.273219e-19, 3.246651e-19, 3.236526e-19, 
    3.232211e-19, 3.22844e-19, 3.219254e-19, 3.225598e-19, 3.223097e-19, 
    3.229048e-19, 3.232826e-19, 3.230958e-19, 3.242486e-19, 3.238005e-19, 
    3.261585e-19, 3.251435e-19, 3.277885e-19, 3.271562e-19, 3.2794e-19, 
    3.275402e-19, 3.282251e-19, 3.276087e-19, 3.286764e-19, 3.289086e-19, 
    3.2875e-19, 3.293598e-19, 3.275745e-19, 3.282604e-19, 3.230905e-19, 
    3.23121e-19, 3.23263e-19, 3.226385e-19, 3.226004e-19, 3.220282e-19, 
    3.225374e-19, 3.227542e-19, 3.233046e-19, 3.236298e-19, 3.23939e-19, 
    3.246185e-19, 3.253767e-19, 3.264364e-19, 3.271972e-19, 3.277068e-19, 
    3.273944e-19, 3.276702e-19, 3.273619e-19, 3.272173e-19, 3.288216e-19, 
    3.27921e-19, 3.292721e-19, 3.291975e-19, 3.285861e-19, 3.292059e-19, 
    3.231424e-19, 3.229671e-19, 3.223578e-19, 3.228346e-19, 3.219658e-19, 
    3.224521e-19, 3.227315e-19, 3.238096e-19, 3.240466e-19, 3.24266e-19, 
    3.246994e-19, 3.252553e-19, 3.262296e-19, 3.270769e-19, 3.278499e-19, 
    3.277933e-19, 3.278132e-19, 3.279857e-19, 3.275582e-19, 3.280559e-19, 
    3.281392e-19, 3.27921e-19, 3.291875e-19, 3.288258e-19, 3.291959e-19, 
    3.289604e-19, 3.230241e-19, 3.233191e-19, 3.231597e-19, 3.234594e-19, 
    3.232482e-19, 3.241869e-19, 3.244682e-19, 3.257837e-19, 3.252443e-19, 
    3.26103e-19, 3.253316e-19, 3.254683e-19, 3.261306e-19, 3.253734e-19, 
    3.2703e-19, 3.259067e-19, 3.279924e-19, 3.268713e-19, 3.280626e-19, 
    3.278465e-19, 3.282043e-19, 3.285245e-19, 3.289274e-19, 3.296701e-19, 
    3.294982e-19, 3.301192e-19, 3.237589e-19, 3.241412e-19, 3.241078e-19, 
    3.245079e-19, 3.248037e-19, 3.254448e-19, 3.26472e-19, 3.260859e-19, 
    3.267948e-19, 3.26937e-19, 3.2586e-19, 3.265212e-19, 3.243972e-19, 
    3.247404e-19, 3.245362e-19, 3.23789e-19, 3.261746e-19, 3.249508e-19, 
    3.272097e-19, 3.265476e-19, 3.284788e-19, 3.275186e-19, 3.294036e-19, 
    3.302077e-19, 3.309649e-19, 3.31848e-19, 3.243501e-19, 3.240903e-19, 
    3.245556e-19, 3.251985e-19, 3.257953e-19, 3.26588e-19, 3.266691e-19, 
    3.268175e-19, 3.272019e-19, 3.275249e-19, 3.268642e-19, 3.276059e-19, 
    3.248196e-19, 3.262808e-19, 3.239919e-19, 3.246814e-19, 3.251607e-19, 
    3.249507e-19, 3.260418e-19, 3.262987e-19, 3.273421e-19, 3.26803e-19, 
    3.300091e-19, 3.285919e-19, 3.325204e-19, 3.314241e-19, 3.239995e-19, 
    3.243493e-19, 3.255654e-19, 3.24987e-19, 3.26641e-19, 3.270476e-19, 
    3.273782e-19, 3.278004e-19, 3.278461e-19, 3.280962e-19, 3.276864e-19, 
    3.280801e-19, 3.265896e-19, 3.27256e-19, 3.254267e-19, 3.258721e-19, 
    3.256673e-19, 3.254425e-19, 3.261362e-19, 3.268746e-19, 3.268906e-19, 
    3.271272e-19, 3.27793e-19, 3.266477e-19, 3.301913e-19, 3.280037e-19, 
    3.247305e-19, 3.254033e-19, 3.254997e-19, 3.252391e-19, 3.270068e-19, 
    3.263666e-19, 3.280902e-19, 3.276247e-19, 3.283873e-19, 3.280084e-19, 
    3.279526e-19, 3.274658e-19, 3.271625e-19, 3.263959e-19, 3.257719e-19, 
    3.25277e-19, 3.253921e-19, 3.259357e-19, 3.269198e-19, 3.278501e-19, 
    3.276463e-19, 3.283294e-19, 3.265211e-19, 3.272796e-19, 3.269864e-19, 
    3.277507e-19, 3.260756e-19, 3.275012e-19, 3.257107e-19, 3.258679e-19, 
    3.263539e-19, 3.273307e-19, 3.275472e-19, 3.277778e-19, 3.276356e-19, 
    3.269448e-19, 3.268317e-19, 3.263422e-19, 3.262068e-19, 3.258337e-19, 
    3.255245e-19, 3.258069e-19, 3.261033e-19, 3.269452e-19, 3.277032e-19, 
    3.28529e-19, 3.287312e-19, 3.296942e-19, 3.289099e-19, 3.302034e-19, 
    3.291031e-19, 3.310074e-19, 3.275843e-19, 3.290714e-19, 3.263761e-19, 
    3.266669e-19, 3.271923e-19, 3.28397e-19, 3.277472e-19, 3.285073e-19, 
    3.268273e-19, 3.259543e-19, 3.257287e-19, 3.25307e-19, 3.257383e-19, 
    3.257033e-19, 3.261158e-19, 3.259833e-19, 3.269732e-19, 3.264416e-19, 
    3.279511e-19, 3.285014e-19, 3.30054e-19, 3.310044e-19, 3.319715e-19, 
    3.323979e-19, 3.325277e-19, 3.325819e-19 ;

 CWDN_vr =
  1.02207e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.02207e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.02207e-07, 1.02207e-07, 1.02207e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.02207e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.02207e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.02207e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 1.022069e-07, 
    1.022069e-07, 1.022069e-07, 1.022069e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADCROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DEADSTEMC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 DEADSTEMN =
  6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 6.149015e-05, 
    6.149015e-05, 6.149015e-05, 6.149015e-05 ;

 DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.605194e-45, 0, 4.551417e-42, 
    2.802597e-45, 1.913193e-41, 3.698027e-42, 4.768479e-40, 1.216804e-40, 
    4.618803e-38, 8.893803e-40, 8.562508e-37, 1.82806e-38, 3.377825e-38, 
    7.783162e-40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.403934e-43, 3.363116e-44, 1.288718e-40, 1.736209e-41, 1.174148e-40, 
    6.60418e-41, 1.182948e-40, 6.143292e-42, 2.207185e-41, 1.56525e-42, 0, 
    1.401298e-45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 
    1.146262e-42, 3.783506e-43, 2.455075e-42, 1.418815e-41, 2.508002e-40, 
    1.572887e-40, 5.453685e-40, 2.337366e-42, 9.083777e-41, 1.989844e-43, 
    1.108427e-42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.802597e-45, 0, 
    1.158313e-41, 4.750402e-43, 2.451432e-41, 3.343498e-42, 9.89597e-41, 
    4.718172e-42, 8.623619e-40, 2.577666e-39, 1.221582e-39, 2.076547e-38, 
    3.974082e-42, 1.174288e-40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.121039e-44, 5.857428e-43, 7.708543e-42, 1.600283e-42, 6.42075e-42, 
    1.356457e-42, 6.488012e-43, 1.713117e-39, 2.23367e-41, 1.389566e-38, 
    9.852799e-39, 5.616474e-40, 1.024267e-38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4.203895e-45, 3.152922e-43, 1.569594e-41, 1.185358e-41, 
    1.308673e-41, 3.069544e-41, 3.661593e-42, 4.331554e-41, 6.516038e-41, 
    2.232128e-41, 9.408437e-39, 1.745448e-39, 9.780899e-39, 3.279918e-39, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 0, 0, 2.802597e-45, 0, 
    2.480298e-43, 0, 3.1724e-41, 1.093013e-43, 4.476448e-41, 1.543811e-41, 
    8.93538e-41, 4.185454e-40, 2.811773e-39, 8.485865e-38, 3.902624e-38, 
    6.231172e-37, 0, 0, 0, 0, 0, 0, 1.261169e-44, 1.401298e-45, 7.286752e-44, 
    1.527415e-43, 0, 1.681558e-44, 0, 0, 0, 0, 2.802597e-45, 0, 6.249791e-43, 
    1.961818e-44, 3.363915e-40, 3.005785e-42, 2.536987e-38, 9.203849e-37, 
    2.340174e-35, 8.675964e-34, 0, 0, 0, 0, 0, 2.522337e-44, 3.783506e-44, 
    8.267661e-44, 5.997557e-43, 3.09687e-42, 1.050974e-43, 4.652311e-42, 0, 
    4.203895e-45, 0, 0, 0, 0, 1.401298e-45, 5.605194e-45, 1.228939e-42, 
    7.567012e-44, 3.850611e-37, 5.781982e-40, 1.20543e-32, 1.566253e-34, 0, 
    0, 0, 0, 3.222986e-44, 2.718519e-43, 1.474166e-42, 1.229499e-41, 
    1.541148e-41, 5.278831e-41, 6.960249e-42, 4.876519e-41, 2.522337e-44, 
    7.917336e-43, 0, 0, 0, 0, 2.802597e-45, 1.107026e-43, 1.205117e-43, 
    4.091792e-43, 1.193206e-41, 3.363116e-44, 8.600233e-37, 3.375868e-41, 0, 
    0, 0, 0, 2.200039e-43, 7.006492e-45, 5.123568e-41, 5.111937e-42, 
    2.165973e-40, 3.4315e-41, 2.608517e-41, 2.298129e-42, 4.904545e-43, 
    8.407791e-45, 0, 0, 0, 1.401298e-45, 1.401298e-43, 1.573378e-41, 
    5.706087e-42, 1.638048e-40, 1.681558e-44, 8.940284e-43, 1.975831e-43, 
    9.598894e-42, 1.401298e-45, 2.766163e-42, 0, 0, 7.006492e-45, 
    1.161676e-42, 3.465411e-42, 1.098618e-41, 5.399203e-42, 1.59748e-43, 
    8.82818e-44, 7.006492e-45, 2.802597e-45, 0, 0, 0, 1.401298e-45, 
    1.59748e-43, 7.578222e-42, 4.277912e-40, 1.117072e-39, 9.486179e-38, 
    2.598732e-39, 9.070593e-37, 6.421963e-39, 2.808711e-35, 4.191284e-42, 
    5.521899e-39, 8.407791e-45, 3.783506e-44, 5.717298e-43, 2.275709e-40, 
    9.427936e-42, 3.860339e-40, 8.68805e-44, 1.401298e-45, 0, 0, 0, 0, 
    1.401298e-45, 1.401298e-45, 1.849714e-43, 1.121039e-44, 2.590861e-41, 
    3.750631e-40, 4.682267e-37, 2.766208e-35, 1.414291e-33, 7.510774e-33, 
    1.238513e-32, 1.524886e-32 ;

 DISPVEGC =
  0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 0.1735653, 
    0.1735653, 0.1735653 ;

 DISPVEGN =
  0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997, 0.003631997, 0.003631997, 
    0.003631997, 0.003631997, 0.003631997 ;

 DSTDEP =
  2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 2.653438e-12, 
    2.653438e-12, 2.653438e-12, 2.653438e-12 ;

 DSTFLXT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_CONV_NFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD100N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10C_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_PROD10N_GAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDC_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_DEADSTEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 DWT_SEEDN_TO_LEAF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 EFLX_GRND_LAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 EFLX_LH_TOT =
  22.01506, 22.07914, 22.0667, 22.11838, 22.08974, 22.12356, 22.02809, 
    22.08165, 22.04748, 22.02089, 22.21867, 22.12069, 22.32102, 22.25834, 
    22.41604, 22.31121, 22.43722, 22.41311, 22.48593, 22.46507, 22.55809, 
    22.49556, 22.60652, 22.54321, 22.55307, 22.49348, 22.14049, 22.20643, 
    22.13656, 22.14597, 22.14177, 22.0903, 22.06432, 22.01023, 22.02006, 
    22.05983, 22.1502, 22.11957, 22.19697, 22.19522, 22.28147, 22.24257, 
    22.38778, 22.34649, 22.46594, 22.43586, 22.46451, 22.45584, 22.46462, 
    22.42053, 22.43941, 22.40065, 22.24983, 22.29409, 22.16215, 22.08282, 
    22.03042, 21.9932, 21.99846, 22.00847, 22.06006, 22.10869, 22.14574, 
    22.17053, 22.19497, 22.2688, 22.30812, 22.39608, 22.38028, 22.40711, 
    22.43288, 22.47605, 22.46895, 22.48796, 22.40646, 22.46058, 22.37126, 
    22.39567, 22.2013, 22.12784, 22.09637, 22.06908, 22.0025, 22.04845, 
    22.03032, 22.07353, 22.10095, 22.0874, 22.17121, 22.1386, 22.31045, 
    22.23636, 22.42987, 22.38353, 22.441, 22.41168, 22.46189, 22.4167, 
    22.49506, 22.5121, 22.50045, 22.54532, 22.41419, 22.46448, 22.08701, 
    22.08921, 22.09954, 22.05416, 22.0514, 22.00994, 22.04686, 22.06256, 
    22.10257, 22.12618, 22.14866, 22.19812, 22.25337, 22.33079, 22.38653, 
    22.4239, 22.401, 22.42121, 22.39861, 22.38803, 22.50569, 22.43957, 
    22.53886, 22.53338, 22.4884, 22.53399, 22.09077, 22.07805, 22.03383, 
    22.06844, 22.00544, 22.04065, 22.06089, 22.13921, 22.15651, 22.17245, 
    22.20403, 22.24456, 22.31569, 22.37769, 22.43439, 22.43024, 22.4317, 
    22.44434, 22.41299, 22.44949, 22.45559, 22.4396, 22.53264, 22.50605, 
    22.53326, 22.51595, 22.0822, 22.10361, 22.09203, 22.11379, 22.09844, 
    22.16664, 22.1871, 22.28306, 22.24374, 22.30642, 22.25013, 22.26008, 
    22.30833, 22.25319, 22.37421, 22.29202, 22.44483, 22.36253, 22.44998, 
    22.43414, 22.4604, 22.48389, 22.51352, 22.56812, 22.55548, 22.60122, 
    22.13558, 22.16335, 22.16096, 22.19008, 22.21162, 22.2584, 22.33343, 
    22.30522, 22.35708, 22.36747, 22.28873, 22.33701, 22.18199, 22.20694, 
    22.19213, 22.13773, 22.31164, 22.22228, 22.38744, 22.33897, 22.48053, 
    22.41003, 22.54851, 22.60764, 22.66362, 22.72877, 22.17858, 22.15969, 
    22.19356, 22.24035, 22.28397, 22.34191, 22.34788, 22.35872, 22.38689, 
    22.41056, 22.36209, 22.4165, 22.21261, 22.31943, 22.1525, 22.20263, 
    22.23762, 22.22233, 22.30201, 22.32079, 22.39711, 22.35768, 22.59299, 
    22.48877, 22.77861, 22.69745, 22.15308, 22.17854, 22.26715, 22.22499, 
    22.34582, 22.37557, 22.39981, 22.43073, 22.43411, 22.45244, 22.4224, 
    22.45127, 22.34204, 22.39084, 22.25709, 22.28958, 22.27465, 22.25824, 
    22.30891, 22.36284, 22.36409, 22.38137, 22.42994, 22.34631, 22.60628, 
    22.44543, 22.20631, 22.25528, 22.26239, 22.2434, 22.37258, 22.32573, 
    22.45201, 22.41787, 22.47383, 22.44601, 22.44191, 22.40622, 22.38399, 
    22.32786, 22.28225, 22.24616, 22.25456, 22.29421, 22.36616, 22.43437, 
    22.41941, 22.46958, 22.33704, 22.39253, 22.37105, 22.4271, 22.30445, 
    22.40859, 22.27782, 22.2893, 22.3248, 22.39623, 22.41219, 22.42906, 
    22.41867, 22.36801, 22.35975, 22.32396, 22.31403, 22.28681, 22.26423, 
    22.28483, 22.30646, 22.36807, 22.42359, 22.48421, 22.49909, 22.56977, 
    22.5121, 22.60715, 22.52612, 22.66655, 22.41477, 22.52394, 22.32645, 
    22.34772, 22.38611, 22.47445, 22.42684, 22.48256, 22.35944, 22.29553, 
    22.27913, 22.24834, 22.27983, 22.27728, 22.30742, 22.29774, 22.37012, 
    22.33123, 22.44179, 22.48215, 22.59639, 22.66646, 22.73801, 22.76957, 
    22.77918, 22.7832 ;

 EFLX_LH_TOT_R =
  22.01506, 22.07914, 22.0667, 22.11838, 22.08974, 22.12356, 22.02809, 
    22.08165, 22.04748, 22.02089, 22.21867, 22.12069, 22.32102, 22.25834, 
    22.41604, 22.31121, 22.43722, 22.41311, 22.48593, 22.46507, 22.55809, 
    22.49556, 22.60652, 22.54321, 22.55307, 22.49348, 22.14049, 22.20643, 
    22.13656, 22.14597, 22.14177, 22.0903, 22.06432, 22.01023, 22.02006, 
    22.05983, 22.1502, 22.11957, 22.19697, 22.19522, 22.28147, 22.24257, 
    22.38778, 22.34649, 22.46594, 22.43586, 22.46451, 22.45584, 22.46462, 
    22.42053, 22.43941, 22.40065, 22.24983, 22.29409, 22.16215, 22.08282, 
    22.03042, 21.9932, 21.99846, 22.00847, 22.06006, 22.10869, 22.14574, 
    22.17053, 22.19497, 22.2688, 22.30812, 22.39608, 22.38028, 22.40711, 
    22.43288, 22.47605, 22.46895, 22.48796, 22.40646, 22.46058, 22.37126, 
    22.39567, 22.2013, 22.12784, 22.09637, 22.06908, 22.0025, 22.04845, 
    22.03032, 22.07353, 22.10095, 22.0874, 22.17121, 22.1386, 22.31045, 
    22.23636, 22.42987, 22.38353, 22.441, 22.41168, 22.46189, 22.4167, 
    22.49506, 22.5121, 22.50045, 22.54532, 22.41419, 22.46448, 22.08701, 
    22.08921, 22.09954, 22.05416, 22.0514, 22.00994, 22.04686, 22.06256, 
    22.10257, 22.12618, 22.14866, 22.19812, 22.25337, 22.33079, 22.38653, 
    22.4239, 22.401, 22.42121, 22.39861, 22.38803, 22.50569, 22.43957, 
    22.53886, 22.53338, 22.4884, 22.53399, 22.09077, 22.07805, 22.03383, 
    22.06844, 22.00544, 22.04065, 22.06089, 22.13921, 22.15651, 22.17245, 
    22.20403, 22.24456, 22.31569, 22.37769, 22.43439, 22.43024, 22.4317, 
    22.44434, 22.41299, 22.44949, 22.45559, 22.4396, 22.53264, 22.50605, 
    22.53326, 22.51595, 22.0822, 22.10361, 22.09203, 22.11379, 22.09844, 
    22.16664, 22.1871, 22.28306, 22.24374, 22.30642, 22.25013, 22.26008, 
    22.30833, 22.25319, 22.37421, 22.29202, 22.44483, 22.36253, 22.44998, 
    22.43414, 22.4604, 22.48389, 22.51352, 22.56812, 22.55548, 22.60122, 
    22.13558, 22.16335, 22.16096, 22.19008, 22.21162, 22.2584, 22.33343, 
    22.30522, 22.35708, 22.36747, 22.28873, 22.33701, 22.18199, 22.20694, 
    22.19213, 22.13773, 22.31164, 22.22228, 22.38744, 22.33897, 22.48053, 
    22.41003, 22.54851, 22.60764, 22.66362, 22.72877, 22.17858, 22.15969, 
    22.19356, 22.24035, 22.28397, 22.34191, 22.34788, 22.35872, 22.38689, 
    22.41056, 22.36209, 22.4165, 22.21261, 22.31943, 22.1525, 22.20263, 
    22.23762, 22.22233, 22.30201, 22.32079, 22.39711, 22.35768, 22.59299, 
    22.48877, 22.77861, 22.69745, 22.15308, 22.17854, 22.26715, 22.22499, 
    22.34582, 22.37557, 22.39981, 22.43073, 22.43411, 22.45244, 22.4224, 
    22.45127, 22.34204, 22.39084, 22.25709, 22.28958, 22.27465, 22.25824, 
    22.30891, 22.36284, 22.36409, 22.38137, 22.42994, 22.34631, 22.60628, 
    22.44543, 22.20631, 22.25528, 22.26239, 22.2434, 22.37258, 22.32573, 
    22.45201, 22.41787, 22.47383, 22.44601, 22.44191, 22.40622, 22.38399, 
    22.32786, 22.28225, 22.24616, 22.25456, 22.29421, 22.36616, 22.43437, 
    22.41941, 22.46958, 22.33704, 22.39253, 22.37105, 22.4271, 22.30445, 
    22.40859, 22.27782, 22.2893, 22.3248, 22.39623, 22.41219, 22.42906, 
    22.41867, 22.36801, 22.35975, 22.32396, 22.31403, 22.28681, 22.26423, 
    22.28483, 22.30646, 22.36807, 22.42359, 22.48421, 22.49909, 22.56977, 
    22.5121, 22.60715, 22.52612, 22.66655, 22.41477, 22.52394, 22.32645, 
    22.34772, 22.38611, 22.47445, 22.42684, 22.48256, 22.35944, 22.29553, 
    22.27913, 22.24834, 22.27983, 22.27728, 22.30742, 22.29774, 22.37012, 
    22.33123, 22.44179, 22.48215, 22.59639, 22.66646, 22.73801, 22.76957, 
    22.77918, 22.7832 ;

 EFLX_LH_TOT_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 ELAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 ER =
  6.191209e-08, 6.218511e-08, 6.213204e-08, 6.235225e-08, 6.22301e-08, 
    6.237429e-08, 6.196745e-08, 6.219594e-08, 6.205008e-08, 6.193667e-08, 
    6.277961e-08, 6.236208e-08, 6.321343e-08, 6.29471e-08, 6.361618e-08, 
    6.317198e-08, 6.370576e-08, 6.360339e-08, 6.391155e-08, 6.382326e-08, 
    6.421742e-08, 6.39523e-08, 6.442178e-08, 6.415411e-08, 6.419598e-08, 
    6.394355e-08, 6.244612e-08, 6.272763e-08, 6.242944e-08, 6.246958e-08, 
    6.245157e-08, 6.223262e-08, 6.212228e-08, 6.189123e-08, 6.193318e-08, 
    6.210288e-08, 6.248763e-08, 6.235703e-08, 6.26862e-08, 6.267877e-08, 
    6.304526e-08, 6.288002e-08, 6.349605e-08, 6.332096e-08, 6.382695e-08, 
    6.369969e-08, 6.382097e-08, 6.37842e-08, 6.382145e-08, 6.363481e-08, 
    6.371478e-08, 6.355055e-08, 6.291096e-08, 6.309892e-08, 6.253835e-08, 
    6.220129e-08, 6.197747e-08, 6.181863e-08, 6.184109e-08, 6.188389e-08, 
    6.210387e-08, 6.231072e-08, 6.246836e-08, 6.25738e-08, 6.267771e-08, 
    6.299219e-08, 6.315867e-08, 6.353144e-08, 6.346419e-08, 6.357814e-08, 
    6.368703e-08, 6.386984e-08, 6.383975e-08, 6.392029e-08, 6.357515e-08, 
    6.380452e-08, 6.342587e-08, 6.352943e-08, 6.27059e-08, 6.239227e-08, 
    6.225892e-08, 6.214224e-08, 6.185834e-08, 6.205439e-08, 6.19771e-08, 
    6.216099e-08, 6.227782e-08, 6.222004e-08, 6.257669e-08, 6.243803e-08, 
    6.316854e-08, 6.285387e-08, 6.367434e-08, 6.347799e-08, 6.372139e-08, 
    6.359719e-08, 6.381001e-08, 6.361848e-08, 6.395027e-08, 6.402251e-08, 
    6.397314e-08, 6.41628e-08, 6.360786e-08, 6.382096e-08, 6.221842e-08, 
    6.222784e-08, 6.227175e-08, 6.207874e-08, 6.206693e-08, 6.189008e-08, 
    6.204745e-08, 6.211446e-08, 6.22846e-08, 6.238523e-08, 6.248089e-08, 
    6.269123e-08, 6.292615e-08, 6.325467e-08, 6.349072e-08, 6.364895e-08, 
    6.355192e-08, 6.363758e-08, 6.354183e-08, 6.349695e-08, 6.399544e-08, 
    6.371552e-08, 6.413553e-08, 6.411229e-08, 6.39222e-08, 6.411491e-08, 
    6.223446e-08, 6.218023e-08, 6.199193e-08, 6.213929e-08, 6.187082e-08, 
    6.202109e-08, 6.210749e-08, 6.244091e-08, 6.251418e-08, 6.258211e-08, 
    6.271628e-08, 6.288847e-08, 6.319055e-08, 6.34534e-08, 6.369337e-08, 
    6.367579e-08, 6.368198e-08, 6.373558e-08, 6.36028e-08, 6.375738e-08, 
    6.378333e-08, 6.371549e-08, 6.410917e-08, 6.39967e-08, 6.411179e-08, 
    6.403856e-08, 6.219786e-08, 6.228911e-08, 6.22398e-08, 6.233252e-08, 
    6.22672e-08, 6.255767e-08, 6.264477e-08, 6.305234e-08, 6.288508e-08, 
    6.315129e-08, 6.291213e-08, 6.29545e-08, 6.315996e-08, 6.292505e-08, 
    6.34389e-08, 6.30905e-08, 6.373767e-08, 6.338972e-08, 6.375947e-08, 
    6.369233e-08, 6.38035e-08, 6.390305e-08, 6.402831e-08, 6.425942e-08, 
    6.420591e-08, 6.43992e-08, 6.242516e-08, 6.254352e-08, 6.25331e-08, 
    6.265698e-08, 6.27486e-08, 6.294718e-08, 6.326568e-08, 6.314591e-08, 
    6.33658e-08, 6.340995e-08, 6.307588e-08, 6.328098e-08, 6.262274e-08, 
    6.272907e-08, 6.266577e-08, 6.243449e-08, 6.317349e-08, 6.279422e-08, 
    6.349462e-08, 6.328914e-08, 6.388886e-08, 6.359058e-08, 6.417645e-08, 
    6.442689e-08, 6.466265e-08, 6.493813e-08, 6.260812e-08, 6.25277e-08, 
    6.267172e-08, 6.287096e-08, 6.305586e-08, 6.330166e-08, 6.332682e-08, 
    6.337287e-08, 6.349217e-08, 6.359246e-08, 6.338743e-08, 6.361761e-08, 
    6.275372e-08, 6.320642e-08, 6.249729e-08, 6.27108e-08, 6.285921e-08, 
    6.279412e-08, 6.313223e-08, 6.321191e-08, 6.353574e-08, 6.336835e-08, 
    6.436507e-08, 6.392407e-08, 6.514793e-08, 6.480587e-08, 6.249959e-08, 
    6.260785e-08, 6.298463e-08, 6.280536e-08, 6.331808e-08, 6.344429e-08, 
    6.35469e-08, 6.367805e-08, 6.369222e-08, 6.376993e-08, 6.364259e-08, 
    6.376491e-08, 6.330219e-08, 6.350896e-08, 6.294157e-08, 6.307966e-08, 
    6.301614e-08, 6.294646e-08, 6.316152e-08, 6.339064e-08, 6.339556e-08, 
    6.346902e-08, 6.367603e-08, 6.332016e-08, 6.442196e-08, 6.374147e-08, 
    6.27259e-08, 6.293441e-08, 6.296421e-08, 6.288344e-08, 6.343164e-08, 
    6.3233e-08, 6.376804e-08, 6.362344e-08, 6.386038e-08, 6.374263e-08, 
    6.372531e-08, 6.357409e-08, 6.347994e-08, 6.32421e-08, 6.304859e-08, 
    6.289515e-08, 6.293084e-08, 6.309938e-08, 6.340467e-08, 6.36935e-08, 
    6.363022e-08, 6.384236e-08, 6.32809e-08, 6.351632e-08, 6.342533e-08, 
    6.36626e-08, 6.314273e-08, 6.358538e-08, 6.302958e-08, 6.307831e-08, 
    6.322905e-08, 6.353228e-08, 6.359939e-08, 6.367102e-08, 6.362682e-08, 
    6.341242e-08, 6.33773e-08, 6.322539e-08, 6.318344e-08, 6.30677e-08, 
    6.297188e-08, 6.305942e-08, 6.315137e-08, 6.341251e-08, 6.364786e-08, 
    6.390447e-08, 6.396727e-08, 6.426707e-08, 6.4023e-08, 6.442575e-08, 
    6.40833e-08, 6.467612e-08, 6.361105e-08, 6.407326e-08, 6.323592e-08, 
    6.332613e-08, 6.348927e-08, 6.386351e-08, 6.366148e-08, 6.389776e-08, 
    6.337593e-08, 6.310519e-08, 6.303516e-08, 6.290448e-08, 6.303815e-08, 
    6.302728e-08, 6.315518e-08, 6.311409e-08, 6.342119e-08, 6.325622e-08, 
    6.372487e-08, 6.38959e-08, 6.437893e-08, 6.467506e-08, 6.497654e-08, 
    6.510964e-08, 6.515015e-08, 6.516709e-08 ;

 ERRH2O =
  -22914.72, -22949.22, -22942.46, -22970.67, -22954.97, -22973.52, 
    -22921.65, -22950.6, -22932.06, -22917.79, -23026.66, -22971.94, 
    -23085.22, -23049.03, -23140.62, -23079.54, -23153.16, -23138.82, 
    -23182.37, -23169.77, -23226.81, -23188.21, -23257.21, -23217.5, 
    -23223.65, -23186.96, -22982.84, -23019.78, -22980.67, -22985.89, 
    -22983.55, -22955.29, -22941.22, -22912.11, -22917.35, -22938.75, 
    -22988.25, -22971.29, -23014.3, -23013.32, -23062.28, -23040.03, 
    -23123.93, -23099.93, -23170.29, -23152.3, -23169.44, -23164.23, 
    -23169.51, -23143.21, -23154.43, -23131.48, -23044.17, -23069.57, 
    -22994.88, -22951.29, -22922.91, -22903.05, -22905.85, -22911.19, 
    -22938.88, -22965.31, -22985.73, -22999.53, -23013.18, -23055.11, 
    -23077.72, -23128.83, -23119.54, -23135.31, -23150.53, -23176.4, 
    -23172.11, -23183.62, -23134.89, -23167.11, -23114.27, -23128.55, 
    -23016.91, -22975.85, -22958.67, -22943.75, -22908, -22932.61, -22922.87, 
    -22946.14, -22961.08, -22953.68, -22999.91, -22981.79, -23079.07, 
    -23036.53, -23148.74, -23121.44, -23155.36, -23137.96, -23167.89, 
    -23140.93, -23187.92, -23198.34, -23191.21, -23218.77, -23139.45, 
    -23169.45, -22953.47, -22954.68, -22960.3, -22935.69, -22934.2, 
    -22911.96, -22931.73, -22940.22, -22961.95, -22974.93, -22987.37, 
    -23014.96, -23046.21, -23090.89, -23123.2, -23145.19, -23131.66, 
    -23143.6, -23130.26, -23124.05, -23194.43, -23154.53, -23214.78, 
    -23211.38, -23183.89, -23211.77, -22955.53, -22948.59, -22924.73, 
    -22943.38, -22909.56, -22928.41, -22939.34, -22982.16, -22991.71, 
    -23000.62, -23018.26, -23041.16, -23082.08, -23118.05, -23151.41, 
    -23148.95, -23149.81, -23157.36, -23138.74, -23160.43, -23164.11, 
    -23154.53, -23210.93, -23194.61, -23211.31, -23200.66, -22950.84, 
    -22962.54, -22956.21, -22968.12, -22959.72, -22997.42, -23008.86, 
    -23063.25, -23040.7, -23076.71, -23044.33, -23050.02, -23077.9, 
    -23046.06, -23116.06, -23068.43, -23157.65, -23109.33, -23160.73, 
    -23151.27, -23166.96, -23181.15, -23199.18, -23233, -23225.11, -23253.81, 
    -22980.11, -22995.56, -22994.19, -23010.45, -23022.54, -23049.03, 
    -23092.4, -23075.97, -23106.04, -23112.08, -23066.44, -23094.51, 
    -23005.96, -23019.96, -23011.61, -22981.33, -23079.74, -23028.59, 
    -23123.73, -23095.61, -23179.12, -23137.04, -23220.78, -23257.98, 
    -23293.79, -23336.3, -23004.04, -22993.48, -23012.39, -23038.82, 
    -23063.72, -23097.31, -23100.73, -23107.01, -23123.39, -23137.3, -23109, 
    -23140.8, -23023.23, -23084.25, -22989.51, -23017.55, -23037.25, 
    -23028.57, -23074.1, -23085, -23129.43, -23106.39, -23248.72, -23184.17, 
    -23369, -23315.91, -22989.81, -23004.01, -23054.08, -23030.07, -23099.54, 
    -23116.8, -23130.97, -23149.27, -23151.25, -23162.21, -23144.29, 
    -23161.5, -23097.38, -23125.71, -23048.28, -23066.95, -23058.33, 
    -23048.93, -23078.1, -23109.45, -23110.11, -23120.21, -23149.01, 
    -23099.82, -23257.26, -23158.21, -23019.54, -23047.32, -23051.33, 
    -23040.48, -23115.06, -23087.9, -23161.94, -23141.62, -23175.05, 
    -23158.35, -23155.91, -23134.74, -23121.71, -23089.15, -23062.73, 
    -23042.05, -23046.83, -23069.63, -23111.37, -23151.44, -23142.57, 
    -23172.48, -23094.49, -23126.74, -23114.2, -23147.1, -23075.54, 
    -23136.33, -23060.15, -23066.77, -23087.36, -23128.95, -23138.27, 
    -23148.28, -23142.09, -23112.43, -23107.62, -23086.85, -23081.1, 
    -23065.32, -23052.36, -23064.2, -23076.72, -23112.44, -23145.04, 
    -23181.35, -23190.37, -23234.15, -23198.42, -23257.83, -23207.19, 
    -23295.87, -23139.9, -23205.72, -23088.3, -23100.63, -23123, -23175.51, 
    -23146.94, -23180.4, -23107.43, -23070.42, -23060.91, -23043.3, 
    -23061.31, -23059.84, -23077.23, -23071.63, -23113.63, -23091.1, 
    -23155.85, -23180.13, -23250.78, -23295.7, -23342.25, -23362.99, 
    -23369.35, -23372.02 ;

 ERRH2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ERRSEB =
  -3.69623e-15, -1.825747e-14, -1.721879e-14, -7.622824e-16, -1.55312e-14, 
    -1.452947e-14, -1.036944e-14, -1.0717e-14, -8.234834e-15, -6.096844e-15, 
    -1.71979e-14, -1.147303e-14, -1.520852e-14, -8.090092e-15, -8.807115e-15, 
    -1.425185e-14, -1.411845e-14, -1.010249e-14, -1.016985e-14, 
    -1.476563e-14, -1.370004e-14, -1.386352e-14, -9.035011e-15, 
    -1.280079e-14, -1.486754e-14, -1.847101e-14, -4.051385e-15, 
    -1.397247e-14, -1.379838e-14, -7.17749e-15, -1.876687e-14, -1.556624e-14, 
    -1.065504e-14, -1.406412e-14, -1.367741e-14, -2.661137e-14, 
    -4.045202e-15, -1.141416e-14, -9.542579e-15, -1.043118e-14, 
    -1.526382e-14, -1.709295e-14, -1.444489e-14, -1.046805e-14, 
    -1.274266e-14, -1.081076e-14, -1.020118e-14, -1.191644e-14, -9.57687e-15, 
    -1.480755e-14, -8.995957e-15, -1.798401e-14, -1.166187e-14, 
    -3.955393e-15, -1.274391e-14, -1.716705e-14, -1.274966e-14, 
    -1.919981e-14, -1.568019e-14, -1.432844e-14, -1.362768e-14, 
    -1.683234e-14, -1.641454e-14, -9.907561e-15, -2.153159e-14, 
    -8.326927e-15, -1.286919e-14, -9.412899e-15, -1.085405e-14, -1.57262e-14, 
    -1.344885e-14, -1.277875e-14, -1.547907e-14, -9.929894e-15, 
    -1.805241e-14, -1.052545e-14, -1.121561e-14, -1.701246e-14, 
    -9.819214e-15, -2.053319e-14, -8.921068e-15, -1.440345e-14, 
    -1.336695e-14, -1.104143e-14, -1.674323e-14, -7.633535e-15, 
    -1.752675e-14, -1.760593e-14, -1.240587e-14, -1.180665e-14, 
    -1.358607e-14, -9.015188e-15, -6.530687e-15, -9.860106e-15, 
    -1.704353e-14, -1.664606e-14, -6.896837e-15, -9.780361e-15, 
    -9.733629e-15, -1.770362e-14, -1.836367e-14, -9.245e-15, -1.181823e-14, 
    -8.663179e-15, -1.352073e-14, -1.238647e-14, -1.380019e-14, 
    -1.401537e-14, -1.785767e-14, -9.979645e-15, -1.339391e-14, 
    -8.359703e-15, -4.465242e-15, -1.677656e-14, -5.957505e-15, 
    -1.144583e-14, -6.895012e-15, -1.427644e-14, -1.128186e-14, 
    -1.673588e-14, -1.796106e-14, -1.040077e-14, -1.878576e-14, 
    -1.549168e-14, -9.482453e-15, -7.845855e-15, -4.620991e-15, 
    -1.512153e-14, -1.272148e-14, -9.655602e-15, -1.113067e-14, 
    -2.314057e-14, -1.115813e-14, -1.424841e-14, -1.314417e-14, 
    -8.625826e-15, -1.77725e-14, -7.33242e-15, -1.667812e-14, -1.365832e-14, 
    -1.434651e-14, -1.446715e-14, -1.504208e-14, -7.945884e-15, 
    -1.761263e-14, -1.636425e-14, -1.000198e-14, -1.600193e-14, 
    -7.196956e-15, -1.610871e-14, -1.291347e-14, -1.504552e-14, 
    -2.063049e-14, -1.218103e-14, -1.649066e-14, -1.347743e-14, -4.34998e-15, 
    -1.342924e-14, -1.190755e-14, -1.735072e-14, -9.623951e-15, 
    -1.139567e-14, -2.032091e-14, -1.44174e-14, -2.048e-14, -1.153205e-14, 
    -1.185282e-14, -4.837422e-15, -2.090579e-14, -8.189484e-15, 
    -1.777406e-14, -8.148349e-15, -1.411741e-14, -1.094856e-14, 
    -1.044494e-14, -1.250438e-14, -7.555389e-15, -3.961245e-15, 
    -2.326999e-14, -1.389602e-14, -1.629071e-14, -1.347704e-14, 
    -2.053143e-14, -1.447479e-14, -9.98056e-15, -1.791968e-14, -1.6565e-14, 
    -1.749311e-14, -1.388391e-14, -1.030316e-14, -1.348947e-14, 
    -1.334491e-14, -2.019836e-14, -1.489847e-14, -2.014948e-14, 
    -1.927088e-14, -1.282554e-14, -1.127396e-14, -1.179896e-14, 
    -1.266552e-14, -1.321973e-14, -2.20493e-14, -8.092408e-15, -8.070557e-15, 
    -1.140537e-14, -7.218851e-15, -1.521204e-14, -2.279371e-14, 
    -1.590301e-14, -1.330593e-14, -1.393993e-14, -1.204009e-14, 
    -6.995837e-15, -1.933286e-14, -6.457949e-15, -6.870978e-15, 
    -1.346024e-14, -1.397426e-14, -1.12293e-14, -1.409705e-14, -1.126178e-14, 
    -1.075268e-14, -1.354274e-14, -1.892903e-14, -1.520079e-14, 
    -1.701361e-14, -1.023798e-14, -1.356102e-14, -1.211717e-14, 
    -2.062239e-14, -8.996677e-15, -1.695179e-14, -2.001127e-14, 
    -1.350331e-14, -8.978899e-15, -1.636707e-14, -9.551864e-15, -1.85274e-14, 
    -9.758201e-15, -7.751616e-15, -1.991044e-14, -1.030175e-14, -3.2275e-15, 
    -2.075219e-14, -1.719797e-14, -6.762134e-15, -1.189739e-14, 
    -1.706374e-14, -1.344383e-14, -1.965388e-14, -9.215571e-15, 
    -1.580628e-14, -8.376374e-15, -1.957694e-14, -1.720067e-14, 
    -5.093208e-15, -1.201266e-14, -8.425178e-15, -1.571778e-14, 
    -1.152465e-14, -1.914996e-14, -1.642859e-14, -1.148552e-14, 
    -5.706656e-15, -1.149579e-14, -2.493366e-14, -1.38365e-14, -1.647694e-14, 
    -2.014839e-14, -8.450903e-15, -1.128869e-14, -6.123346e-15, 
    -1.918924e-14, -8.553228e-15, -1.440029e-14, -1.244701e-14, 
    -1.408765e-14, -5.829819e-15, -1.131035e-14, -1.158487e-14, 
    -1.254433e-14, -1.898336e-14, -1.12609e-14, -1.923557e-14, -1.40939e-14, 
    -2.08602e-14, -9.764827e-15, -1.751272e-14, -6.007919e-15, -5.549935e-15, 
    -1.621309e-14, -1.780459e-14, -1.676058e-14, -1.838318e-14, 
    -1.255588e-14, -1.621191e-14, -7.743195e-15, -1.777625e-14, 
    -1.630536e-14, -1.493004e-14, -1.365761e-14, -1.101351e-14, 
    -1.467731e-14, -1.206812e-14, -1.00365e-14, -1.701146e-14, -1.563223e-14, 
    -1.910873e-14, -7.263286e-15, -1.553212e-14, -3.886367e-15, 
    -1.013623e-14, -1.57934e-14, -1.233619e-14, -5.644678e-15, -9.882703e-15, 
    -1.432925e-14, -5.698745e-15, -9.509276e-15, -1.901094e-14, 
    -1.312846e-14, -1.118442e-14, -1.369828e-14, -9.575321e-15, 
    -1.392922e-14, -8.614011e-15, -1.225686e-14, -1.673357e-14, 
    -1.974655e-14, -1.382981e-14, -1.62863e-14, -1.766018e-14, -9.089834e-15, 
    -2.093336e-14, -1.843198e-14, -1.766276e-14, -2.007472e-14, -2.525328e-14 ;

 ERRSOI =
  -6.059664e-10, -2.65541e-10, -4.444999e-10, -5.545744e-10, -2.299209e-10, 
    -4.435606e-10, -3.092726e-10, -4.954416e-10, -3.04193e-10, -3.904443e-10, 
    -3.825851e-10, -5.266568e-10, -4.300805e-10, -5.644635e-10, 
    -3.972198e-10, -3.844842e-10, -3.128045e-10, -3.744132e-10, 
    -4.299585e-10, -3.309238e-10, -4.609651e-10, -4.017794e-10, 
    -3.400238e-10, -4.615505e-10, -4.241322e-10, -2.763393e-10, 
    -2.774838e-10, -3.473827e-10, -3.915616e-10, -2.077853e-10, 
    -6.633894e-11, -3.008595e-10, -1.401217e-10, -2.787947e-10, -2.42861e-10, 
    -4.16945e-10, -3.388025e-10, -4.776252e-10, -3.454774e-10, -3.304016e-10, 
    -2.748863e-10, -4.6299e-10, -3.393218e-10, -1.973746e-10, -4.29863e-10, 
    -5.441061e-10, -2.066919e-10, -4.155568e-10, -3.21095e-10, -3.528947e-10, 
    -1.922169e-10, -3.354406e-10, -3.941893e-10, -5.547997e-10, 
    -5.157296e-10, -2.483766e-10, -3.265712e-10, -2.43831e-10, -4.20851e-10, 
    -4.375464e-10, -5.009591e-10, -2.951822e-10, -4.104719e-10, 
    -4.338005e-10, -4.281794e-10, -3.75954e-10, -1.484226e-10, -4.238665e-10, 
    -2.67039e-10, -3.122391e-10, -3.800536e-10, -3.215867e-10, -2.911265e-10, 
    -2.078463e-10, -3.681941e-10, -4.318703e-10, -3.143291e-10, -4.83292e-10, 
    -3.178882e-10, -3.690696e-10, -4.392083e-10, -6.565616e-10, 
    -4.176046e-10, -3.842969e-10, -3.243021e-10, -2.218467e-10, 
    -1.956927e-10, -4.180391e-10, -6.371884e-10, -4.296098e-10, 
    -4.451499e-10, -4.759553e-10, -3.184837e-10, -3.640886e-10, 
    -3.383617e-10, -3.992676e-10, -3.220045e-10, -3.012073e-10, 
    -4.173475e-10, -3.08951e-10, -1.155039e-10, -3.878317e-10, -4.419906e-10, 
    -3.51117e-10, -1.768444e-10, -1.44089e-10, -4.458635e-10, -3.735647e-10, 
    -2.711618e-10, -4.088145e-10, -4.068392e-10, -3.60322e-10, -2.738159e-10, 
    -3.85917e-10, -3.620755e-10, -4.616852e-10, -4.194593e-10, -4.71451e-10, 
    -3.059978e-10, -4.86537e-10, -4.0218e-10, -2.881927e-10, -4.710867e-10, 
    -3.080053e-10, -1.632396e-10, -2.634554e-10, -3.305864e-10, 
    -5.359851e-10, -3.085346e-10, -3.600895e-10, -3.46719e-10, -3.255556e-10, 
    -4.89723e-10, -3.228495e-10, -4.564235e-10, -3.845572e-10, -3.762644e-10, 
    -2.900543e-10, -4.381435e-10, -3.493712e-10, -1.48886e-10, -2.703051e-10, 
    -4.04227e-10, -3.744694e-10, -2.459127e-10, -3.931404e-10, -2.865442e-10, 
    -3.342947e-10, -4.065997e-10, -2.752003e-10, -3.501266e-10, 
    -3.285581e-10, -3.424742e-10, -4.159968e-10, -3.400094e-10, 
    -3.429415e-10, -2.918896e-10, -2.807982e-10, -3.624691e-10, 
    -3.347523e-10, -3.185245e-10, -3.331865e-10, -5.140963e-10, 
    -2.948015e-10, -4.884481e-10, -3.866196e-10, -3.425386e-10, 
    -5.523539e-10, -1.800778e-10, -4.759738e-10, -2.014841e-10, 
    -2.310215e-10, -1.248378e-10, -3.761141e-10, -3.641673e-10, 
    -4.199343e-10, -4.737953e-10, -3.623271e-10, -1.439912e-10, 
    -3.030762e-10, -2.791351e-10, -1.85686e-10, -2.874746e-10, -4.084153e-10, 
    -3.76715e-10, -3.561863e-10, -2.063277e-10, -4.326963e-10, -3.852988e-10, 
    -4.313484e-10, -3.909582e-10, -4.162494e-10, -4.904799e-10, 
    -3.607568e-10, -3.655407e-10, -4.319168e-10, -4.156493e-10, 
    -4.593205e-10, -4.045407e-10, -2.811871e-10, -2.352772e-10, 
    -3.225023e-10, -4.165989e-10, -2.874007e-10, -3.304397e-10, 
    -2.424198e-10, -2.148901e-10, -1.323107e-10, -4.587811e-10, 
    -4.703961e-10, -4.452684e-10, -3.855995e-10, -3.610559e-10, 
    -5.181783e-10, -3.034779e-10, -4.498827e-10, -2.769145e-10, 
    -3.974375e-10, -3.455204e-10, -3.366207e-10, -4.116497e-10, 
    -3.547811e-10, -4.130707e-10, -3.958862e-10, -5.299808e-10, 
    -5.262787e-10, -4.532259e-10, -3.141543e-10, -2.176958e-10, 
    -3.555623e-10, -3.630757e-10, -4.223187e-10, -3.187437e-10, 
    -3.306907e-10, -3.855362e-10, -4.476343e-10, -3.320258e-10, 
    -3.182135e-10, -2.157871e-10, -3.648882e-10, -4.372937e-10, 
    -3.035454e-10, -3.627248e-10, -4.90213e-10, -4.03577e-10, -4.749612e-10, 
    -3.215468e-10, -3.758893e-10, -4.064221e-10, -2.68319e-10, -3.549235e-10, 
    -3.535987e-10, -1.193173e-10, -5.090046e-10, -4.916704e-10, 
    -3.628255e-10, -5.06914e-10, -3.650969e-10, -1.347439e-10, -4.613222e-10, 
    -3.275436e-10, -4.167389e-10, -5.266396e-10, -2.150074e-10, 
    -2.815042e-11, -5.331251e-10, -3.294446e-10, -4.963067e-10, 
    -5.372303e-10, -2.312761e-10, -3.528938e-10, -4.381973e-10, -5.59736e-10, 
    -4.976978e-10, -2.589961e-10, -4.329071e-10, -4.499967e-10, 
    -3.337578e-10, -2.172619e-10, -3.983813e-10, -2.263774e-10, 
    -2.782026e-10, -6.058163e-10, -4.889112e-10, -1.841427e-10, 
    -4.099594e-10, -2.204361e-10, -3.057805e-10, -4.198624e-10, 
    -4.175777e-10, -3.92619e-10, -4.86209e-10, -2.232574e-10, -2.662007e-10, 
    -3.959935e-10, -4.984593e-10, -2.726948e-10, -3.11961e-10, -3.328753e-10, 
    -2.131604e-10, -4.606004e-10, -3.63162e-10, -4.39232e-10, -4.104112e-10, 
    -2.510055e-10, -1.749772e-10, -2.3317e-10, -5.302349e-10, -3.448641e-10, 
    -3.700363e-10, -1.848209e-10, -2.53134e-10, -4.669389e-10, -2.772576e-10, 
    -3.208243e-10, -2.622511e-10, -2.343212e-10, -4.497265e-10, 
    -3.272826e-10, -2.329953e-10, -2.406143e-10, -1.702121e-10, 
    -2.808037e-10, -5.196868e-10, -3.799712e-10, -3.297522e-10, 
    -3.322842e-10, -5.86238e-10, -4.717205e-10, -3.372673e-10, -3.518416e-10, 
    -3.978016e-10, -3.020076e-10, -2.918538e-10, -1.132868e-10, 
    -1.799326e-10, -1.359175e-10, -3.232596e-10 ;

 ERRSOL =
  1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 1.387779e-17, 
    1.387779e-17, 1.387779e-17, 1.387779e-17 ;

 ESAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 FAREA_BURNED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCEV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4 =
  1.89762e-16, 1.846676e-16, 1.856581e-16, 1.815484e-16, 1.838283e-16, 
    1.811371e-16, 1.887294e-16, 1.844652e-16, 1.871875e-16, 1.893036e-16, 
    1.735704e-16, 1.813651e-16, 1.654721e-16, 1.704452e-16, 1.579503e-16, 
    1.662459e-16, 1.562772e-16, 1.5819e-16, 1.524331e-16, 1.540825e-16, 
    1.467162e-16, 1.516717e-16, 1.428968e-16, 1.479e-16, 1.471173e-16, 
    1.518351e-16, 1.797969e-16, 1.745409e-16, 1.801082e-16, 1.793588e-16, 
    1.796952e-16, 1.837811e-16, 1.858397e-16, 1.901515e-16, 1.893688e-16, 
    1.86202e-16, 1.790218e-16, 1.814596e-16, 1.753159e-16, 1.754547e-16, 
    1.686127e-16, 1.716979e-16, 1.601947e-16, 1.634649e-16, 1.540137e-16, 
    1.56391e-16, 1.541253e-16, 1.548124e-16, 1.541164e-16, 1.576028e-16, 
    1.561091e-16, 1.591768e-16, 1.7112e-16, 1.676107e-16, 1.780754e-16, 
    1.843649e-16, 1.885423e-16, 1.91506e-16, 1.91087e-16, 1.902883e-16, 
    1.861835e-16, 1.823239e-16, 1.79382e-16, 1.774139e-16, 1.754746e-16, 
    1.696026e-16, 1.664946e-16, 1.595333e-16, 1.6079e-16, 1.586611e-16, 
    1.566275e-16, 1.532123e-16, 1.537745e-16, 1.522696e-16, 1.587175e-16, 
    1.544324e-16, 1.615058e-16, 1.595714e-16, 1.749463e-16, 1.80802e-16, 
    1.832896e-16, 1.854677e-16, 1.907649e-16, 1.871068e-16, 1.885489e-16, 
    1.851181e-16, 1.829378e-16, 1.840162e-16, 1.773601e-16, 1.79948e-16, 
    1.663104e-16, 1.721857e-16, 1.568647e-16, 1.605321e-16, 1.559856e-16, 
    1.583058e-16, 1.5433e-16, 1.579082e-16, 1.517096e-16, 1.503594e-16, 
    1.51282e-16, 1.477378e-16, 1.581065e-16, 1.541252e-16, 1.840464e-16, 
    1.838705e-16, 1.830512e-16, 1.866525e-16, 1.868728e-16, 1.901729e-16, 
    1.872366e-16, 1.85986e-16, 1.828115e-16, 1.809334e-16, 1.79148e-16, 
    1.752219e-16, 1.708362e-16, 1.647022e-16, 1.602944e-16, 1.573391e-16, 
    1.591514e-16, 1.575513e-16, 1.593399e-16, 1.601782e-16, 1.508652e-16, 
    1.560951e-16, 1.482477e-16, 1.48682e-16, 1.522338e-16, 1.486331e-16, 
    1.83747e-16, 1.847591e-16, 1.882725e-16, 1.85523e-16, 1.905323e-16, 
    1.877283e-16, 1.861159e-16, 1.798937e-16, 1.785267e-16, 1.772587e-16, 
    1.747544e-16, 1.7154e-16, 1.658998e-16, 1.609912e-16, 1.565092e-16, 
    1.568377e-16, 1.56722e-16, 1.557205e-16, 1.58201e-16, 1.553133e-16, 
    1.548285e-16, 1.560959e-16, 1.487402e-16, 1.50842e-16, 1.486913e-16, 
    1.500598e-16, 1.844302e-16, 1.827272e-16, 1.836474e-16, 1.819169e-16, 
    1.83136e-16, 1.777144e-16, 1.760886e-16, 1.6848e-16, 1.716032e-16, 
    1.666326e-16, 1.710984e-16, 1.703071e-16, 1.6647e-16, 1.708572e-16, 
    1.612617e-16, 1.677672e-16, 1.556816e-16, 1.621797e-16, 1.552743e-16, 
    1.565286e-16, 1.544519e-16, 1.525917e-16, 1.502513e-16, 1.459318e-16, 
    1.469322e-16, 1.433193e-16, 1.801882e-16, 1.779788e-16, 1.781736e-16, 
    1.758614e-16, 1.741511e-16, 1.704441e-16, 1.644969e-16, 1.667336e-16, 
    1.626274e-16, 1.618029e-16, 1.680412e-16, 1.64211e-16, 1.765002e-16, 
    1.74515e-16, 1.756972e-16, 1.800138e-16, 1.662179e-16, 1.73299e-16, 
    1.602215e-16, 1.640591e-16, 1.528569e-16, 1.584286e-16, 1.474828e-16, 
    1.428007e-16, 1.383937e-16, 1.332407e-16, 1.767732e-16, 1.782745e-16, 
    1.755864e-16, 1.718665e-16, 1.684149e-16, 1.63825e-16, 1.633554e-16, 
    1.624953e-16, 1.602676e-16, 1.583942e-16, 1.622232e-16, 1.579245e-16, 
    1.740542e-16, 1.656033e-16, 1.788419e-16, 1.74856e-16, 1.720859e-16, 
    1.733013e-16, 1.669893e-16, 1.655012e-16, 1.594531e-16, 1.6258e-16, 
    1.439563e-16, 1.521985e-16, 1.293166e-16, 1.357147e-16, 1.78799e-16, 
    1.767784e-16, 1.697445e-16, 1.730916e-16, 1.635187e-16, 1.611615e-16, 
    1.592452e-16, 1.56795e-16, 1.565306e-16, 1.550787e-16, 1.574578e-16, 
    1.551728e-16, 1.638152e-16, 1.599536e-16, 1.705489e-16, 1.679705e-16, 
    1.691568e-16, 1.704578e-16, 1.664422e-16, 1.621629e-16, 1.620717e-16, 
    1.606993e-16, 1.568307e-16, 1.634799e-16, 1.428915e-16, 1.556088e-16, 
    1.745749e-16, 1.706817e-16, 1.701259e-16, 1.716341e-16, 1.613978e-16, 
    1.651074e-16, 1.551142e-16, 1.578156e-16, 1.533892e-16, 1.555889e-16, 
    1.559125e-16, 1.587372e-16, 1.604956e-16, 1.649372e-16, 1.685505e-16, 
    1.714154e-16, 1.707493e-16, 1.676021e-16, 1.619011e-16, 1.565065e-16, 
    1.576883e-16, 1.537257e-16, 1.642129e-16, 1.59816e-16, 1.615154e-16, 
    1.570839e-16, 1.66793e-16, 1.585245e-16, 1.689057e-16, 1.679958e-16, 
    1.65181e-16, 1.595175e-16, 1.582648e-16, 1.569265e-16, 1.577523e-16, 
    1.617565e-16, 1.624125e-16, 1.652495e-16, 1.660326e-16, 1.68194e-16, 
    1.699831e-16, 1.683484e-16, 1.666314e-16, 1.617549e-16, 1.57359e-16, 
    1.525652e-16, 1.51392e-16, 1.457878e-16, 1.503495e-16, 1.428206e-16, 
    1.492211e-16, 1.3814e-16, 1.580457e-16, 1.4941e-16, 1.65053e-16, 
    1.633685e-16, 1.603209e-16, 1.533298e-16, 1.571048e-16, 1.526901e-16, 
    1.624382e-16, 1.674934e-16, 1.688015e-16, 1.712412e-16, 1.687457e-16, 
    1.689487e-16, 1.665605e-16, 1.67328e-16, 1.61593e-16, 1.646738e-16, 
    1.559205e-16, 1.52725e-16, 1.436978e-16, 1.38161e-16, 1.325231e-16, 
    1.300332e-16, 1.292753e-16, 1.289584e-16 ;

 FCH4TOCO2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCH4_DFSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FCOV =
  0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584 ;

 FCTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FGEV =
  22.01506, 22.07914, 22.0667, 22.11838, 22.08974, 22.12356, 22.02809, 
    22.08165, 22.04748, 22.02089, 22.21867, 22.12069, 22.32102, 22.25834, 
    22.41604, 22.31121, 22.43722, 22.41311, 22.48593, 22.46507, 22.55809, 
    22.49556, 22.60652, 22.54321, 22.55307, 22.49348, 22.14049, 22.20643, 
    22.13656, 22.14597, 22.14177, 22.0903, 22.06432, 22.01023, 22.02006, 
    22.05983, 22.1502, 22.11957, 22.19697, 22.19522, 22.28147, 22.24257, 
    22.38778, 22.34649, 22.46594, 22.43586, 22.46451, 22.45584, 22.46462, 
    22.42053, 22.43941, 22.40065, 22.24983, 22.29409, 22.16215, 22.08282, 
    22.03042, 21.9932, 21.99846, 22.00847, 22.06006, 22.10869, 22.14574, 
    22.17053, 22.19497, 22.2688, 22.30812, 22.39608, 22.38028, 22.40711, 
    22.43288, 22.47605, 22.46895, 22.48796, 22.40646, 22.46058, 22.37126, 
    22.39567, 22.2013, 22.12784, 22.09637, 22.06908, 22.0025, 22.04845, 
    22.03032, 22.07353, 22.10095, 22.0874, 22.17121, 22.1386, 22.31045, 
    22.23636, 22.42987, 22.38353, 22.441, 22.41168, 22.46189, 22.4167, 
    22.49506, 22.5121, 22.50045, 22.54532, 22.41419, 22.46448, 22.08701, 
    22.08921, 22.09954, 22.05416, 22.0514, 22.00994, 22.04686, 22.06256, 
    22.10257, 22.12618, 22.14866, 22.19812, 22.25337, 22.33079, 22.38653, 
    22.4239, 22.401, 22.42121, 22.39861, 22.38803, 22.50569, 22.43957, 
    22.53886, 22.53338, 22.4884, 22.53399, 22.09077, 22.07805, 22.03383, 
    22.06844, 22.00544, 22.04065, 22.06089, 22.13921, 22.15651, 22.17245, 
    22.20403, 22.24456, 22.31569, 22.37769, 22.43439, 22.43024, 22.4317, 
    22.44434, 22.41299, 22.44949, 22.45559, 22.4396, 22.53264, 22.50605, 
    22.53326, 22.51595, 22.0822, 22.10361, 22.09203, 22.11379, 22.09844, 
    22.16664, 22.1871, 22.28306, 22.24374, 22.30642, 22.25013, 22.26008, 
    22.30833, 22.25319, 22.37421, 22.29202, 22.44483, 22.36253, 22.44998, 
    22.43414, 22.4604, 22.48389, 22.51352, 22.56812, 22.55548, 22.60122, 
    22.13558, 22.16335, 22.16096, 22.19008, 22.21162, 22.2584, 22.33343, 
    22.30522, 22.35708, 22.36747, 22.28873, 22.33701, 22.18199, 22.20694, 
    22.19213, 22.13773, 22.31164, 22.22228, 22.38744, 22.33897, 22.48053, 
    22.41003, 22.54851, 22.60764, 22.66362, 22.72877, 22.17858, 22.15969, 
    22.19356, 22.24035, 22.28397, 22.34191, 22.34788, 22.35872, 22.38689, 
    22.41056, 22.36209, 22.4165, 22.21261, 22.31943, 22.1525, 22.20263, 
    22.23762, 22.22233, 22.30201, 22.32079, 22.39711, 22.35768, 22.59299, 
    22.48877, 22.77861, 22.69745, 22.15308, 22.17854, 22.26715, 22.22499, 
    22.34582, 22.37557, 22.39981, 22.43073, 22.43411, 22.45244, 22.4224, 
    22.45127, 22.34204, 22.39084, 22.25709, 22.28958, 22.27465, 22.25824, 
    22.30891, 22.36284, 22.36409, 22.38137, 22.42994, 22.34631, 22.60628, 
    22.44543, 22.20631, 22.25528, 22.26239, 22.2434, 22.37258, 22.32573, 
    22.45201, 22.41787, 22.47383, 22.44601, 22.44191, 22.40622, 22.38399, 
    22.32786, 22.28225, 22.24616, 22.25456, 22.29421, 22.36616, 22.43437, 
    22.41941, 22.46958, 22.33704, 22.39253, 22.37105, 22.4271, 22.30445, 
    22.40859, 22.27782, 22.2893, 22.3248, 22.39623, 22.41219, 22.42906, 
    22.41867, 22.36801, 22.35975, 22.32396, 22.31403, 22.28681, 22.26423, 
    22.28483, 22.30646, 22.36807, 22.42359, 22.48421, 22.49909, 22.56977, 
    22.5121, 22.60715, 22.52612, 22.66655, 22.41477, 22.52394, 22.32645, 
    22.34772, 22.38611, 22.47445, 22.42684, 22.48256, 22.35944, 22.29553, 
    22.27913, 22.24834, 22.27983, 22.27728, 22.30742, 22.29774, 22.37012, 
    22.33123, 22.44179, 22.48215, 22.59639, 22.66646, 22.73801, 22.76957, 
    22.77918, 22.7832 ;

 FGR =
  -386.0582, -387.156, -386.9427, -387.8278, -387.3371, -387.9164, -386.2811, 
    -387.1993, -386.6133, -386.1574, -389.5446, -387.8674, -391.2898, 
    -390.2197, -392.9088, -391.1229, -393.269, -392.858, -394.0968, -393.742, 
    -395.3248, -394.2606, -396.1464, -395.071, -395.239, -394.2254, 
    -388.2056, -389.3355, -388.1385, -388.2996, -388.2275, -387.347, 
    -386.9028, -385.9748, -386.1434, -386.8253, -388.3721, -387.8475, 
    -389.1711, -389.1412, -390.6143, -389.9502, -392.4266, -391.7229, 
    -393.7568, -393.2452, -393.7327, -393.585, -393.7346, -392.9843, 
    -393.3057, -392.6458, -390.0744, -390.8299, -388.5762, -387.2201, 
    -386.3212, -385.6828, -385.773, -385.9449, -386.8293, -387.6613, 
    -388.2952, -388.7191, -389.1369, -390.3997, -391.0697, -392.5685, 
    -392.2986, -392.7563, -393.1944, -393.929, -393.8082, -394.1317, 
    -392.7447, -393.6663, -392.1448, -392.5609, -389.2481, -387.9891, 
    -387.452, -386.9836, -385.8424, -386.6304, -386.3197, -387.0593, 
    -387.529, -387.2968, -388.7307, -388.1731, -391.1094, -389.8447, 
    -393.1433, -392.3541, -393.3325, -392.8334, -393.6884, -392.9189, 
    -394.2523, -394.5423, -394.3441, -395.1064, -392.8762, -393.7324, 
    -387.2902, -387.328, -387.5047, -386.7282, -386.6808, -385.97, -386.6027, 
    -386.8719, -387.5564, -387.9608, -388.3454, -389.1911, -390.1352, 
    -391.456, -392.4052, -393.0414, -392.6515, -392.9957, -392.6108, 
    -392.4305, -394.4335, -393.3086, -394.9968, -394.9034, -394.1393, 
    -394.914, -387.3546, -387.1367, -386.3794, -386.9721, -385.8926, 
    -386.4966, -386.8437, -388.1843, -388.4794, -388.7523, -389.2919, 
    -389.9841, -391.1982, -392.255, -393.22, -393.1493, -393.1742, -393.3895, 
    -392.8558, -393.4771, -393.5811, -393.3087, -394.8909, -394.439, 
    -394.9015, -394.6072, -387.2076, -387.5744, -387.3762, -387.7488, 
    -387.4861, -388.6536, -389.0036, -390.6422, -389.9704, -391.0403, 
    -390.0793, -390.2494, -391.0742, -390.1313, -392.1963, -390.7954, 
    -393.3978, -391.998, -393.4855, -393.2158, -393.6626, -394.0624, 
    -394.5659, -395.4942, -395.2794, -396.056, -388.1214, -388.597, 
    -388.5555, -389.0535, -389.4217, -390.2202, -391.5005, -391.0192, 
    -391.9033, -392.0806, -390.7378, -391.5618, -388.9156, -389.3426, 
    -389.0887, -388.1587, -391.1295, -389.6046, -392.4208, -391.5949, 
    -394.0054, -392.8062, -395.161, -396.1663, -397.1144, -398.2197, 
    -388.857, -388.5338, -389.1129, -389.9131, -390.657, -391.6452, 
    -391.7465, -391.9315, -392.4112, -392.8143, -391.9895, -392.9154, 
    -389.4407, -391.2621, -388.4112, -389.269, -389.8662, -389.6047, 
    -390.9643, -391.2846, -392.5859, -391.9135, -395.9178, -394.1463, 
    -399.0627, -397.6889, -388.4208, -388.8561, -390.3704, -389.6499, 
    -391.7114, -392.2186, -392.6313, -393.1581, -393.2153, -393.5274, 
    -393.0158, -393.5074, -391.6473, -392.4786, -390.1978, -390.7527, 
    -390.4976, -390.2174, -391.0821, -392.0024, -392.0228, -392.3178, 
    -393.1477, -391.7198, -396.145, -393.411, -389.3307, -390.1681, 
    -390.2886, -389.9641, -392.1677, -391.3692, -393.5199, -392.9388, 
    -393.8911, -393.4178, -393.3482, -392.7405, -392.3619, -391.4056, 
    -390.6277, -390.0112, -390.1546, -390.8319, -392.0589, -393.2201, 
    -392.9656, -393.8188, -391.5619, -392.5079, -392.142, -393.0961, 
    -391.0063, -392.7837, -390.5517, -390.7475, -391.3533, -392.5715, 
    -392.8422, -393.1298, -392.9525, -392.0902, -391.9492, -391.3388, 
    -391.1699, -390.7049, -390.3197, -390.6715, -391.0408, -392.0909, 
    -393.0367, -394.068, -394.3207, -395.5237, -394.5434, -396.1601, 
    -394.7841, -397.1666, -392.8878, -394.7451, -391.3811, -391.7438, 
    -392.3988, -393.9028, -393.0916, -394.0406, -391.9438, -390.8549, 
    -390.574, -390.0486, -390.5861, -390.5424, -391.0566, -390.8914, 
    -392.1257, -391.4627, -393.3463, -394.0333, -395.9743, -397.1635, 
    -398.3749, -398.9093, -399.072, -399.14 ;

 FGR12 =
  -50.28005, -50.34876, -50.33542, -50.39087, -50.36014, -50.39644, 
    -50.29401, -50.35144, -50.3148, -50.28629, -50.49866, -50.39338, 
    -50.60887, -50.54137, -50.71137, -50.59832, -50.73425, -50.70823, 
    -50.7869, -50.76435, -50.86497, -50.79732, -50.91743, -50.84887, 
    -50.85953, -50.79507, -50.41463, -50.4855, -50.41041, -50.42051, 
    -50.41599, -50.36074, -50.33285, -50.27487, -50.28541, -50.32804, 
    -50.42506, -50.39216, -50.47535, -50.47347, -50.56627, -50.5244, 
    -50.68087, -50.63634, -50.76529, -50.7328, -50.76374, -50.75437, 
    -50.76387, -50.71624, -50.73662, -50.69477, -50.53221, -50.57985, 
    -50.4379, -50.35271, -50.2965, -50.25662, -50.26225, -50.27298, 
    -50.32829, -50.38047, -50.42028, -50.44691, -50.47321, -50.55262, 
    -50.59497, -50.68983, -50.67279, -50.70174, -50.72957, -50.77621, 
    -50.76855, -50.78909, -50.70105, -50.7595, -50.66306, -50.68939, 
    -50.47999, -50.40105, -50.36725, -50.33797, -50.26658, -50.31583, 
    -50.2964, -50.34274, -50.37217, -50.35763, -50.44764, -50.41261, 
    -50.59747, -50.51772, -50.72631, -50.67629, -50.73833, -50.70668, 
    -50.76091, -50.7121, -50.79677, -50.8152, -50.8026, -50.85114, -50.70939, 
    -50.76371, -50.35721, -50.35957, -50.37065, -50.32196, -50.319, 
    -50.27457, -50.31414, -50.33097, -50.37391, -50.39927, -50.42342, 
    -50.47658, -50.53602, -50.6194, -50.67953, -50.71986, -50.69515, 
    -50.71697, -50.69257, -50.68115, -50.80826, -50.7368, -50.84416, 
    -50.83822, -50.78957, -50.83889, -50.36124, -50.3476, -50.30016, 
    -50.33728, -50.26973, -50.30748, -50.32919, -50.41325, -50.43185, 
    -50.44898, -50.48294, -50.52653, -50.60313, -50.66998, -50.7312, 
    -50.72672, -50.72829, -50.74195, -50.7081, -50.74751, -50.7541, 
    -50.73683, -50.83742, -50.80866, -50.83809, -50.81937, -50.35205, 
    -50.37503, -50.3626, -50.38595, -50.36948, -50.44273, -50.46474, 
    -50.56797, -50.52566, -50.59314, -50.53253, -50.54324, -50.5952, 
    -50.53583, -50.66622, -50.57763, -50.74247, -50.65365, -50.74804, 
    -50.73094, -50.7593, -50.78469, -50.81674, -50.87583, -50.86216, 
    -50.91169, -50.40936, -50.43919, -50.43663, -50.46793, -50.4911, 
    -50.54143, -50.62225, -50.59186, -50.64775, -50.65897, -50.57409, 
    -50.62611, -50.45924, -50.48606, -50.47013, -50.41168, -50.59876, 
    -50.50257, -50.6805, -50.62823, -50.78106, -50.7049, -50.85461, 
    -50.91865, -50.97929, -51.04989, -50.45556, -50.43527, -50.47168, 
    -50.52201, -50.56897, -50.6314, -50.63784, -50.64953, -50.67992, 
    -50.70547, -50.65317, -50.71187, -50.49217, -50.60715, -50.42755, 
    -50.48142, -50.51907, -50.50262, -50.5884, -50.60863, -50.69095, 
    -50.64841, -50.90277, -50.78997, -51.10397, -51.01594, -50.42817, 
    -50.45553, -50.55085, -50.50548, -50.63561, -50.6677, -50.69387, 
    -50.72724, -50.7309, -50.7507, -50.71825, -50.74944, -50.63154, 
    -50.68417, -50.54003, -50.57501, -50.55893, -50.54126, -50.59584, 
    -50.65396, -50.65532, -50.67397, -50.72638, -50.63615, -50.91716, 
    -50.74314, -50.48539, -50.53806, -50.54573, -50.52529, -50.66447, 
    -50.61396, -50.75023, -50.71337, -50.77382, -50.74376, -50.73933, 
    -50.70079, -50.67678, -50.61626, -50.56711, -50.52827, -50.5373, -50.58, 
    -50.65756, -50.73117, -50.71503, -50.76922, -50.62616, -50.68601, 
    -50.66284, -50.72333, -50.59103, -50.70332, -50.56235, -50.5747, 
    -50.61296, -50.68999, -50.70724, -50.72544, -50.71422, -50.65955, 
    -50.65064, -50.61205, -50.60135, -50.57202, -50.54771, -50.56989, 
    -50.59319, -50.65961, -50.71954, -50.78503, -50.80114, -50.87761, 
    -50.8152, -50.91811, -50.83039, -50.98244, -50.71002, -50.828, -50.61474, 
    -50.63766, -50.67908, -50.77447, -50.72305, -50.78325, -50.6503, 
    -50.58142, -50.56375, -50.53061, -50.56451, -50.56176, -50.59423, 
    -50.5838, -50.66182, -50.6199, -50.73919, -50.78281, -50.90646, 
    -50.98235, -51.05991, -51.09416, -51.1046, -51.10896 ;

 FGR_R =
  -386.0582, -387.156, -386.9427, -387.8278, -387.3371, -387.9164, -386.2811, 
    -387.1993, -386.6133, -386.1574, -389.5446, -387.8674, -391.2898, 
    -390.2197, -392.9088, -391.1229, -393.269, -392.858, -394.0968, -393.742, 
    -395.3248, -394.2606, -396.1464, -395.071, -395.239, -394.2254, 
    -388.2056, -389.3355, -388.1385, -388.2996, -388.2275, -387.347, 
    -386.9028, -385.9748, -386.1434, -386.8253, -388.3721, -387.8475, 
    -389.1711, -389.1412, -390.6143, -389.9502, -392.4266, -391.7229, 
    -393.7568, -393.2452, -393.7327, -393.585, -393.7346, -392.9843, 
    -393.3057, -392.6458, -390.0744, -390.8299, -388.5762, -387.2201, 
    -386.3212, -385.6828, -385.773, -385.9449, -386.8293, -387.6613, 
    -388.2952, -388.7191, -389.1369, -390.3997, -391.0697, -392.5685, 
    -392.2986, -392.7563, -393.1944, -393.929, -393.8082, -394.1317, 
    -392.7447, -393.6663, -392.1448, -392.5609, -389.2481, -387.9891, 
    -387.452, -386.9836, -385.8424, -386.6304, -386.3197, -387.0593, 
    -387.529, -387.2968, -388.7307, -388.1731, -391.1094, -389.8447, 
    -393.1433, -392.3541, -393.3325, -392.8334, -393.6884, -392.9189, 
    -394.2523, -394.5423, -394.3441, -395.1064, -392.8762, -393.7324, 
    -387.2902, -387.328, -387.5047, -386.7282, -386.6808, -385.97, -386.6027, 
    -386.8719, -387.5564, -387.9608, -388.3454, -389.1911, -390.1352, 
    -391.456, -392.4052, -393.0414, -392.6515, -392.9957, -392.6108, 
    -392.4305, -394.4335, -393.3086, -394.9968, -394.9034, -394.1393, 
    -394.914, -387.3546, -387.1367, -386.3794, -386.9721, -385.8926, 
    -386.4966, -386.8437, -388.1843, -388.4794, -388.7523, -389.2919, 
    -389.9841, -391.1982, -392.255, -393.22, -393.1493, -393.1742, -393.3895, 
    -392.8558, -393.4771, -393.5811, -393.3087, -394.8909, -394.439, 
    -394.9015, -394.6072, -387.2076, -387.5744, -387.3762, -387.7488, 
    -387.4861, -388.6536, -389.0036, -390.6422, -389.9704, -391.0403, 
    -390.0793, -390.2494, -391.0742, -390.1313, -392.1963, -390.7954, 
    -393.3978, -391.998, -393.4855, -393.2158, -393.6626, -394.0624, 
    -394.5659, -395.4942, -395.2794, -396.056, -388.1214, -388.597, 
    -388.5555, -389.0535, -389.4217, -390.2202, -391.5005, -391.0192, 
    -391.9033, -392.0806, -390.7378, -391.5618, -388.9156, -389.3426, 
    -389.0887, -388.1587, -391.1295, -389.6046, -392.4208, -391.5949, 
    -394.0054, -392.8062, -395.161, -396.1663, -397.1144, -398.2197, 
    -388.857, -388.5338, -389.1129, -389.9131, -390.657, -391.6452, 
    -391.7465, -391.9315, -392.4112, -392.8143, -391.9895, -392.9154, 
    -389.4407, -391.2621, -388.4112, -389.269, -389.8662, -389.6047, 
    -390.9643, -391.2846, -392.5859, -391.9135, -395.9178, -394.1463, 
    -399.0627, -397.6889, -388.4208, -388.8561, -390.3704, -389.6499, 
    -391.7114, -392.2186, -392.6313, -393.1581, -393.2153, -393.5274, 
    -393.0158, -393.5074, -391.6473, -392.4786, -390.1978, -390.7527, 
    -390.4976, -390.2174, -391.0821, -392.0024, -392.0228, -392.3178, 
    -393.1477, -391.7198, -396.145, -393.411, -389.3307, -390.1681, 
    -390.2886, -389.9641, -392.1677, -391.3692, -393.5199, -392.9388, 
    -393.8911, -393.4178, -393.3482, -392.7405, -392.3619, -391.4056, 
    -390.6277, -390.0112, -390.1546, -390.8319, -392.0589, -393.2201, 
    -392.9656, -393.8188, -391.5619, -392.5079, -392.142, -393.0961, 
    -391.0063, -392.7837, -390.5517, -390.7475, -391.3533, -392.5715, 
    -392.8422, -393.1298, -392.9525, -392.0902, -391.9492, -391.3388, 
    -391.1699, -390.7049, -390.3197, -390.6715, -391.0408, -392.0909, 
    -393.0367, -394.068, -394.3207, -395.5237, -394.5434, -396.1601, 
    -394.7841, -397.1666, -392.8878, -394.7451, -391.3811, -391.7438, 
    -392.3988, -393.9028, -393.0916, -394.0406, -391.9438, -390.8549, 
    -390.574, -390.0486, -390.5861, -390.5424, -391.0566, -390.8914, 
    -392.1257, -391.4627, -393.3463, -394.0333, -395.9743, -397.1635, 
    -398.3749, -398.9093, -399.072, -399.14 ;

 FGR_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FINUNDATED_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FIRA =
  46.2159, 46.29252, 46.27764, 46.3394, 46.30516, 46.34559, 46.23146, 
    46.29554, 46.25465, 46.22283, 46.45919, 46.34217, 46.58097, 46.50631, 
    46.69393, 46.56932, 46.71907, 46.69039, 46.77682, 46.75207, 46.86248, 
    46.78825, 46.91981, 46.84479, 46.8565, 46.78579, 46.36577, 46.44461, 
    46.36109, 46.37233, 46.3673, 46.30585, 46.27485, 46.21008, 46.22185, 
    46.26944, 46.37739, 46.34078, 46.43315, 46.43106, 46.53385, 46.4875, 
    46.66029, 46.6112, 46.7531, 46.71741, 46.75142, 46.74111, 46.75155, 
    46.6992, 46.72163, 46.67558, 46.49617, 46.54889, 46.39164, 46.29699, 
    46.23426, 46.1897, 46.196, 46.208, 46.26971, 46.32779, 46.37202, 
    46.40161, 46.43076, 46.51886, 46.56561, 46.67019, 46.65136, 46.68329, 
    46.71386, 46.76511, 46.75668, 46.77925, 46.68248, 46.74678, 46.64063, 
    46.66966, 46.4385, 46.35067, 46.31317, 46.28049, 46.20084, 46.25583, 
    46.23415, 46.28578, 46.31855, 46.30235, 46.40242, 46.36351, 46.56838, 
    46.48014, 46.71029, 46.65523, 46.7235, 46.68867, 46.74833, 46.69464, 
    46.78767, 46.8079, 46.79407, 46.84726, 46.69166, 46.7514, 46.30189, 
    46.30453, 46.31686, 46.26266, 46.25936, 46.20975, 46.25391, 46.2727, 
    46.32047, 46.34869, 46.37553, 46.43454, 46.50041, 46.59257, 46.6588, 
    46.70319, 46.67598, 46.7, 46.67315, 46.66056, 46.8003, 46.72183, 
    46.83961, 46.8331, 46.77978, 46.83383, 46.30639, 46.29118, 46.23832, 
    46.27969, 46.20435, 46.2465, 46.27072, 46.36428, 46.38488, 46.40392, 
    46.44158, 46.48988, 46.57458, 46.64832, 46.71564, 46.71072, 46.71245, 
    46.72747, 46.69024, 46.73359, 46.74084, 46.72184, 46.83223, 46.80069, 
    46.83296, 46.81244, 46.29613, 46.32172, 46.30789, 46.33389, 46.31556, 
    46.39703, 46.42146, 46.53579, 46.48891, 46.56357, 46.49651, 46.50838, 
    46.56592, 46.50015, 46.64421, 46.54647, 46.72805, 46.63038, 46.73417, 
    46.71535, 46.74652, 46.77442, 46.80955, 46.87431, 46.85932, 46.91351, 
    46.3599, 46.39308, 46.39019, 46.42494, 46.45063, 46.50635, 46.59568, 
    46.5621, 46.62378, 46.63615, 46.54246, 46.59995, 46.41531, 46.44511, 
    46.42739, 46.3625, 46.56979, 46.46339, 46.65989, 46.60226, 46.77044, 
    46.68677, 46.85106, 46.92119, 46.98735, 47.06445, 46.41123, 46.38868, 
    46.42908, 46.48492, 46.53682, 46.60577, 46.61284, 46.62575, 46.65922, 
    46.68734, 46.6298, 46.6944, 46.45195, 46.57904, 46.38012, 46.43998, 
    46.48164, 46.4634, 46.55827, 46.58062, 46.6714, 46.62449, 46.90385, 
    46.78027, 47.12326, 47.02742, 46.38079, 46.41117, 46.51682, 46.46656, 
    46.61039, 46.64577, 46.67457, 46.71132, 46.71532, 46.73709, 46.7014, 
    46.7357, 46.60592, 46.66392, 46.50479, 46.5435, 46.5257, 46.50616, 
    46.56648, 46.63069, 46.63212, 46.6527, 46.71058, 46.61097, 46.9197, 
    46.72895, 46.44428, 46.50271, 46.51112, 46.48848, 46.64223, 46.58651, 
    46.73657, 46.69603, 46.76247, 46.72945, 46.72459, 46.68219, 46.65578, 
    46.58906, 46.53478, 46.49177, 46.50177, 46.54902, 46.63463, 46.71565, 
    46.6979, 46.75742, 46.59996, 46.66596, 46.64043, 46.707, 46.56119, 
    46.68519, 46.52948, 46.54314, 46.58541, 46.6704, 46.68929, 46.70935, 
    46.69698, 46.63682, 46.62698, 46.58439, 46.57261, 46.54017, 46.51329, 
    46.53783, 46.5636, 46.63686, 46.70285, 46.77481, 46.79244, 46.87636, 
    46.80797, 46.92075, 46.82475, 46.99097, 46.69246, 46.82204, 46.58735, 
    46.61265, 46.65835, 46.76328, 46.70669, 46.7729, 46.6266, 46.55062, 
    46.53104, 46.49437, 46.53188, 46.52883, 46.56471, 46.55318, 46.6393, 
    46.59304, 46.72445, 46.77239, 46.90781, 46.99076, 47.07528, 47.11256, 
    47.12391, 47.12865 ;

 FIRA_R =
  46.2159, 46.29252, 46.27764, 46.3394, 46.30516, 46.34559, 46.23146, 
    46.29554, 46.25465, 46.22283, 46.45919, 46.34217, 46.58097, 46.50631, 
    46.69393, 46.56932, 46.71907, 46.69039, 46.77682, 46.75207, 46.86248, 
    46.78825, 46.91981, 46.84479, 46.8565, 46.78579, 46.36577, 46.44461, 
    46.36109, 46.37233, 46.3673, 46.30585, 46.27485, 46.21008, 46.22185, 
    46.26944, 46.37739, 46.34078, 46.43315, 46.43106, 46.53385, 46.4875, 
    46.66029, 46.6112, 46.7531, 46.71741, 46.75142, 46.74111, 46.75155, 
    46.6992, 46.72163, 46.67558, 46.49617, 46.54889, 46.39164, 46.29699, 
    46.23426, 46.1897, 46.196, 46.208, 46.26971, 46.32779, 46.37202, 
    46.40161, 46.43076, 46.51886, 46.56561, 46.67019, 46.65136, 46.68329, 
    46.71386, 46.76511, 46.75668, 46.77925, 46.68248, 46.74678, 46.64063, 
    46.66966, 46.4385, 46.35067, 46.31317, 46.28049, 46.20084, 46.25583, 
    46.23415, 46.28578, 46.31855, 46.30235, 46.40242, 46.36351, 46.56838, 
    46.48014, 46.71029, 46.65523, 46.7235, 46.68867, 46.74833, 46.69464, 
    46.78767, 46.8079, 46.79407, 46.84726, 46.69166, 46.7514, 46.30189, 
    46.30453, 46.31686, 46.26266, 46.25936, 46.20975, 46.25391, 46.2727, 
    46.32047, 46.34869, 46.37553, 46.43454, 46.50041, 46.59257, 46.6588, 
    46.70319, 46.67598, 46.7, 46.67315, 46.66056, 46.8003, 46.72183, 
    46.83961, 46.8331, 46.77978, 46.83383, 46.30639, 46.29118, 46.23832, 
    46.27969, 46.20435, 46.2465, 46.27072, 46.36428, 46.38488, 46.40392, 
    46.44158, 46.48988, 46.57458, 46.64832, 46.71564, 46.71072, 46.71245, 
    46.72747, 46.69024, 46.73359, 46.74084, 46.72184, 46.83223, 46.80069, 
    46.83296, 46.81244, 46.29613, 46.32172, 46.30789, 46.33389, 46.31556, 
    46.39703, 46.42146, 46.53579, 46.48891, 46.56357, 46.49651, 46.50838, 
    46.56592, 46.50015, 46.64421, 46.54647, 46.72805, 46.63038, 46.73417, 
    46.71535, 46.74652, 46.77442, 46.80955, 46.87431, 46.85932, 46.91351, 
    46.3599, 46.39308, 46.39019, 46.42494, 46.45063, 46.50635, 46.59568, 
    46.5621, 46.62378, 46.63615, 46.54246, 46.59995, 46.41531, 46.44511, 
    46.42739, 46.3625, 46.56979, 46.46339, 46.65989, 46.60226, 46.77044, 
    46.68677, 46.85106, 46.92119, 46.98735, 47.06445, 46.41123, 46.38868, 
    46.42908, 46.48492, 46.53682, 46.60577, 46.61284, 46.62575, 46.65922, 
    46.68734, 46.6298, 46.6944, 46.45195, 46.57904, 46.38012, 46.43998, 
    46.48164, 46.4634, 46.55827, 46.58062, 46.6714, 46.62449, 46.90385, 
    46.78027, 47.12326, 47.02742, 46.38079, 46.41117, 46.51682, 46.46656, 
    46.61039, 46.64577, 46.67457, 46.71132, 46.71532, 46.73709, 46.7014, 
    46.7357, 46.60592, 46.66392, 46.50479, 46.5435, 46.5257, 46.50616, 
    46.56648, 46.63069, 46.63212, 46.6527, 46.71058, 46.61097, 46.9197, 
    46.72895, 46.44428, 46.50271, 46.51112, 46.48848, 46.64223, 46.58651, 
    46.73657, 46.69603, 46.76247, 46.72945, 46.72459, 46.68219, 46.65578, 
    46.58906, 46.53478, 46.49177, 46.50177, 46.54902, 46.63463, 46.71565, 
    46.6979, 46.75742, 46.59996, 46.66596, 46.64043, 46.707, 46.56119, 
    46.68519, 46.52948, 46.54314, 46.58541, 46.6704, 46.68929, 46.70935, 
    46.69698, 46.63682, 46.62698, 46.58439, 46.57261, 46.54017, 46.51329, 
    46.53783, 46.5636, 46.63686, 46.70285, 46.77481, 46.79244, 46.87636, 
    46.80797, 46.92075, 46.82475, 46.99097, 46.69246, 46.82204, 46.58735, 
    46.61265, 46.65835, 46.76328, 46.70669, 46.7729, 46.6266, 46.55062, 
    46.53104, 46.49437, 46.53188, 46.52883, 46.56471, 46.55318, 46.6393, 
    46.59304, 46.72445, 46.77239, 46.90781, 46.99076, 47.07528, 47.11256, 
    47.12391, 47.12865 ;

 FIRA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FIRE =
  260.562, 260.6387, 260.6238, 260.6855, 260.6513, 260.6917, 260.5776, 
    260.6417, 260.6008, 260.569, 260.8053, 260.6883, 260.9271, 260.8524, 
    261.0401, 260.9155, 261.0652, 261.0365, 261.123, 261.0982, 261.2086, 
    261.1344, 261.266, 261.1909, 261.2026, 261.1319, 260.7119, 260.7907, 
    260.7072, 260.7185, 260.7134, 260.652, 260.621, 260.5562, 260.568, 
    260.6156, 260.7235, 260.6869, 260.7793, 260.7772, 260.88, 260.8336, 
    261.0064, 260.9573, 261.0992, 261.0635, 261.0976, 261.0872, 261.0977, 
    261.0453, 261.0678, 261.0217, 260.8423, 260.895, 260.7378, 260.6431, 
    260.5804, 260.5359, 260.5421, 260.5541, 260.6158, 260.6739, 260.7182, 
    260.7477, 260.7769, 260.865, 260.9117, 261.0163, 260.9975, 261.0294, 
    261.06, 261.1113, 261.1028, 261.1254, 261.0286, 261.0929, 260.9868, 
    261.0158, 260.7846, 260.6968, 260.6593, 260.6266, 260.547, 260.602, 
    260.5803, 260.6319, 260.6647, 260.6485, 260.7486, 260.7097, 260.9145, 
    260.8263, 261.0564, 261.0014, 261.0696, 261.0348, 261.0945, 261.0408, 
    261.1338, 261.1541, 261.1402, 261.1934, 261.0378, 261.0975, 260.648, 
    260.6507, 260.663, 260.6088, 260.6055, 260.5559, 260.6, 260.6188, 
    260.6666, 260.6948, 260.7217, 260.7807, 260.8466, 260.9387, 261.0049, 
    261.0493, 261.0221, 261.0461, 261.0193, 261.0067, 261.1465, 261.068, 
    261.1858, 261.1792, 261.1259, 261.18, 260.6525, 260.6373, 260.5845, 
    260.6258, 260.5505, 260.5927, 260.6169, 260.7104, 260.731, 260.7501, 
    260.7877, 260.836, 260.9207, 260.9944, 261.0618, 261.0569, 261.0586, 
    261.0736, 261.0364, 261.0797, 261.087, 261.068, 261.1784, 261.1469, 
    261.1791, 261.1586, 260.6423, 260.6679, 260.654, 260.68, 260.6617, 
    260.7432, 260.7676, 260.8819, 260.8351, 260.9097, 260.8427, 260.8545, 
    260.9121, 260.8463, 260.9904, 260.8926, 261.0742, 260.9765, 261.0803, 
    261.0615, 261.0927, 261.1206, 261.1557, 261.2205, 261.2055, 261.2596, 
    260.7061, 260.7392, 260.7363, 260.7711, 260.7968, 260.8525, 260.9418, 
    260.9082, 260.9699, 260.9823, 260.8886, 260.9461, 260.7614, 260.7913, 
    260.7735, 260.7086, 260.9159, 260.8095, 261.006, 260.9484, 261.1166, 
    261.0329, 261.1972, 261.2673, 261.3335, 261.4106, 260.7574, 260.7348, 
    260.7752, 260.8311, 260.883, 260.9519, 260.959, 260.9719, 261.0054, 
    261.0335, 260.976, 261.0405, 260.7981, 260.9252, 260.7263, 260.7861, 
    260.8278, 260.8095, 260.9044, 260.9268, 261.0175, 260.9706, 261.25, 
    261.1264, 261.4694, 261.3736, 260.7269, 260.7573, 260.863, 260.8127, 
    260.9565, 260.9919, 261.0207, 261.0575, 261.0615, 261.0833, 261.0475, 
    261.0818, 260.9521, 261.0101, 260.8509, 260.8896, 260.8719, 260.8523, 
    260.9126, 260.9768, 260.9783, 260.9988, 261.0567, 260.9571, 261.2658, 
    261.0751, 260.7904, 260.8488, 260.8573, 260.8346, 260.9884, 260.9326, 
    261.0827, 261.0422, 261.1086, 261.0756, 261.0707, 261.0284, 261.0019, 
    260.9352, 260.8809, 260.8379, 260.8479, 260.8952, 260.9808, 261.0618, 
    261.044, 261.1036, 260.9461, 261.0121, 260.9866, 261.0532, 260.9073, 
    261.0313, 260.8756, 260.8893, 260.9315, 261.0165, 261.0354, 261.0555, 
    261.0431, 260.983, 260.9731, 260.9305, 260.9188, 260.8863, 260.8594, 
    260.884, 260.9098, 260.983, 261.049, 261.1209, 261.1386, 261.2225, 
    261.1541, 261.2669, 261.1709, 261.3371, 261.0386, 261.1682, 260.9335, 
    260.9588, 261.0045, 261.1094, 261.0528, 261.119, 260.9727, 260.8968, 
    260.8772, 260.8405, 260.878, 260.875, 260.9109, 260.8993, 260.9854, 
    260.9392, 261.0706, 261.1185, 261.2539, 261.3369, 261.4214, 261.4587, 
    261.4701, 261.4748 ;

 FIRE_R =
  260.562, 260.6387, 260.6238, 260.6855, 260.6513, 260.6917, 260.5776, 
    260.6417, 260.6008, 260.569, 260.8053, 260.6883, 260.9271, 260.8524, 
    261.0401, 260.9155, 261.0652, 261.0365, 261.123, 261.0982, 261.2086, 
    261.1344, 261.266, 261.1909, 261.2026, 261.1319, 260.7119, 260.7907, 
    260.7072, 260.7185, 260.7134, 260.652, 260.621, 260.5562, 260.568, 
    260.6156, 260.7235, 260.6869, 260.7793, 260.7772, 260.88, 260.8336, 
    261.0064, 260.9573, 261.0992, 261.0635, 261.0976, 261.0872, 261.0977, 
    261.0453, 261.0678, 261.0217, 260.8423, 260.895, 260.7378, 260.6431, 
    260.5804, 260.5359, 260.5421, 260.5541, 260.6158, 260.6739, 260.7182, 
    260.7477, 260.7769, 260.865, 260.9117, 261.0163, 260.9975, 261.0294, 
    261.06, 261.1113, 261.1028, 261.1254, 261.0286, 261.0929, 260.9868, 
    261.0158, 260.7846, 260.6968, 260.6593, 260.6266, 260.547, 260.602, 
    260.5803, 260.6319, 260.6647, 260.6485, 260.7486, 260.7097, 260.9145, 
    260.8263, 261.0564, 261.0014, 261.0696, 261.0348, 261.0945, 261.0408, 
    261.1338, 261.1541, 261.1402, 261.1934, 261.0378, 261.0975, 260.648, 
    260.6507, 260.663, 260.6088, 260.6055, 260.5559, 260.6, 260.6188, 
    260.6666, 260.6948, 260.7217, 260.7807, 260.8466, 260.9387, 261.0049, 
    261.0493, 261.0221, 261.0461, 261.0193, 261.0067, 261.1465, 261.068, 
    261.1858, 261.1792, 261.1259, 261.18, 260.6525, 260.6373, 260.5845, 
    260.6258, 260.5505, 260.5927, 260.6169, 260.7104, 260.731, 260.7501, 
    260.7877, 260.836, 260.9207, 260.9944, 261.0618, 261.0569, 261.0586, 
    261.0736, 261.0364, 261.0797, 261.087, 261.068, 261.1784, 261.1469, 
    261.1791, 261.1586, 260.6423, 260.6679, 260.654, 260.68, 260.6617, 
    260.7432, 260.7676, 260.8819, 260.8351, 260.9097, 260.8427, 260.8545, 
    260.9121, 260.8463, 260.9904, 260.8926, 261.0742, 260.9765, 261.0803, 
    261.0615, 261.0927, 261.1206, 261.1557, 261.2205, 261.2055, 261.2596, 
    260.7061, 260.7392, 260.7363, 260.7711, 260.7968, 260.8525, 260.9418, 
    260.9082, 260.9699, 260.9823, 260.8886, 260.9461, 260.7614, 260.7913, 
    260.7735, 260.7086, 260.9159, 260.8095, 261.006, 260.9484, 261.1166, 
    261.0329, 261.1972, 261.2673, 261.3335, 261.4106, 260.7574, 260.7348, 
    260.7752, 260.8311, 260.883, 260.9519, 260.959, 260.9719, 261.0054, 
    261.0335, 260.976, 261.0405, 260.7981, 260.9252, 260.7263, 260.7861, 
    260.8278, 260.8095, 260.9044, 260.9268, 261.0175, 260.9706, 261.25, 
    261.1264, 261.4694, 261.3736, 260.7269, 260.7573, 260.863, 260.8127, 
    260.9565, 260.9919, 261.0207, 261.0575, 261.0615, 261.0833, 261.0475, 
    261.0818, 260.9521, 261.0101, 260.8509, 260.8896, 260.8719, 260.8523, 
    260.9126, 260.9768, 260.9783, 260.9988, 261.0567, 260.9571, 261.2658, 
    261.0751, 260.7904, 260.8488, 260.8573, 260.8346, 260.9884, 260.9326, 
    261.0827, 261.0422, 261.1086, 261.0756, 261.0707, 261.0284, 261.0019, 
    260.9352, 260.8809, 260.8379, 260.8479, 260.8952, 260.9808, 261.0618, 
    261.044, 261.1036, 260.9461, 261.0121, 260.9866, 261.0532, 260.9073, 
    261.0313, 260.8756, 260.8893, 260.9315, 261.0165, 261.0354, 261.0555, 
    261.0431, 260.983, 260.9731, 260.9305, 260.9188, 260.8863, 260.8594, 
    260.884, 260.9098, 260.983, 261.049, 261.1209, 261.1386, 261.2225, 
    261.1541, 261.2669, 261.1709, 261.3371, 261.0386, 261.1682, 260.9335, 
    260.9588, 261.0045, 261.1094, 261.0528, 261.119, 260.9727, 260.8968, 
    260.8772, 260.8405, 260.878, 260.875, 260.9109, 260.8993, 260.9854, 
    260.9392, 261.0706, 261.1185, 261.2539, 261.3369, 261.4214, 261.4587, 
    261.4701, 261.4748 ;

 FIRE_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FLDS =
  214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 214.3461, 
    214.3461, 214.3461 ;

 FPG =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 FPI_vr =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WJ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FPSN_WP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTC_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FROST_TABLE =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 FSA =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 FSAT =
  0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 0.04295584, 
    0.04295584, 0.04295584 ;

 FSA_R =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 FSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSDS =
  1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 1.20347, 
    1.20347, 1.20347 ;

 FSDSND =
  0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 0.1797532, 
    0.1797532, 0.1797532 ;

 FSDSNDLN =
  0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495 ;

 FSDSNI =
  0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 0.4219819, 
    0.4219819, 0.4219819 ;

 FSDSVD =
  0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 0.1076128, 
    0.1076128, 0.1076128 ;

 FSDSVDLN =
  0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609 ;

 FSDSVI =
  0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 0.4941223, 
    0.4941223, 0.4941223 ;

 FSDSVILN =
  0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 0.7227376, 
    0.7227376, 0.7227376 ;

 FSH =
  317.8795, 318.8366, 318.6507, 319.4223, 318.9945, 319.4996, 318.0738, 
    318.8744, 318.3635, 317.966, 320.919, 319.4568, 322.4401, 321.5073, 
    323.8511, 322.2946, 324.1651, 323.8068, 324.8864, 324.5771, 325.9565, 
    325.0291, 326.6723, 325.7354, 325.8817, 324.9984, 319.7516, 320.7368, 
    319.6931, 319.8336, 319.7707, 319.0031, 318.6159, 317.8067, 317.9538, 
    318.5483, 319.8968, 319.4394, 320.5933, 320.5672, 321.8513, 321.2724, 
    323.4308, 322.8175, 324.5901, 324.1443, 324.569, 324.4403, 324.5707, 
    323.9169, 324.197, 323.6218, 321.3807, 322.0392, 320.0747, 318.8926, 
    318.1088, 317.5522, 317.6309, 317.7808, 318.5518, 319.2771, 319.8297, 
    320.1993, 320.5635, 321.6644, 322.2483, 323.5545, 323.3193, 323.7182, 
    324.0999, 324.7401, 324.6348, 324.9167, 323.708, 324.5112, 323.1852, 
    323.5478, 320.6606, 319.5629, 319.0947, 318.6863, 317.6913, 318.3784, 
    318.1075, 318.7523, 319.1618, 318.9594, 320.2094, 319.7233, 322.2829, 
    321.1805, 324.0554, 323.3676, 324.2203, 323.7853, 324.5305, 323.8599, 
    325.0218, 325.2746, 325.1018, 325.7661, 323.8226, 324.5688, 318.9536, 
    318.9866, 319.1406, 318.4637, 318.4224, 317.8026, 318.3542, 318.589, 
    319.1857, 319.5382, 319.8735, 320.6107, 321.4337, 322.5849, 323.4122, 
    323.9666, 323.6268, 323.9268, 323.5913, 323.4342, 325.1797, 324.1995, 
    325.6706, 325.5893, 324.9234, 325.5984, 319.0098, 318.8198, 318.1596, 
    318.6763, 317.7351, 318.2617, 318.5643, 319.7331, 319.9903, 320.2282, 
    320.6986, 321.302, 322.3603, 323.2813, 324.1222, 324.0606, 324.0823, 
    324.27, 323.8049, 324.3463, 324.437, 324.1996, 325.5783, 325.1845, 
    325.5875, 325.3311, 318.8816, 319.2014, 319.0286, 319.3534, 319.1244, 
    320.1422, 320.4474, 321.8757, 321.29, 322.2227, 321.3849, 321.5332, 
    322.2523, 321.4303, 323.2301, 322.0092, 324.2773, 323.0574, 324.3536, 
    324.1186, 324.5079, 324.8564, 325.2952, 326.1041, 325.9168, 326.5935, 
    319.6782, 320.0928, 320.0567, 320.4908, 320.8117, 321.5078, 322.6237, 
    322.2042, 322.9747, 323.1292, 321.9589, 322.6771, 320.3705, 320.7429, 
    320.5215, 319.7107, 322.3004, 320.9712, 323.4258, 322.7059, 324.8067, 
    323.7617, 325.8137, 326.6897, 327.5157, 328.4788, 320.3195, 320.0377, 
    320.5425, 321.2402, 321.8885, 322.7498, 322.8381, 322.9993, 323.4174, 
    323.7687, 323.05, 323.8568, 320.8285, 322.4159, 319.9309, 320.6787, 
    321.1992, 320.9713, 322.1563, 322.4355, 323.5697, 322.9836, 326.4732, 
    324.9295, 329.2132, 328.0163, 319.9392, 320.3187, 321.6387, 321.0107, 
    322.8075, 323.2495, 323.6092, 324.0683, 324.1181, 324.3902, 323.9443, 
    324.3727, 322.7516, 323.4761, 321.4883, 321.9719, 321.7495, 321.5053, 
    322.2589, 323.0612, 323.0789, 323.336, 324.0594, 322.8148, 326.6713, 
    324.2889, 320.7324, 321.4624, 321.5674, 321.2845, 323.2052, 322.5092, 
    324.3836, 323.8772, 324.7071, 324.2947, 324.234, 323.7044, 323.3745, 
    322.541, 321.863, 321.3256, 321.4506, 322.0409, 323.1104, 324.1224, 
    323.9006, 324.644, 322.6772, 323.5017, 323.1828, 324.0143, 322.1929, 
    323.7422, 321.7967, 321.9674, 322.4954, 323.5572, 323.793, 324.0436, 
    323.8891, 323.1376, 323.0148, 322.4827, 322.3355, 321.9303, 321.5945, 
    321.9011, 322.2231, 323.1382, 323.9625, 324.8613, 325.0815, 326.1299, 
    325.2756, 326.6844, 325.4855, 327.5613, 323.8328, 325.4514, 322.5196, 
    322.8357, 323.4067, 324.7173, 324.0104, 324.8374, 323.01, 322.061, 
    321.8162, 321.3582, 321.8266, 321.7886, 322.2368, 322.0928, 323.1686, 
    322.5908, 324.2323, 324.8311, 326.5224, 327.5585, 328.6139, 329.0795, 
    329.2212, 329.2804 ;

 FSH_G =
  324.5388, 325.4964, 325.3104, 326.0825, 325.6544, 326.1598, 324.7332, 
    325.5342, 325.023, 324.6253, 327.58, 326.117, 329.102, 328.1687, 
    330.5138, 328.9565, 330.8279, 330.4695, 331.5497, 331.2403, 332.6204, 
    331.6925, 333.3366, 332.3991, 332.5456, 331.6617, 326.412, 327.3977, 
    326.3534, 326.494, 326.4311, 325.663, 325.2756, 324.466, 324.6131, 
    325.2079, 326.5573, 326.0996, 327.2541, 327.2281, 328.5129, 327.9336, 
    330.0933, 329.4796, 331.2532, 330.8071, 331.2321, 331.1034, 331.2338, 
    330.5796, 330.8599, 330.2844, 328.042, 328.7009, 326.7353, 325.5525, 
    324.7682, 324.2113, 324.29, 324.44, 325.2114, 325.9372, 326.4901, 
    326.8599, 327.2243, 328.3258, 328.91, 330.2171, 329.9817, 330.3808, 
    330.7628, 331.4034, 331.298, 331.5801, 330.3706, 331.1743, 329.8475, 
    330.2104, 327.3214, 326.2232, 325.7547, 325.3461, 324.3505, 325.0379, 
    324.7669, 325.4121, 325.8218, 325.6193, 326.87, 326.3837, 328.9446, 
    327.8416, 330.7182, 330.0301, 330.8832, 330.448, 331.1936, 330.5226, 
    331.6852, 331.9381, 331.7653, 332.4299, 330.4853, 331.232, 325.6135, 
    325.6465, 325.8006, 325.1233, 325.0819, 324.4619, 325.0138, 325.2487, 
    325.8457, 326.1985, 326.5339, 327.2715, 328.095, 329.2469, 330.0746, 
    330.6294, 330.2893, 330.5895, 330.2539, 330.0966, 331.8432, 330.8624, 
    332.3343, 332.253, 331.5867, 332.2621, 325.6697, 325.4796, 324.819, 
    325.336, 324.3943, 324.9212, 325.224, 326.3934, 326.6508, 326.8889, 
    327.3595, 327.9632, 329.0221, 329.9436, 330.7851, 330.7235, 330.7451, 
    330.9329, 330.4675, 331.0093, 331.1, 330.8625, 332.2421, 331.848, 
    332.2512, 331.9947, 325.5415, 325.8614, 325.6885, 326.0135, 325.7844, 
    326.8028, 327.1081, 328.5373, 327.9512, 328.8844, 328.0462, 328.1946, 
    328.914, 328.0916, 329.8925, 328.6708, 330.9402, 329.7197, 331.0166, 
    330.7814, 331.171, 331.5197, 331.9587, 332.7681, 332.5807, 333.2578, 
    326.3385, 326.7534, 326.7172, 327.1516, 327.4727, 328.1692, 329.2857, 
    328.866, 329.6369, 329.7915, 328.6205, 329.3391, 327.0312, 327.4037, 
    327.1822, 326.3711, 328.9622, 327.6322, 330.0883, 329.368, 331.4699, 
    330.4243, 332.4775, 333.354, 334.1805, 335.1442, 326.9801, 326.6982, 
    327.2033, 327.9014, 328.5501, 329.4118, 329.5002, 329.6615, 330.0799, 
    330.4314, 329.7122, 330.5195, 327.4894, 329.0778, 326.5913, 327.3396, 
    327.8604, 327.6323, 328.8181, 329.0974, 330.2322, 329.6458, 333.1374, 
    331.5928, 335.879, 334.6814, 326.5997, 326.9793, 328.3001, 327.6718, 
    329.4696, 329.9119, 330.2717, 330.7311, 330.781, 331.0532, 330.6071, 
    331.0357, 329.4137, 330.1386, 328.1496, 328.6335, 328.411, 328.1667, 
    328.9207, 329.7234, 329.7411, 329.9984, 330.7222, 329.4769, 333.3356, 
    330.9518, 327.3933, 328.1237, 328.2288, 327.9457, 329.8675, 329.1711, 
    331.0467, 330.5399, 331.3703, 330.9576, 330.8969, 330.367, 330.0369, 
    329.203, 328.5245, 327.9868, 328.1119, 328.7026, 329.7726, 330.7852, 
    330.5634, 331.3072, 329.3392, 330.1642, 329.8452, 330.6771, 328.8547, 
    330.4048, 328.4582, 328.629, 329.1573, 330.2197, 330.4557, 330.7065, 
    330.5518, 329.7999, 329.677, 329.1446, 328.9973, 328.5919, 328.2559, 
    328.5627, 328.8848, 329.8005, 330.6253, 331.5246, 331.7449, 332.7939, 
    331.9391, 333.3488, 332.1491, 334.2262, 330.4955, 332.115, 329.1816, 
    329.4978, 330.0691, 331.3805, 330.6732, 331.5007, 329.6722, 328.7227, 
    328.4777, 328.0194, 328.4882, 328.4501, 328.8986, 328.7545, 329.8309, 
    329.2527, 330.8952, 331.4943, 333.1866, 334.2234, 335.2794, 335.7452, 
    335.887, 335.9463 ;

 FSH_NODYNLNDUSE =
  317.8795, 318.8366, 318.6507, 319.4223, 318.9945, 319.4996, 318.0738, 
    318.8744, 318.3635, 317.966, 320.919, 319.4568, 322.4401, 321.5073, 
    323.8511, 322.2946, 324.1651, 323.8068, 324.8864, 324.5771, 325.9565, 
    325.0291, 326.6723, 325.7354, 325.8817, 324.9984, 319.7516, 320.7368, 
    319.6931, 319.8336, 319.7707, 319.0031, 318.6159, 317.8067, 317.9538, 
    318.5483, 319.8968, 319.4394, 320.5933, 320.5672, 321.8513, 321.2724, 
    323.4308, 322.8175, 324.5901, 324.1443, 324.569, 324.4403, 324.5707, 
    323.9169, 324.197, 323.6218, 321.3807, 322.0392, 320.0747, 318.8926, 
    318.1088, 317.5522, 317.6309, 317.7808, 318.5518, 319.2771, 319.8297, 
    320.1993, 320.5635, 321.6644, 322.2483, 323.5545, 323.3193, 323.7182, 
    324.0999, 324.7401, 324.6348, 324.9167, 323.708, 324.5112, 323.1852, 
    323.5478, 320.6606, 319.5629, 319.0947, 318.6863, 317.6913, 318.3784, 
    318.1075, 318.7523, 319.1618, 318.9594, 320.2094, 319.7233, 322.2829, 
    321.1805, 324.0554, 323.3676, 324.2203, 323.7853, 324.5305, 323.8599, 
    325.0218, 325.2746, 325.1018, 325.7661, 323.8226, 324.5688, 318.9536, 
    318.9866, 319.1406, 318.4637, 318.4224, 317.8026, 318.3542, 318.589, 
    319.1857, 319.5382, 319.8735, 320.6107, 321.4337, 322.5849, 323.4122, 
    323.9666, 323.6268, 323.9268, 323.5913, 323.4342, 325.1797, 324.1995, 
    325.6706, 325.5893, 324.9234, 325.5984, 319.0098, 318.8198, 318.1596, 
    318.6763, 317.7351, 318.2617, 318.5643, 319.7331, 319.9903, 320.2282, 
    320.6986, 321.302, 322.3603, 323.2813, 324.1222, 324.0606, 324.0823, 
    324.27, 323.8049, 324.3463, 324.437, 324.1996, 325.5783, 325.1845, 
    325.5875, 325.3311, 318.8816, 319.2014, 319.0286, 319.3534, 319.1244, 
    320.1422, 320.4474, 321.8757, 321.29, 322.2227, 321.3849, 321.5332, 
    322.2523, 321.4303, 323.2301, 322.0092, 324.2773, 323.0574, 324.3536, 
    324.1186, 324.5079, 324.8564, 325.2952, 326.1041, 325.9168, 326.5935, 
    319.6782, 320.0928, 320.0567, 320.4908, 320.8117, 321.5078, 322.6237, 
    322.2042, 322.9747, 323.1292, 321.9589, 322.6771, 320.3705, 320.7429, 
    320.5215, 319.7107, 322.3004, 320.9712, 323.4258, 322.7059, 324.8067, 
    323.7617, 325.8137, 326.6897, 327.5157, 328.4788, 320.3195, 320.0377, 
    320.5425, 321.2402, 321.8885, 322.7498, 322.8381, 322.9993, 323.4174, 
    323.7687, 323.05, 323.8568, 320.8285, 322.4159, 319.9309, 320.6787, 
    321.1992, 320.9713, 322.1563, 322.4355, 323.5697, 322.9836, 326.4732, 
    324.9295, 329.2132, 328.0163, 319.9392, 320.3187, 321.6387, 321.0107, 
    322.8075, 323.2495, 323.6092, 324.0683, 324.1181, 324.3902, 323.9443, 
    324.3727, 322.7516, 323.4761, 321.4883, 321.9719, 321.7495, 321.5053, 
    322.2589, 323.0612, 323.0789, 323.336, 324.0594, 322.8148, 326.6713, 
    324.2889, 320.7324, 321.4624, 321.5674, 321.2845, 323.2052, 322.5092, 
    324.3836, 323.8772, 324.7071, 324.2947, 324.234, 323.7044, 323.3745, 
    322.541, 321.863, 321.3256, 321.4506, 322.0409, 323.1104, 324.1224, 
    323.9006, 324.644, 322.6772, 323.5017, 323.1828, 324.0143, 322.1929, 
    323.7422, 321.7967, 321.9674, 322.4954, 323.5572, 323.793, 324.0436, 
    323.8891, 323.1376, 323.0148, 322.4827, 322.3355, 321.9303, 321.5945, 
    321.9011, 322.2231, 323.1382, 323.9625, 324.8613, 325.0815, 326.1299, 
    325.2756, 326.6844, 325.4855, 327.5613, 323.8328, 325.4514, 322.5196, 
    322.8357, 323.4067, 324.7173, 324.0104, 324.8374, 323.01, 322.061, 
    321.8162, 321.3582, 321.8266, 321.7886, 322.2368, 322.0928, 323.1686, 
    322.5908, 324.2323, 324.8311, 326.5224, 327.5585, 328.6139, 329.0795, 
    329.2212, 329.2804 ;

 FSH_R =
  317.8795, 318.8366, 318.6507, 319.4223, 318.9945, 319.4996, 318.0738, 
    318.8744, 318.3635, 317.966, 320.919, 319.4568, 322.4401, 321.5073, 
    323.8511, 322.2946, 324.1651, 323.8068, 324.8864, 324.5771, 325.9565, 
    325.0291, 326.6723, 325.7354, 325.8817, 324.9984, 319.7516, 320.7368, 
    319.6931, 319.8336, 319.7707, 319.0031, 318.6159, 317.8067, 317.9538, 
    318.5483, 319.8968, 319.4394, 320.5933, 320.5672, 321.8513, 321.2724, 
    323.4308, 322.8175, 324.5901, 324.1443, 324.569, 324.4403, 324.5707, 
    323.9169, 324.197, 323.6218, 321.3807, 322.0392, 320.0747, 318.8926, 
    318.1088, 317.5522, 317.6309, 317.7808, 318.5518, 319.2771, 319.8297, 
    320.1993, 320.5635, 321.6644, 322.2483, 323.5545, 323.3193, 323.7182, 
    324.0999, 324.7401, 324.6348, 324.9167, 323.708, 324.5112, 323.1852, 
    323.5478, 320.6606, 319.5629, 319.0947, 318.6863, 317.6913, 318.3784, 
    318.1075, 318.7523, 319.1618, 318.9594, 320.2094, 319.7233, 322.2829, 
    321.1805, 324.0554, 323.3676, 324.2203, 323.7853, 324.5305, 323.8599, 
    325.0218, 325.2746, 325.1018, 325.7661, 323.8226, 324.5688, 318.9536, 
    318.9866, 319.1406, 318.4637, 318.4224, 317.8026, 318.3542, 318.589, 
    319.1857, 319.5382, 319.8735, 320.6107, 321.4337, 322.5849, 323.4122, 
    323.9666, 323.6268, 323.9268, 323.5913, 323.4342, 325.1797, 324.1995, 
    325.6706, 325.5893, 324.9234, 325.5984, 319.0098, 318.8198, 318.1596, 
    318.6763, 317.7351, 318.2617, 318.5643, 319.7331, 319.9903, 320.2282, 
    320.6986, 321.302, 322.3603, 323.2813, 324.1222, 324.0606, 324.0823, 
    324.27, 323.8049, 324.3463, 324.437, 324.1996, 325.5783, 325.1845, 
    325.5875, 325.3311, 318.8816, 319.2014, 319.0286, 319.3534, 319.1244, 
    320.1422, 320.4474, 321.8757, 321.29, 322.2227, 321.3849, 321.5332, 
    322.2523, 321.4303, 323.2301, 322.0092, 324.2773, 323.0574, 324.3536, 
    324.1186, 324.5079, 324.8564, 325.2952, 326.1041, 325.9168, 326.5935, 
    319.6782, 320.0928, 320.0567, 320.4908, 320.8117, 321.5078, 322.6237, 
    322.2042, 322.9747, 323.1292, 321.9589, 322.6771, 320.3705, 320.7429, 
    320.5215, 319.7107, 322.3004, 320.9712, 323.4258, 322.7059, 324.8067, 
    323.7617, 325.8137, 326.6897, 327.5157, 328.4788, 320.3195, 320.0377, 
    320.5425, 321.2402, 321.8885, 322.7498, 322.8381, 322.9993, 323.4174, 
    323.7687, 323.05, 323.8568, 320.8285, 322.4159, 319.9309, 320.6787, 
    321.1992, 320.9713, 322.1563, 322.4355, 323.5697, 322.9836, 326.4732, 
    324.9295, 329.2132, 328.0163, 319.9392, 320.3187, 321.6387, 321.0107, 
    322.8075, 323.2495, 323.6092, 324.0683, 324.1181, 324.3902, 323.9443, 
    324.3727, 322.7516, 323.4761, 321.4883, 321.9719, 321.7495, 321.5053, 
    322.2589, 323.0612, 323.0789, 323.336, 324.0594, 322.8148, 326.6713, 
    324.2889, 320.7324, 321.4624, 321.5674, 321.2845, 323.2052, 322.5092, 
    324.3836, 323.8772, 324.7071, 324.2947, 324.234, 323.7044, 323.3745, 
    322.541, 321.863, 321.3256, 321.4506, 322.0409, 323.1104, 324.1224, 
    323.9006, 324.644, 322.6772, 323.5017, 323.1828, 324.0143, 322.1929, 
    323.7422, 321.7967, 321.9674, 322.4954, 323.5572, 323.793, 324.0436, 
    323.8891, 323.1376, 323.0148, 322.4827, 322.3355, 321.9303, 321.5945, 
    321.9011, 322.2231, 323.1382, 323.9625, 324.8613, 325.0815, 326.1299, 
    325.2756, 326.6844, 325.4855, 327.5613, 323.8328, 325.4514, 322.5196, 
    322.8357, 323.4067, 324.7173, 324.0104, 324.8374, 323.01, 322.061, 
    321.8162, 321.3582, 321.8266, 321.7886, 322.2368, 322.0928, 323.1686, 
    322.5908, 324.2323, 324.8311, 326.5224, 327.5585, 328.6139, 329.0795, 
    329.2212, 329.2804 ;

 FSH_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSH_V =
  -6.659277, -6.659824, -6.659721, -6.660156, -6.659919, -6.660201, 
    -6.659393, -6.659842, -6.659558, -6.659333, -6.660989, -6.660177, 
    -6.66188, -6.661354, -6.662693, -6.661792, -6.662877, -6.662678, 
    -6.663304, -6.663125, -6.663904, -6.663386, -6.664327, -6.663786, 
    -6.663867, -6.663368, -6.660351, -6.660884, -6.660317, -6.660393, 
    -6.660361, -6.65992, -6.65969, -6.659243, -6.659327, -6.659659, 
    -6.660428, -6.660174, -6.660836, -6.660821, -6.661552, -6.661222, 
    -6.662461, -6.662111, -6.663133, -6.662874, -6.663118, -6.663046, 
    -6.663119, -6.66274, -6.662902, -6.662572, -6.661282, -6.661657, 
    -6.660533, -6.659842, -6.659411, -6.659097, -6.659142, -6.659224, 
    -6.65966, -6.660081, -6.660398, -6.66061, -6.660819, -6.661425, -6.66177, 
    -6.662526, -6.662399, -6.662622, -6.662848, -6.663216, -6.663157, 
    -6.663317, -6.662623, -6.663081, -6.662324, -6.66253, -6.660839, 
    -6.660244, -6.65996, -6.659739, -6.659174, -6.659563, -6.659409, 
    -6.659782, -6.660015, -6.659902, -6.660615, -6.660336, -6.66179, 
    -6.661164, -6.662822, -6.662426, -6.662918, -6.662669, -6.663094, 
    -6.662711, -6.66338, -6.663521, -6.663424, -6.663811, -6.662689, 
    -6.663115, -6.659896, -6.659914, -6.660004, -6.65961, -6.659588, 
    -6.659239, -6.659553, -6.659684, -6.660031, -6.66023, -6.660421, 
    -6.660842, -6.661307, -6.661969, -6.662451, -6.662773, -6.662578, 
    -6.66275, -6.662556, -6.662467, -6.663465, -6.662901, -6.663755, 
    -6.663709, -6.66332, -6.663714, -6.659928, -6.659822, -6.659441, 
    -6.659739, -6.659202, -6.659498, -6.659666, -6.660334, -6.66049, 
    -6.660623, -6.660894, -6.661239, -6.661841, -6.662372, -6.662863, 
    -6.662828, -6.66284, -6.662946, -6.662678, -6.66299, -6.663039, 
    -6.662906, -6.663702, -6.663475, -6.663708, -6.663561, -6.659857, 
    -6.660038, -6.65994, -6.660122, -6.659991, -6.660566, -6.660738, 
    -6.661557, -6.66123, -6.66176, -6.661287, -6.661368, -6.661762, 
    -6.661314, -6.662336, -6.661629, -6.66295, -6.662228, -6.662994, 
    -6.662861, -6.663085, -6.663283, -6.663538, -6.664, -6.663894, -6.664287, 
    -6.660311, -6.660542, -6.660529, -6.660776, -6.660957, -6.661358, 
    -6.661995, -6.661758, -6.662202, -6.662289, -6.661619, -6.662023, 
    -6.660702, -6.660908, -6.66079, -6.660325, -6.661803, -6.661039, 
    -6.662458, -6.662045, -6.663254, -6.662645, -6.663835, -6.664327, 
    -6.664824, -6.665367, -6.660676, -6.660518, -6.660807, -6.661194, 
    -6.661574, -6.662068, -6.662123, -6.662213, -6.662457, -6.662659, 
    -6.662235, -6.66271, -6.660942, -6.661873, -6.660452, -6.66087, 
    -6.661175, -6.661048, -6.661733, -6.661892, -6.662537, -6.662207, 
    -6.664199, -6.663315, -6.665804, -6.665102, -6.660461, -6.660678, 
    -6.661427, -6.661071, -6.662105, -6.662357, -6.662568, -6.662827, 
    -6.662859, -6.663014, -6.66276, -6.663006, -6.662069, -6.662489, 
    -6.661349, -6.661622, -6.661499, -6.661358, -6.661791, -6.662241, 
    -6.662261, -6.662404, -6.662785, -6.662109, -6.664293, -6.662923, 
    -6.660915, -6.661319, -6.661391, -6.661232, -6.662331, -6.661931, 
    -6.663012, -6.662722, -6.6632, -6.662961, -6.662925, -6.662621, -6.66243, 
    -6.661947, -6.661558, -6.661256, -6.661327, -6.66166, -6.662271, 
    -6.662858, -6.662727, -6.663164, -6.66203, -6.662499, -6.662313, 
    -6.662798, -6.661749, -6.662609, -6.661526, -6.661623, -6.661923, 
    -6.662523, -6.662673, -6.662812, -6.662728, -6.662288, -6.662221, 
    -6.661919, -6.661829, -6.661603, -6.66141, -6.661583, -6.661763, 
    -6.662293, -6.662765, -6.663284, -6.663416, -6.663996, -6.663508, 
    -6.664298, -6.663603, -6.664819, -6.662675, -6.663605, -6.661941, 
    -6.662122, -6.662439, -6.663191, -6.662796, -6.663263, -6.66222, 
    -6.661665, -6.661536, -6.661273, -6.661542, -6.661521, -6.661778, 
    -6.661696, -6.662311, -6.661981, -6.662921, -6.663262, -6.664241, 
    -6.664836, -6.665461, -6.665731, -6.665814, -6.665849 ;

 FSM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSM_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 FSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSNO_EFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 FSR =
  1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 1.151179, 
    1.151179, 1.151179 ;

 FSRND =
  0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 0.1719234, 
    0.1719234, 0.1719234 ;

 FSRNDLN =
  0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 0.2642495, 
    0.2642495, 0.2642495 ;

 FSRNI =
  0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 0.403666, 
    0.403666, 0.403666 ;

 FSRVD =
  0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 0.1029223, 
    0.1029223, 0.1029223 ;

 FSRVDLN =
  0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 0.1583609, 
    0.1583609, 0.1583609 ;

 FSRVI =
  0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 0.4726671, 
    0.4726671, 0.4726671 ;

 FUELC =
  0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 0.8953806, 
    0.8953806, 0.8953806 ;

 F_DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.605194e-45, 0, 4.551417e-42, 
    2.802597e-45, 1.913193e-41, 3.698027e-42, 4.768479e-40, 1.216804e-40, 
    4.618803e-38, 8.893803e-40, 8.562508e-37, 1.82806e-38, 3.377825e-38, 
    7.783162e-40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.403934e-43, 3.363116e-44, 1.288718e-40, 1.736209e-41, 1.174148e-40, 
    6.60418e-41, 1.182948e-40, 6.143292e-42, 2.207185e-41, 1.56525e-42, 0, 
    1.401298e-45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 
    1.146262e-42, 3.783506e-43, 2.455075e-42, 1.418815e-41, 2.508002e-40, 
    1.572887e-40, 5.453685e-40, 2.337366e-42, 9.083777e-41, 1.989844e-43, 
    1.108427e-42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.802597e-45, 0, 
    1.158313e-41, 4.750402e-43, 2.451432e-41, 3.343498e-42, 9.89597e-41, 
    4.718172e-42, 8.623619e-40, 2.577666e-39, 1.221582e-39, 2.076547e-38, 
    3.974082e-42, 1.174288e-40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.121039e-44, 5.857428e-43, 7.708543e-42, 1.600283e-42, 6.42075e-42, 
    1.356457e-42, 6.488012e-43, 1.713117e-39, 2.23367e-41, 1.389566e-38, 
    9.852799e-39, 5.616474e-40, 1.024267e-38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4.203895e-45, 3.152922e-43, 1.569594e-41, 1.185358e-41, 
    1.308673e-41, 3.069544e-41, 3.661593e-42, 4.331554e-41, 6.516038e-41, 
    2.232128e-41, 9.408437e-39, 1.745448e-39, 9.780899e-39, 3.279918e-39, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 0, 0, 2.802597e-45, 0, 
    2.480298e-43, 0, 3.1724e-41, 1.093013e-43, 4.476448e-41, 1.543811e-41, 
    8.93538e-41, 4.185454e-40, 2.811773e-39, 8.485865e-38, 3.902624e-38, 
    6.231172e-37, 0, 0, 0, 0, 0, 0, 1.261169e-44, 1.401298e-45, 7.286752e-44, 
    1.527415e-43, 0, 1.681558e-44, 0, 0, 0, 0, 2.802597e-45, 0, 6.249791e-43, 
    1.961818e-44, 3.363915e-40, 3.005785e-42, 2.536987e-38, 9.203849e-37, 
    2.340174e-35, 8.675964e-34, 0, 0, 0, 0, 0, 2.522337e-44, 3.783506e-44, 
    8.267661e-44, 5.997557e-43, 3.09687e-42, 1.050974e-43, 4.652311e-42, 0, 
    4.203895e-45, 0, 0, 0, 0, 1.401298e-45, 5.605194e-45, 1.228939e-42, 
    7.567012e-44, 3.850611e-37, 5.781982e-40, 1.20543e-32, 1.566253e-34, 0, 
    0, 0, 0, 3.222986e-44, 2.718519e-43, 1.474166e-42, 1.229499e-41, 
    1.541148e-41, 5.278831e-41, 6.960249e-42, 4.876519e-41, 2.522337e-44, 
    7.917336e-43, 0, 0, 0, 0, 2.802597e-45, 1.107026e-43, 1.205117e-43, 
    4.091792e-43, 1.193206e-41, 3.363116e-44, 8.600233e-37, 3.375868e-41, 0, 
    0, 0, 0, 2.200039e-43, 7.006492e-45, 5.123568e-41, 5.111937e-42, 
    2.165973e-40, 3.4315e-41, 2.608517e-41, 2.298129e-42, 4.904545e-43, 
    8.407791e-45, 0, 0, 0, 1.401298e-45, 1.401298e-43, 1.573378e-41, 
    5.706087e-42, 1.638048e-40, 1.681558e-44, 8.940284e-43, 1.975831e-43, 
    9.598894e-42, 1.401298e-45, 2.766163e-42, 0, 0, 7.006492e-45, 
    1.161676e-42, 3.465411e-42, 1.098618e-41, 5.399203e-42, 1.59748e-43, 
    8.82818e-44, 7.006492e-45, 2.802597e-45, 0, 0, 0, 1.401298e-45, 
    1.59748e-43, 7.578222e-42, 4.277912e-40, 1.117072e-39, 9.486179e-38, 
    2.598732e-39, 9.070593e-37, 6.421963e-39, 2.808711e-35, 4.191284e-42, 
    5.521899e-39, 8.407791e-45, 3.783506e-44, 5.717298e-43, 2.275709e-40, 
    9.427936e-42, 3.860339e-40, 8.68805e-44, 1.401298e-45, 0, 0, 0, 0, 
    1.401298e-45, 1.401298e-45, 1.849714e-43, 1.121039e-44, 2.590861e-41, 
    3.750631e-40, 4.682267e-37, 2.766208e-35, 1.414291e-33, 7.510774e-33, 
    1.238513e-32, 1.524886e-32 ;

 F_DENIT_vr =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.344025e-44, 0, 3.682192e-41, 
    2.101948e-44, 1.54793e-40, 2.991492e-41, 3.857985e-39, 9.84464e-40, 
    3.736885e-37, 7.195609e-39, 6.927575e-36, 1.479009e-37, 2.73286e-37, 
    6.297036e-39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.802597e-45, 0, 
    5.176397e-42, 2.760558e-43, 1.042645e-39, 1.404676e-40, 9.499542e-40, 
    5.343207e-40, 9.570784e-40, 4.969845e-41, 1.785731e-40, 1.266634e-41, 0, 
    5.605194e-45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 
    1.681558e-44, 9.268188e-42, 3.056232e-42, 1.986761e-41, 1.147916e-40, 
    2.029124e-39, 1.27256e-39, 4.412358e-39, 1.891333e-41, 7.349306e-40, 
    1.614296e-42, 8.962705e-42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.961818e-44, 0, 9.371043e-41, 3.840959e-42, 1.983314e-40, 2.705487e-41, 
    8.006403e-40, 3.817838e-41, 6.977017e-39, 2.085484e-38, 9.883324e-39, 
    1.680049e-37, 3.2157e-41, 9.500734e-40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8.82818e-44, 4.740593e-42, 6.236899e-41, 1.29508e-41, 5.195174e-41, 
    1.098057e-41, 5.252067e-42, 1.386012e-38, 1.807171e-40, 1.124241e-37, 
    7.971497e-38, 4.544063e-39, 8.286928e-38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2.942727e-44, 2.555968e-42, 1.269885e-40, 9.590206e-41, 
    1.058765e-40, 2.483451e-40, 2.962905e-41, 3.504493e-40, 5.271867e-40, 
    1.805909e-40, 7.611982e-38, 1.41217e-38, 7.913326e-38, 2.653648e-38, 0, 
    0, 0, 0, 0, 0, 0, 2.802597e-45, 0, 1.541428e-44, 0, 0, 1.681558e-44, 0, 
    2.008061e-42, 5.605194e-45, 2.566702e-40, 8.82818e-43, 3.621684e-40, 
    1.249047e-40, 7.229229e-40, 3.386277e-39, 2.27489e-38, 6.865567e-37, 
    3.157454e-37, 5.041387e-36, 0, 0, 0, 0, 0, 0, 1.079e-43, 1.401298e-44, 
    5.899467e-43, 1.237347e-42, 4.203895e-45, 1.401298e-43, 0, 0, 0, 0, 
    2.242078e-44, 0, 5.055885e-42, 1.59748e-43, 2.721612e-39, 2.432094e-41, 
    2.052572e-37, 7.446458e-36, 1.893339e-34, 7.019368e-33, 0, 0, 0, 0, 
    2.802597e-45, 1.989844e-43, 3.054831e-43, 6.642155e-43, 4.854098e-42, 
    2.505662e-41, 8.491869e-43, 3.764308e-41, 0, 3.923636e-44, 0, 0, 0, 0, 
    1.121039e-44, 4.203895e-44, 9.943614e-42, 6.1517e-43, 3.115371e-36, 
    4.677963e-39, 9.75264e-32, 1.267191e-33, 0, 0, 1.401298e-45, 0, 
    2.620428e-43, 2.195835e-42, 1.192925e-41, 9.947538e-41, 1.246903e-40, 
    4.270905e-40, 5.630978e-41, 3.945342e-40, 2.003857e-43, 6.403934e-42, 0, 
    4.203895e-45, 1.401298e-45, 0, 1.821688e-44, 8.954297e-43, 9.725011e-43, 
    3.31267e-42, 9.653545e-41, 2.718519e-43, 6.958096e-36, 2.731271e-40, 0, 
    0, 0, 0, 1.778248e-42, 6.165713e-44, 4.145223e-40, 4.135932e-41, 
    1.752395e-39, 2.776281e-40, 2.110412e-40, 1.859103e-41, 3.967076e-42, 
    7.146622e-44, 2.802597e-45, 0, 0, 5.605194e-45, 1.13365e-42, 
    1.272911e-40, 4.616858e-41, 1.325272e-39, 1.387285e-43, 7.229299e-42, 
    1.601684e-42, 7.765576e-41, 1.261169e-44, 2.238434e-41, 1.401298e-45, 
    4.203895e-45, 5.745324e-44, 9.398509e-42, 2.803438e-41, 8.888716e-41, 
    4.368128e-41, 1.290596e-42, 7.160635e-43, 5.324934e-44, 2.662467e-44, 
    2.802597e-45, 0, 2.802597e-45, 1.541428e-44, 1.291997e-42, 6.131381e-41, 
    3.461081e-39, 9.037766e-39, 7.674879e-37, 2.102527e-38, 7.338646e-36, 
    5.195748e-38, 2.272414e-34, 3.390582e-41, 4.467543e-38, 6.445973e-44, 
    3.012792e-43, 4.631291e-42, 1.841181e-39, 7.627968e-41, 3.123243e-39, 
    6.992479e-43, 7.006492e-45, 1.401298e-45, 0, 1.401298e-45, 1.401298e-45, 
    1.541428e-44, 7.006492e-45, 1.493784e-42, 9.10844e-44, 2.096146e-40, 
    3.034485e-39, 3.788231e-36, 2.238026e-34, 1.144245e-32, 6.07666e-32, 
    1.00203e-31, 1.233723e-31,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 F_N2O_DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.809089e-44, 0, 4.13383e-43, 
    7.987401e-44, 1.030235e-41, 2.628836e-42, 9.97866e-40, 1.92146e-41, 
    1.849882e-38, 3.94942e-40, 7.297598e-40, 1.681558e-41, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-44, 1.401298e-45, 2.78438e-42, 
    3.75548e-43, 2.53635e-42, 1.426522e-42, 2.555968e-42, 1.331234e-43, 
    4.764415e-43, 3.363116e-44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.522337e-44, 8.407791e-45, 5.324934e-44, 3.068844e-43, 5.418821e-42, 
    3.398149e-42, 1.178212e-41, 5.044674e-44, 1.961818e-42, 4.203895e-45, 
    2.382207e-44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.508324e-43, 
    9.809089e-45, 5.296908e-43, 7.286752e-44, 2.138381e-42, 1.022948e-43, 
    1.863026e-41, 5.5689e-41, 2.639206e-41, 4.486257e-40, 8.547921e-44, 
    2.53635e-42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.261169e-44, 
    1.667545e-43, 3.503246e-44, 1.387285e-43, 2.942727e-44, 1.401298e-44, 
    3.70111e-41, 4.820467e-43, 3.002072e-40, 2.128642e-40, 1.213384e-41, 
    2.212874e-40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.006492e-45, 
    3.391142e-43, 2.564376e-43, 2.830623e-43, 6.628142e-43, 7.847271e-44, 
    9.360674e-43, 1.408305e-42, 4.820467e-43, 2.032639e-40, 3.770894e-41, 
    2.113102e-40, 7.086086e-41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5.605194e-45, 0, 6.852349e-43, 2.802597e-45, 9.668959e-43, 3.33509e-43, 
    1.930989e-42, 9.042579e-42, 6.074629e-41, 1.833323e-39, 8.431403e-40, 
    1.34621e-38, 0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 2.802597e-45, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.401298e-44, 0, 7.267134e-42, 6.445973e-44, 5.481011e-40, 
    1.98844e-38, 5.055816e-37, 1.874394e-35, 0, 0, 0, 0, 0, 0, 1.401298e-45, 
    1.401298e-45, 1.261169e-44, 6.726233e-44, 2.802597e-45, 1.008935e-43, 0, 
    0, 0, 0, 0, 0, 0, 0, 2.662467e-44, 1.401298e-45, 8.319027e-39, 
    1.249117e-41, 2.604265e-34, 3.383802e-36, 0, 0, 0, 0, 1.401298e-45, 
    5.605194e-45, 3.222986e-44, 2.662467e-43, 3.33509e-43, 1.140657e-42, 
    1.499389e-43, 1.053776e-42, 0, 1.681558e-44, 0, 0, 0, 0, 0, 2.802597e-45, 
    2.802597e-45, 8.407791e-45, 2.578389e-43, 1.401298e-45, 1.858032e-38, 
    7.286752e-43, 0, 0, 0, 0, 4.203895e-45, 0, 1.107026e-42, 1.107026e-43, 
    4.678936e-42, 7.412869e-43, 5.63322e-43, 4.904545e-44, 1.121039e-44, 0, 
    0, 0, 0, 0, 2.802597e-45, 3.405155e-43, 1.233143e-43, 3.538279e-42, 0, 
    1.961818e-44, 4.203895e-45, 2.073922e-43, 0, 6.025583e-44, 0, 0, 0, 
    2.522337e-44, 7.426882e-44, 2.368194e-43, 1.163078e-43, 2.802597e-45, 
    1.401298e-45, 0, 0, 0, 0, 0, 0, 2.802597e-45, 1.639519e-43, 9.241563e-42, 
    2.413316e-41, 2.049435e-39, 5.614442e-41, 1.959651e-38, 1.387426e-40, 
    6.068065e-37, 9.10844e-44, 1.192981e-40, 0, 1.401298e-45, 1.261169e-44, 
    4.917156e-42, 2.031883e-43, 8.340528e-42, 1.401298e-45, 0, 0, 0, 0, 0, 0, 
    0, 4.203895e-45, 0, 5.591181e-43, 8.103709e-42, 1.011577e-38, 
    5.976238e-37, 3.055498e-35, 1.622661e-34, 2.675739e-34, 3.294431e-34 ;

 F_N2O_NIT =
  2.298773e-14, 2.318585e-14, 2.314727e-14, 2.330757e-14, 2.321858e-14, 
    2.332364e-14, 2.302782e-14, 2.319372e-14, 2.308774e-14, 2.300552e-14, 
    2.362028e-14, 2.331471e-14, 2.393994e-14, 2.374342e-14, 2.42387e-14, 
    2.390929e-14, 2.430541e-14, 2.422917e-14, 2.445902e-14, 2.439305e-14, 
    2.468827e-14, 2.448949e-14, 2.484205e-14, 2.464072e-14, 2.467215e-14, 
    2.448293e-14, 2.337607e-14, 2.358214e-14, 2.336388e-14, 2.33932e-14, 
    2.338004e-14, 2.32204e-14, 2.314015e-14, 2.297261e-14, 2.300298e-14, 
    2.312606e-14, 2.340637e-14, 2.331102e-14, 2.355173e-14, 2.354628e-14, 
    2.381574e-14, 2.369404e-14, 2.414937e-14, 2.401949e-14, 2.43958e-14, 
    2.430087e-14, 2.439133e-14, 2.436388e-14, 2.439168e-14, 2.425254e-14, 
    2.431209e-14, 2.418985e-14, 2.371684e-14, 2.385535e-14, 2.344347e-14, 
    2.31976e-14, 2.303507e-14, 2.292009e-14, 2.293632e-14, 2.296729e-14, 
    2.312677e-14, 2.327726e-14, 2.339228e-14, 2.346938e-14, 2.354549e-14, 
    2.377661e-14, 2.389944e-14, 2.417566e-14, 2.41257e-14, 2.421038e-14, 
    2.429143e-14, 2.442782e-14, 2.440535e-14, 2.446553e-14, 2.420813e-14, 
    2.437903e-14, 2.409724e-14, 2.417414e-14, 2.356619e-14, 2.333674e-14, 
    2.323954e-14, 2.315466e-14, 2.294881e-14, 2.309086e-14, 2.30348e-14, 
    2.316827e-14, 2.325329e-14, 2.321122e-14, 2.347149e-14, 2.337012e-14, 
    2.390673e-14, 2.367481e-14, 2.428197e-14, 2.413594e-14, 2.431704e-14, 
    2.422454e-14, 2.438313e-14, 2.424037e-14, 2.448795e-14, 2.454203e-14, 
    2.450506e-14, 2.464723e-14, 2.423245e-14, 2.43913e-14, 2.321005e-14, 
    2.321691e-14, 2.324887e-14, 2.310852e-14, 2.309995e-14, 2.297176e-14, 
    2.30858e-14, 2.313446e-14, 2.325821e-14, 2.333157e-14, 2.340142e-14, 
    2.355539e-14, 2.372797e-14, 2.397041e-14, 2.414539e-14, 2.426306e-14, 
    2.419087e-14, 2.425459e-14, 2.418336e-14, 2.415001e-14, 2.452175e-14, 
    2.431264e-14, 2.462674e-14, 2.460931e-14, 2.446694e-14, 2.461126e-14, 
    2.322172e-14, 2.318226e-14, 2.304554e-14, 2.31525e-14, 2.295782e-14, 
    2.306668e-14, 2.312939e-14, 2.337222e-14, 2.342576e-14, 2.347545e-14, 
    2.357376e-14, 2.370024e-14, 2.392298e-14, 2.411768e-14, 2.429614e-14, 
    2.428304e-14, 2.428765e-14, 2.43276e-14, 2.422869e-14, 2.434385e-14, 
    2.43632e-14, 2.431261e-14, 2.460696e-14, 2.452268e-14, 2.460893e-14, 
    2.455402e-14, 2.319508e-14, 2.326151e-14, 2.322559e-14, 2.329314e-14, 
    2.324553e-14, 2.345757e-14, 2.352134e-14, 2.382094e-14, 2.369775e-14, 
    2.389398e-14, 2.371764e-14, 2.374883e-14, 2.390037e-14, 2.372714e-14, 
    2.41069e-14, 2.384907e-14, 2.432914e-14, 2.407041e-14, 2.43454e-14, 
    2.429535e-14, 2.437824e-14, 2.445261e-14, 2.454634e-14, 2.471978e-14, 
    2.467956e-14, 2.482498e-14, 2.336072e-14, 2.344721e-14, 2.34396e-14, 
    2.353028e-14, 2.359747e-14, 2.374345e-14, 2.397855e-14, 2.389e-14, 
    2.40527e-14, 2.408543e-14, 2.383829e-14, 2.398987e-14, 2.350517e-14, 
    2.358312e-14, 2.35367e-14, 2.336749e-14, 2.391036e-14, 2.363093e-14, 
    2.414826e-14, 2.399588e-14, 2.444199e-14, 2.421958e-14, 2.465743e-14, 
    2.484585e-14, 2.50239e-14, 2.523278e-14, 2.34945e-14, 2.343564e-14, 
    2.354108e-14, 2.368736e-14, 2.382353e-14, 2.400519e-14, 2.402382e-14, 
    2.405793e-14, 2.414645e-14, 2.4221e-14, 2.406872e-14, 2.42397e-14, 
    2.36012e-14, 2.393469e-14, 2.341336e-14, 2.35697e-14, 2.367869e-14, 
    2.363085e-14, 2.387985e-14, 2.393873e-14, 2.41788e-14, 2.405454e-14, 
    2.479926e-14, 2.446831e-14, 2.539245e-14, 2.513238e-14, 2.341509e-14, 
    2.349429e-14, 2.377102e-14, 2.363914e-14, 2.401734e-14, 2.411091e-14, 
    2.418712e-14, 2.428472e-14, 2.429527e-14, 2.435321e-14, 2.42583e-14, 
    2.434945e-14, 2.400555e-14, 2.415891e-14, 2.373928e-14, 2.384105e-14, 
    2.37942e-14, 2.374286e-14, 2.390148e-14, 2.407108e-14, 2.407471e-14, 
    2.412923e-14, 2.428318e-14, 2.401882e-14, 2.484212e-14, 2.433193e-14, 
    2.358081e-14, 2.373404e-14, 2.375598e-14, 2.369653e-14, 2.410151e-14, 
    2.395435e-14, 2.43518e-14, 2.424404e-14, 2.442072e-14, 2.433284e-14, 
    2.431992e-14, 2.420732e-14, 2.413735e-14, 2.396106e-14, 2.381813e-14, 
    2.370511e-14, 2.373136e-14, 2.385559e-14, 2.408147e-14, 2.429618e-14, 
    2.424906e-14, 2.440723e-14, 2.398975e-14, 2.416434e-14, 2.409677e-14, 
    2.427315e-14, 2.388764e-14, 2.421574e-14, 2.380414e-14, 2.384008e-14, 
    2.395143e-14, 2.417624e-14, 2.422614e-14, 2.427946e-14, 2.424655e-14, 
    2.408724e-14, 2.406119e-14, 2.39487e-14, 2.391768e-14, 2.383222e-14, 
    2.376158e-14, 2.382611e-14, 2.389397e-14, 2.408729e-14, 2.426219e-14, 
    2.445363e-14, 2.450061e-14, 2.47255e-14, 2.454233e-14, 2.484496e-14, 
    2.458752e-14, 2.503406e-14, 2.423483e-14, 2.458004e-14, 2.395651e-14, 
    2.402327e-14, 2.414429e-14, 2.442306e-14, 2.427235e-14, 2.444865e-14, 
    2.406017e-14, 2.385989e-14, 2.380822e-14, 2.371197e-14, 2.381042e-14, 
    2.38024e-14, 2.389679e-14, 2.386644e-14, 2.409371e-14, 2.397149e-14, 
    2.431955e-14, 2.444723e-14, 2.480968e-14, 2.503326e-14, 2.526194e-14, 
    2.536324e-14, 2.539412e-14, 2.540703e-14 ;

 F_NIT =
  3.831289e-11, 3.864309e-11, 3.857878e-11, 3.884595e-11, 3.869762e-11, 
    3.887273e-11, 3.83797e-11, 3.865619e-11, 3.847956e-11, 3.834253e-11, 
    3.936713e-11, 3.885786e-11, 3.98999e-11, 3.957237e-11, 4.039783e-11, 
    3.984882e-11, 4.050901e-11, 4.038195e-11, 4.076504e-11, 4.065509e-11, 
    4.114711e-11, 4.081582e-11, 4.140342e-11, 4.106787e-11, 4.112025e-11, 
    4.080489e-11, 3.896012e-11, 3.930356e-11, 3.89398e-11, 3.898867e-11, 
    3.896674e-11, 3.870066e-11, 3.856692e-11, 3.828768e-11, 3.833829e-11, 
    3.854343e-11, 3.901062e-11, 3.88517e-11, 3.925288e-11, 3.92438e-11, 
    3.96929e-11, 3.949007e-11, 4.024895e-11, 4.003249e-11, 4.065967e-11, 
    4.050145e-11, 4.065222e-11, 4.060646e-11, 4.06528e-11, 4.04209e-11, 
    4.052016e-11, 4.031641e-11, 3.952807e-11, 3.975893e-11, 3.907245e-11, 
    3.866267e-11, 3.839178e-11, 3.820015e-11, 3.822721e-11, 3.827882e-11, 
    3.854463e-11, 3.879543e-11, 3.898714e-11, 3.911564e-11, 3.924248e-11, 
    3.962769e-11, 3.983241e-11, 4.029277e-11, 4.02095e-11, 4.035063e-11, 
    4.048572e-11, 4.071304e-11, 4.067558e-11, 4.077588e-11, 4.034689e-11, 
    4.063172e-11, 4.016206e-11, 4.029023e-11, 3.927698e-11, 3.889456e-11, 
    3.873256e-11, 3.859109e-11, 3.824802e-11, 3.848476e-11, 3.839133e-11, 
    3.861378e-11, 3.875547e-11, 3.868536e-11, 3.911915e-11, 3.895019e-11, 
    3.984455e-11, 3.945801e-11, 4.046996e-11, 4.022658e-11, 4.052839e-11, 
    4.037424e-11, 4.063855e-11, 4.040062e-11, 4.081325e-11, 4.090338e-11, 
    4.084176e-11, 4.107871e-11, 4.038742e-11, 4.065216e-11, 3.868342e-11, 
    3.869485e-11, 3.874812e-11, 3.85142e-11, 3.849992e-11, 3.828626e-11, 
    3.847634e-11, 3.855742e-11, 3.876369e-11, 3.888595e-11, 3.900237e-11, 
    3.925899e-11, 3.954662e-11, 3.995068e-11, 4.024232e-11, 4.043842e-11, 
    4.031812e-11, 4.042431e-11, 4.030559e-11, 4.025001e-11, 4.086958e-11, 
    4.052106e-11, 4.104457e-11, 4.101551e-11, 4.077823e-11, 4.101878e-11, 
    3.870287e-11, 3.86371e-11, 3.840923e-11, 3.858749e-11, 3.826303e-11, 
    3.844446e-11, 3.854898e-11, 3.89537e-11, 3.904293e-11, 3.912575e-11, 
    3.92896e-11, 3.95004e-11, 3.987164e-11, 4.019613e-11, 4.049357e-11, 
    4.047173e-11, 4.047941e-11, 4.054599e-11, 4.038115e-11, 4.057308e-11, 
    4.060533e-11, 4.052102e-11, 4.101161e-11, 4.087113e-11, 4.101488e-11, 
    4.092338e-11, 3.865847e-11, 3.876918e-11, 3.870932e-11, 3.88219e-11, 
    3.874255e-11, 3.909595e-11, 3.920223e-11, 3.970157e-11, 3.949625e-11, 
    3.98233e-11, 3.95294e-11, 3.958139e-11, 3.983395e-11, 3.954524e-11, 
    4.017817e-11, 3.974846e-11, 4.054857e-11, 4.011736e-11, 4.057567e-11, 
    4.049224e-11, 4.063041e-11, 4.075435e-11, 4.091057e-11, 4.119964e-11, 
    4.11326e-11, 4.137497e-11, 3.893453e-11, 3.907869e-11, 3.9066e-11, 
    3.921714e-11, 3.932911e-11, 3.957241e-11, 3.996426e-11, 3.981666e-11, 
    4.008784e-11, 4.014239e-11, 3.973049e-11, 3.998311e-11, 3.917529e-11, 
    3.93052e-11, 3.922783e-11, 3.894582e-11, 3.985059e-11, 3.938488e-11, 
    4.024709e-11, 3.999313e-11, 4.073665e-11, 4.036597e-11, 4.109572e-11, 
    4.140975e-11, 4.17065e-11, 4.205463e-11, 3.91575e-11, 3.90594e-11, 
    3.923513e-11, 3.947893e-11, 3.970588e-11, 4.000865e-11, 4.003969e-11, 
    4.009656e-11, 4.024408e-11, 4.036834e-11, 4.011453e-11, 4.039951e-11, 
    3.933533e-11, 3.989115e-11, 3.902227e-11, 3.928284e-11, 3.946448e-11, 
    3.938476e-11, 3.979976e-11, 3.989789e-11, 4.029799e-11, 4.009091e-11, 
    4.13321e-11, 4.078051e-11, 4.232075e-11, 4.188729e-11, 3.902515e-11, 
    3.915714e-11, 3.961837e-11, 3.939856e-11, 4.002889e-11, 4.018485e-11, 
    4.031187e-11, 4.047454e-11, 4.049212e-11, 4.058868e-11, 4.04305e-11, 
    4.058242e-11, 4.000924e-11, 4.026485e-11, 3.956547e-11, 3.973508e-11, 
    3.9657e-11, 3.957144e-11, 3.98358e-11, 4.011846e-11, 4.012453e-11, 
    4.021538e-11, 4.047196e-11, 4.003137e-11, 4.140353e-11, 4.055322e-11, 
    3.930135e-11, 3.955673e-11, 3.959329e-11, 3.949421e-11, 4.016919e-11, 
    3.992392e-11, 4.058633e-11, 4.040673e-11, 4.07012e-11, 4.055473e-11, 
    4.053319e-11, 4.034554e-11, 4.022892e-11, 3.993511e-11, 3.969688e-11, 
    3.950852e-11, 3.955227e-11, 3.975932e-11, 4.013578e-11, 4.049364e-11, 
    4.04151e-11, 4.067872e-11, 3.998292e-11, 4.027391e-11, 4.016129e-11, 
    4.045525e-11, 3.981272e-11, 4.035956e-11, 3.967356e-11, 3.973346e-11, 
    3.991905e-11, 4.029374e-11, 4.03769e-11, 4.046577e-11, 4.041092e-11, 
    4.01454e-11, 4.010198e-11, 3.99145e-11, 3.986281e-11, 3.972037e-11, 
    3.960263e-11, 3.971019e-11, 3.982329e-11, 4.014548e-11, 4.043698e-11, 
    4.075606e-11, 4.083435e-11, 4.120916e-11, 4.090388e-11, 4.140826e-11, 
    4.09792e-11, 4.172343e-11, 4.039138e-11, 4.096674e-11, 3.992751e-11, 
    4.003879e-11, 4.024048e-11, 4.070509e-11, 4.045392e-11, 4.074775e-11, 
    4.010028e-11, 3.976648e-11, 3.968037e-11, 3.951995e-11, 3.968403e-11, 
    3.967067e-11, 3.982799e-11, 3.977739e-11, 4.015618e-11, 3.995248e-11, 
    4.053259e-11, 4.074538e-11, 4.134947e-11, 4.172209e-11, 4.210324e-11, 
    4.227207e-11, 4.232353e-11, 4.234505e-11 ;

 F_NIT_vr =
  2.424388e-10, 2.435265e-10, 2.433145e-10, 2.441924e-10, 2.437051e-10, 
    2.442796e-10, 2.426581e-10, 2.435677e-10, 2.429867e-10, 2.425347e-10, 
    2.45896e-10, 2.442295e-10, 2.476323e-10, 2.465661e-10, 2.492463e-10, 
    2.474654e-10, 2.496057e-10, 2.491947e-10, 2.504321e-10, 2.50077e-10, 
    2.516604e-10, 2.505951e-10, 2.524827e-10, 2.514056e-10, 2.515735e-10, 
    2.505586e-10, 2.445669e-10, 2.456901e-10, 2.444998e-10, 2.446599e-10, 
    2.445878e-10, 2.437139e-10, 2.432736e-10, 2.423536e-10, 2.425202e-10, 
    2.431959e-10, 2.4473e-10, 2.442087e-10, 2.455227e-10, 2.454931e-10, 
    2.469579e-10, 2.462969e-10, 2.487638e-10, 2.480615e-10, 2.500915e-10, 
    2.4958e-10, 2.500669e-10, 2.499188e-10, 2.50068e-10, 2.493187e-10, 
    2.496391e-10, 2.489801e-10, 2.464237e-10, 2.471754e-10, 2.44934e-10, 
    2.435883e-10, 2.426968e-10, 2.420647e-10, 2.421535e-10, 2.423237e-10, 
    2.431993e-10, 2.440238e-10, 2.446527e-10, 2.450733e-10, 2.45488e-10, 
    2.467446e-10, 2.47411e-10, 2.489049e-10, 2.486353e-10, 2.490917e-10, 
    2.495289e-10, 2.502625e-10, 2.501416e-10, 2.504646e-10, 2.490786e-10, 
    2.499992e-10, 2.484794e-10, 2.488947e-10, 2.45602e-10, 2.443505e-10, 
    2.438178e-10, 2.433528e-10, 2.422219e-10, 2.430024e-10, 2.426943e-10, 
    2.434266e-10, 2.438922e-10, 2.436615e-10, 2.450845e-10, 2.445305e-10, 
    2.474502e-10, 2.461912e-10, 2.494782e-10, 2.486901e-10, 2.496664e-10, 
    2.49168e-10, 2.500216e-10, 2.492529e-10, 2.505846e-10, 2.508749e-10, 
    2.506759e-10, 2.514387e-10, 2.492086e-10, 2.50064e-10, 2.436566e-10, 
    2.436942e-10, 2.43869e-10, 2.430989e-10, 2.430519e-10, 2.423474e-10, 
    2.429736e-10, 2.432405e-10, 2.439187e-10, 2.443195e-10, 2.44701e-10, 
    2.455411e-10, 2.464797e-10, 2.477945e-10, 2.487408e-10, 2.493753e-10, 
    2.489859e-10, 2.493291e-10, 2.489448e-10, 2.487644e-10, 2.507652e-10, 
    2.496409e-10, 2.513282e-10, 2.512348e-10, 2.504701e-10, 2.512446e-10, 
    2.4372e-10, 2.435035e-10, 2.42753e-10, 2.433398e-10, 2.422702e-10, 
    2.428684e-10, 2.432121e-10, 2.445413e-10, 2.448338e-10, 2.45105e-10, 
    2.456407e-10, 2.463287e-10, 2.475374e-10, 2.485904e-10, 2.495533e-10, 
    2.494823e-10, 2.49507e-10, 2.497217e-10, 2.491886e-10, 2.498087e-10, 
    2.499124e-10, 2.496403e-10, 2.512215e-10, 2.507694e-10, 2.512318e-10, 
    2.509369e-10, 2.435735e-10, 2.439368e-10, 2.437399e-10, 2.441096e-10, 
    2.438484e-10, 2.450074e-10, 2.453548e-10, 2.469842e-10, 2.46315e-10, 
    2.473803e-10, 2.464227e-10, 2.465922e-10, 2.474135e-10, 2.464738e-10, 
    2.485311e-10, 2.471347e-10, 2.497298e-10, 2.483327e-10, 2.498168e-10, 
    2.495469e-10, 2.499929e-10, 2.503927e-10, 2.508956e-10, 2.51825e-10, 
    2.516092e-10, 2.523872e-10, 2.444793e-10, 2.449511e-10, 2.449097e-10, 
    2.45404e-10, 2.457697e-10, 2.465639e-10, 2.478386e-10, 2.473586e-10, 
    2.482392e-10, 2.484162e-10, 2.470774e-10, 2.478985e-10, 2.452648e-10, 
    2.45689e-10, 2.454363e-10, 2.445123e-10, 2.474664e-10, 2.459483e-10, 
    2.487531e-10, 2.47929e-10, 2.503349e-10, 2.491372e-10, 2.514905e-10, 
    2.524979e-10, 2.534481e-10, 2.54558e-10, 2.45209e-10, 2.448876e-10, 
    2.454624e-10, 2.462584e-10, 2.469979e-10, 2.479824e-10, 2.48083e-10, 
    2.482671e-10, 2.487452e-10, 2.491475e-10, 2.483245e-10, 2.492477e-10, 
    2.457866e-10, 2.475984e-10, 2.447624e-10, 2.456149e-10, 2.462079e-10, 
    2.459478e-10, 2.473004e-10, 2.47619e-10, 2.489165e-10, 2.482456e-10, 
    2.522481e-10, 2.504748e-10, 2.554048e-10, 2.540241e-10, 2.44775e-10, 
    2.452069e-10, 2.467125e-10, 2.459958e-10, 2.480476e-10, 2.485535e-10, 
    2.489645e-10, 2.494907e-10, 2.495471e-10, 2.498591e-10, 2.493474e-10, 
    2.498385e-10, 2.479816e-10, 2.488107e-10, 2.465377e-10, 2.470897e-10, 
    2.468355e-10, 2.465562e-10, 2.474167e-10, 2.483343e-10, 2.483541e-10, 
    2.48648e-10, 2.494771e-10, 2.480509e-10, 2.524753e-10, 2.49739e-10, 
    2.456783e-10, 2.46511e-10, 2.466303e-10, 2.463074e-10, 2.485019e-10, 
    2.477059e-10, 2.498515e-10, 2.492707e-10, 2.502216e-10, 2.497488e-10, 
    2.496786e-10, 2.490719e-10, 2.486936e-10, 2.477402e-10, 2.469647e-10, 
    2.463511e-10, 2.464932e-10, 2.471675e-10, 2.483898e-10, 2.495487e-10, 
    2.492943e-10, 2.501459e-10, 2.478931e-10, 2.488367e-10, 2.484711e-10, 
    2.494232e-10, 2.473446e-10, 2.491177e-10, 2.468916e-10, 2.470862e-10, 
    2.476893e-10, 2.489045e-10, 2.491737e-10, 2.49461e-10, 2.492832e-10, 
    2.48423e-10, 2.48282e-10, 2.47673e-10, 2.475044e-10, 2.470413e-10, 
    2.466572e-10, 2.470076e-10, 2.473749e-10, 2.484214e-10, 2.49365e-10, 
    2.50395e-10, 2.506475e-10, 2.518517e-10, 2.508702e-10, 2.524891e-10, 
    2.51111e-10, 2.534978e-10, 2.492205e-10, 2.51077e-10, 2.47717e-10, 
    2.48078e-10, 2.487315e-10, 2.502331e-10, 2.49422e-10, 2.503705e-10, 
    2.482763e-10, 2.47191e-10, 2.469108e-10, 2.463879e-10, 2.469222e-10, 
    2.468788e-10, 2.473905e-10, 2.472255e-10, 2.484554e-10, 2.477944e-10, 
    2.496732e-10, 2.5036e-10, 2.523023e-10, 2.534946e-10, 2.547109e-10, 
    2.552477e-10, 2.554112e-10, 2.554793e-10,
  1.243035e-10, 1.252448e-10, 1.250617e-10, 1.258223e-10, 1.254002e-10, 
    1.258985e-10, 1.244942e-10, 1.252821e-10, 1.24779e-10, 1.243883e-10, 
    1.27303e-10, 1.258563e-10, 1.288132e-10, 1.278856e-10, 1.302207e-10, 
    1.286685e-10, 1.305346e-10, 1.301761e-10, 1.312567e-10, 1.309468e-10, 
    1.323321e-10, 1.313999e-10, 1.330527e-10, 1.321094e-10, 1.322567e-10, 
    1.313691e-10, 1.261471e-10, 1.271225e-10, 1.260893e-10, 1.262283e-10, 
    1.26166e-10, 1.254088e-10, 1.250278e-10, 1.242318e-10, 1.243762e-10, 
    1.24961e-10, 1.262907e-10, 1.258389e-10, 1.269792e-10, 1.269534e-10, 
    1.282272e-10, 1.276523e-10, 1.298005e-10, 1.291886e-10, 1.309598e-10, 
    1.305135e-10, 1.309387e-10, 1.308098e-10, 1.309404e-10, 1.302861e-10, 
    1.305663e-10, 1.299912e-10, 1.277599e-10, 1.284141e-10, 1.264665e-10, 
    1.253004e-10, 1.245287e-10, 1.23982e-10, 1.240593e-10, 1.242065e-10, 
    1.249644e-10, 1.256788e-10, 1.262241e-10, 1.265894e-10, 1.269497e-10, 
    1.280421e-10, 1.286222e-10, 1.299242e-10, 1.296891e-10, 1.300876e-10, 
    1.304691e-10, 1.311102e-10, 1.310047e-10, 1.312874e-10, 1.300773e-10, 
    1.30881e-10, 1.295552e-10, 1.299173e-10, 1.27047e-10, 1.259608e-10, 
    1.254995e-10, 1.250968e-10, 1.241186e-10, 1.247938e-10, 1.245275e-10, 
    1.251616e-10, 1.255651e-10, 1.253655e-10, 1.265994e-10, 1.261191e-10, 
    1.286566e-10, 1.275613e-10, 1.304246e-10, 1.297373e-10, 1.305896e-10, 
    1.301545e-10, 1.309002e-10, 1.30229e-10, 1.313927e-10, 1.316465e-10, 
    1.31473e-10, 1.321401e-10, 1.301918e-10, 1.309387e-10, 1.253599e-10, 
    1.253924e-10, 1.255441e-10, 1.248777e-10, 1.248371e-10, 1.242279e-10, 
    1.247699e-10, 1.25001e-10, 1.255885e-10, 1.259364e-10, 1.262675e-10, 
    1.269966e-10, 1.278126e-10, 1.289571e-10, 1.297818e-10, 1.303357e-10, 
    1.29996e-10, 1.302959e-10, 1.299607e-10, 1.298037e-10, 1.315513e-10, 
    1.305689e-10, 1.320441e-10, 1.319623e-10, 1.31294e-10, 1.319715e-10, 
    1.254152e-10, 1.25228e-10, 1.245786e-10, 1.250867e-10, 1.241616e-10, 
    1.24679e-10, 1.249769e-10, 1.26129e-10, 1.263828e-10, 1.266181e-10, 
    1.270836e-10, 1.276817e-10, 1.287335e-10, 1.296513e-10, 1.304914e-10, 
    1.304298e-10, 1.304514e-10, 1.306393e-10, 1.301741e-10, 1.307157e-10, 
    1.308066e-10, 1.305688e-10, 1.319514e-10, 1.315559e-10, 1.319606e-10, 
    1.31703e-10, 1.252889e-10, 1.256041e-10, 1.254337e-10, 1.257541e-10, 
    1.255283e-10, 1.265333e-10, 1.268353e-10, 1.282517e-10, 1.276699e-10, 
    1.285966e-10, 1.27764e-10, 1.279113e-10, 1.286265e-10, 1.278089e-10, 
    1.296005e-10, 1.283846e-10, 1.306466e-10, 1.294285e-10, 1.30723e-10, 
    1.304877e-10, 1.308775e-10, 1.312268e-10, 1.31667e-10, 1.324802e-10, 
    1.322918e-10, 1.329731e-10, 1.260746e-10, 1.264844e-10, 1.264484e-10, 
    1.268778e-10, 1.271957e-10, 1.278859e-10, 1.289956e-10, 1.285779e-10, 
    1.293453e-10, 1.294995e-10, 1.283339e-10, 1.29049e-10, 1.26759e-10, 
    1.271278e-10, 1.269082e-10, 1.261068e-10, 1.28674e-10, 1.27354e-10, 
    1.297955e-10, 1.290775e-10, 1.31177e-10, 1.301312e-10, 1.321881e-10, 
    1.330706e-10, 1.339037e-10, 1.34879e-10, 1.267083e-10, 1.264297e-10, 
    1.269289e-10, 1.276207e-10, 1.282641e-10, 1.291212e-10, 1.292091e-10, 
    1.293699e-10, 1.297869e-10, 1.301379e-10, 1.294206e-10, 1.302259e-10, 
    1.272131e-10, 1.287888e-10, 1.263242e-10, 1.270643e-10, 1.275799e-10, 
    1.273538e-10, 1.285303e-10, 1.288081e-10, 1.299393e-10, 1.293541e-10, 
    1.328524e-10, 1.313005e-10, 1.356237e-10, 1.344104e-10, 1.263323e-10, 
    1.267075e-10, 1.280161e-10, 1.273928e-10, 1.291786e-10, 1.296195e-10, 
    1.299784e-10, 1.304376e-10, 1.304873e-10, 1.307597e-10, 1.303134e-10, 
    1.307421e-10, 1.29123e-10, 1.298457e-10, 1.278664e-10, 1.28347e-10, 
    1.281259e-10, 1.278834e-10, 1.286324e-10, 1.294319e-10, 1.294492e-10, 
    1.297059e-10, 1.3043e-10, 1.291858e-10, 1.330528e-10, 1.306594e-10, 
    1.27117e-10, 1.278413e-10, 1.279451e-10, 1.276642e-10, 1.295753e-10, 
    1.288816e-10, 1.307531e-10, 1.302464e-10, 1.310771e-10, 1.30664e-10, 
    1.306033e-10, 1.300736e-10, 1.297442e-10, 1.289133e-10, 1.282388e-10, 
    1.27705e-10, 1.278291e-10, 1.284157e-10, 1.294809e-10, 1.304917e-10, 
    1.3027e-10, 1.310139e-10, 1.290488e-10, 1.298713e-10, 1.295531e-10, 
    1.303835e-10, 1.285668e-10, 1.301126e-10, 1.281727e-10, 1.283424e-10, 
    1.288678e-10, 1.29927e-10, 1.301621e-10, 1.304129e-10, 1.302582e-10, 
    1.29508e-10, 1.293854e-10, 1.288551e-10, 1.287087e-10, 1.283055e-10, 
    1.279719e-10, 1.282766e-10, 1.285969e-10, 1.295084e-10, 1.303318e-10, 
    1.312318e-10, 1.314524e-10, 1.325069e-10, 1.31648e-10, 1.330661e-10, 
    1.318596e-10, 1.339509e-10, 1.302027e-10, 1.318247e-10, 1.288918e-10, 
    1.292067e-10, 1.297766e-10, 1.310878e-10, 1.303796e-10, 1.312081e-10, 
    1.293806e-10, 1.284359e-10, 1.281921e-10, 1.277374e-10, 1.282025e-10, 
    1.281647e-10, 1.286103e-10, 1.28467e-10, 1.295387e-10, 1.289627e-10, 
    1.306017e-10, 1.312016e-10, 1.329016e-10, 1.339474e-10, 1.350155e-10, 
    1.354878e-10, 1.356317e-10, 1.356919e-10,
  1.174377e-10, 1.18479e-10, 1.182763e-10, 1.191184e-10, 1.18651e-10, 
    1.192028e-10, 1.176485e-10, 1.185204e-10, 1.179635e-10, 1.175313e-10, 
    1.207598e-10, 1.191561e-10, 1.224358e-10, 1.214058e-10, 1.240003e-10, 
    1.222752e-10, 1.243494e-10, 1.239505e-10, 1.25153e-10, 1.24808e-10, 
    1.263511e-10, 1.253123e-10, 1.271543e-10, 1.261027e-10, 1.262669e-10, 
    1.252781e-10, 1.194782e-10, 1.205596e-10, 1.194142e-10, 1.195681e-10, 
    1.194991e-10, 1.186606e-10, 1.182389e-10, 1.173583e-10, 1.17518e-10, 
    1.18165e-10, 1.196374e-10, 1.191368e-10, 1.204004e-10, 1.203718e-10, 
    1.21785e-10, 1.21147e-10, 1.235328e-10, 1.228527e-10, 1.248224e-10, 
    1.243258e-10, 1.24799e-10, 1.246555e-10, 1.248009e-10, 1.240729e-10, 
    1.243846e-10, 1.237448e-10, 1.212663e-10, 1.219925e-10, 1.198321e-10, 
    1.185408e-10, 1.176867e-10, 1.170821e-10, 1.171675e-10, 1.173303e-10, 
    1.181687e-10, 1.189594e-10, 1.195635e-10, 1.199683e-10, 1.203677e-10, 
    1.215798e-10, 1.222237e-10, 1.236705e-10, 1.234089e-10, 1.238522e-10, 
    1.242764e-10, 1.249899e-10, 1.248724e-10, 1.251871e-10, 1.238406e-10, 
    1.247348e-10, 1.232601e-10, 1.236626e-10, 1.204759e-10, 1.192717e-10, 
    1.187611e-10, 1.183152e-10, 1.172332e-10, 1.179799e-10, 1.176853e-10, 
    1.183869e-10, 1.188335e-10, 1.186126e-10, 1.199793e-10, 1.194472e-10, 
    1.222619e-10, 1.210461e-10, 1.242269e-10, 1.234626e-10, 1.244104e-10, 
    1.239264e-10, 1.247562e-10, 1.240093e-10, 1.253044e-10, 1.255871e-10, 
    1.253938e-10, 1.261369e-10, 1.239679e-10, 1.24799e-10, 1.186063e-10, 
    1.186424e-10, 1.188103e-10, 1.180728e-10, 1.180278e-10, 1.173539e-10, 
    1.179535e-10, 1.182092e-10, 1.188595e-10, 1.192448e-10, 1.196116e-10, 
    1.204197e-10, 1.213249e-10, 1.225956e-10, 1.235121e-10, 1.24128e-10, 
    1.237502e-10, 1.240837e-10, 1.237109e-10, 1.235363e-10, 1.254811e-10, 
    1.243875e-10, 1.260299e-10, 1.259388e-10, 1.251946e-10, 1.259491e-10, 
    1.186677e-10, 1.184604e-10, 1.177418e-10, 1.18304e-10, 1.172806e-10, 
    1.178529e-10, 1.181825e-10, 1.194582e-10, 1.197393e-10, 1.200001e-10, 
    1.205161e-10, 1.211796e-10, 1.223472e-10, 1.23367e-10, 1.243012e-10, 
    1.242326e-10, 1.242567e-10, 1.244657e-10, 1.239482e-10, 1.245508e-10, 
    1.24652e-10, 1.243874e-10, 1.259266e-10, 1.254861e-10, 1.259369e-10, 
    1.256499e-10, 1.185278e-10, 1.188767e-10, 1.186881e-10, 1.190429e-10, 
    1.187929e-10, 1.199062e-10, 1.202409e-10, 1.218123e-10, 1.211665e-10, 
    1.221952e-10, 1.212708e-10, 1.214344e-10, 1.222286e-10, 1.213207e-10, 
    1.233106e-10, 1.219599e-10, 1.244739e-10, 1.231195e-10, 1.245589e-10, 
    1.242971e-10, 1.247308e-10, 1.251197e-10, 1.256098e-10, 1.26516e-10, 
    1.26306e-10, 1.270655e-10, 1.193978e-10, 1.198519e-10, 1.19812e-10, 
    1.202879e-10, 1.206405e-10, 1.214061e-10, 1.226383e-10, 1.221744e-10, 
    1.230268e-10, 1.231982e-10, 1.219034e-10, 1.226976e-10, 1.201563e-10, 
    1.205653e-10, 1.203217e-10, 1.194336e-10, 1.222811e-10, 1.208161e-10, 
    1.235272e-10, 1.227293e-10, 1.250642e-10, 1.239006e-10, 1.261903e-10, 
    1.271743e-10, 1.281037e-10, 1.291928e-10, 1.201001e-10, 1.197912e-10, 
    1.203446e-10, 1.21112e-10, 1.21826e-10, 1.227779e-10, 1.228755e-10, 
    1.230542e-10, 1.235177e-10, 1.23908e-10, 1.231107e-10, 1.240059e-10, 
    1.2066e-10, 1.224087e-10, 1.196745e-10, 1.204949e-10, 1.210667e-10, 
    1.208158e-10, 1.221214e-10, 1.2243e-10, 1.236872e-10, 1.230367e-10, 
    1.269311e-10, 1.252018e-10, 1.30025e-10, 1.286694e-10, 1.196833e-10, 
    1.200991e-10, 1.215507e-10, 1.208591e-10, 1.228416e-10, 1.233316e-10, 
    1.237307e-10, 1.242414e-10, 1.242967e-10, 1.245998e-10, 1.241032e-10, 
    1.245802e-10, 1.227799e-10, 1.23583e-10, 1.213845e-10, 1.21918e-10, 
    1.216725e-10, 1.214033e-10, 1.222348e-10, 1.231232e-10, 1.231423e-10, 
    1.234277e-10, 1.242333e-10, 1.228496e-10, 1.271548e-10, 1.244885e-10, 
    1.205531e-10, 1.213568e-10, 1.214719e-10, 1.211602e-10, 1.232824e-10, 
    1.225117e-10, 1.245924e-10, 1.240286e-10, 1.249529e-10, 1.244933e-10, 
    1.244257e-10, 1.238365e-10, 1.234702e-10, 1.225469e-10, 1.217979e-10, 
    1.212054e-10, 1.21343e-10, 1.219943e-10, 1.231776e-10, 1.243016e-10, 
    1.24055e-10, 1.248826e-10, 1.226974e-10, 1.236116e-10, 1.232579e-10, 
    1.241812e-10, 1.22162e-10, 1.238802e-10, 1.217244e-10, 1.219128e-10, 
    1.224964e-10, 1.236737e-10, 1.23935e-10, 1.24214e-10, 1.240418e-10, 
    1.232078e-10, 1.230714e-10, 1.224822e-10, 1.223197e-10, 1.218718e-10, 
    1.215015e-10, 1.218398e-10, 1.221955e-10, 1.232082e-10, 1.241237e-10, 
    1.251252e-10, 1.253709e-10, 1.265459e-10, 1.255889e-10, 1.271696e-10, 
    1.258249e-10, 1.281567e-10, 1.239803e-10, 1.257857e-10, 1.22523e-10, 
    1.228728e-10, 1.235064e-10, 1.249651e-10, 1.241768e-10, 1.25099e-10, 
    1.230661e-10, 1.220167e-10, 1.21746e-10, 1.212413e-10, 1.217576e-10, 
    1.217155e-10, 1.222103e-10, 1.220512e-10, 1.232418e-10, 1.226017e-10, 
    1.244239e-10, 1.250917e-10, 1.269857e-10, 1.281526e-10, 1.293451e-10, 
    1.29873e-10, 1.300338e-10, 1.301011e-10,
  1.205484e-10, 1.216951e-10, 1.214718e-10, 1.223997e-10, 1.218846e-10, 
    1.224928e-10, 1.207805e-10, 1.217407e-10, 1.211273e-10, 1.206514e-10, 
    1.242102e-10, 1.224412e-10, 1.260609e-10, 1.249231e-10, 1.277908e-10, 
    1.258835e-10, 1.281771e-10, 1.277356e-10, 1.290666e-10, 1.286846e-10, 
    1.303942e-10, 1.292431e-10, 1.312848e-10, 1.301189e-10, 1.303009e-10, 
    1.292052e-10, 1.227962e-10, 1.239892e-10, 1.227257e-10, 1.228955e-10, 
    1.228193e-10, 1.218952e-10, 1.214308e-10, 1.20461e-10, 1.206368e-10, 
    1.213492e-10, 1.229718e-10, 1.224199e-10, 1.238133e-10, 1.237818e-10, 
    1.253419e-10, 1.246373e-10, 1.272736e-10, 1.265216e-10, 1.287006e-10, 
    1.281509e-10, 1.286747e-10, 1.285158e-10, 1.286768e-10, 1.278711e-10, 
    1.28216e-10, 1.275081e-10, 1.247691e-10, 1.255711e-10, 1.231865e-10, 
    1.217633e-10, 1.208225e-10, 1.201571e-10, 1.20251e-10, 1.204302e-10, 
    1.213534e-10, 1.222244e-10, 1.228903e-10, 1.233366e-10, 1.237772e-10, 
    1.251154e-10, 1.258265e-10, 1.274259e-10, 1.271366e-10, 1.276269e-10, 
    1.280963e-10, 1.288861e-10, 1.287559e-10, 1.291045e-10, 1.27614e-10, 
    1.286036e-10, 1.269719e-10, 1.274172e-10, 1.23897e-10, 1.225687e-10, 
    1.22006e-10, 1.215147e-10, 1.203233e-10, 1.211454e-10, 1.20821e-10, 
    1.215936e-10, 1.220857e-10, 1.218422e-10, 1.233489e-10, 1.22762e-10, 
    1.258687e-10, 1.24526e-10, 1.280415e-10, 1.271959e-10, 1.282446e-10, 
    1.27709e-10, 1.286273e-10, 1.278007e-10, 1.292343e-10, 1.295475e-10, 
    1.293334e-10, 1.301567e-10, 1.277549e-10, 1.286747e-10, 1.218354e-10, 
    1.218751e-10, 1.220601e-10, 1.212477e-10, 1.211981e-10, 1.204562e-10, 
    1.211163e-10, 1.213979e-10, 1.221143e-10, 1.225389e-10, 1.229433e-10, 
    1.238347e-10, 1.248338e-10, 1.262375e-10, 1.272507e-10, 1.27932e-10, 
    1.27514e-10, 1.27883e-10, 1.274706e-10, 1.272775e-10, 1.294301e-10, 
    1.282192e-10, 1.300381e-10, 1.299372e-10, 1.291127e-10, 1.299485e-10, 
    1.219029e-10, 1.216746e-10, 1.208832e-10, 1.215023e-10, 1.203755e-10, 
    1.210056e-10, 1.213686e-10, 1.227742e-10, 1.230842e-10, 1.233719e-10, 
    1.23941e-10, 1.246733e-10, 1.259629e-10, 1.270902e-10, 1.281236e-10, 
    1.280478e-10, 1.280745e-10, 1.283058e-10, 1.277331e-10, 1.283999e-10, 
    1.28512e-10, 1.282191e-10, 1.299236e-10, 1.294355e-10, 1.29935e-10, 
    1.296171e-10, 1.217488e-10, 1.221333e-10, 1.219254e-10, 1.223164e-10, 
    1.220409e-10, 1.232683e-10, 1.236375e-10, 1.253721e-10, 1.246589e-10, 
    1.25795e-10, 1.24774e-10, 1.249546e-10, 1.258321e-10, 1.248291e-10, 
    1.270279e-10, 1.255351e-10, 1.283148e-10, 1.268167e-10, 1.28409e-10, 
    1.281191e-10, 1.285992e-10, 1.290298e-10, 1.295726e-10, 1.30577e-10, 
    1.303441e-10, 1.311862e-10, 1.227076e-10, 1.232084e-10, 1.231643e-10, 
    1.236893e-10, 1.240783e-10, 1.249234e-10, 1.262847e-10, 1.257719e-10, 
    1.26714e-10, 1.269035e-10, 1.254726e-10, 1.263502e-10, 1.235441e-10, 
    1.239954e-10, 1.237266e-10, 1.227471e-10, 1.2589e-10, 1.242722e-10, 
    1.272674e-10, 1.263852e-10, 1.289684e-10, 1.276805e-10, 1.30216e-10, 
    1.313071e-10, 1.323382e-10, 1.335479e-10, 1.234821e-10, 1.231414e-10, 
    1.237518e-10, 1.245987e-10, 1.253871e-10, 1.264389e-10, 1.265468e-10, 
    1.267444e-10, 1.272569e-10, 1.276886e-10, 1.268068e-10, 1.277969e-10, 
    1.241001e-10, 1.260309e-10, 1.230127e-10, 1.239178e-10, 1.245487e-10, 
    1.242718e-10, 1.257134e-10, 1.260544e-10, 1.274444e-10, 1.267249e-10, 
    1.310374e-10, 1.291208e-10, 1.344726e-10, 1.329665e-10, 1.230225e-10, 
    1.23481e-10, 1.250831e-10, 1.243196e-10, 1.265093e-10, 1.270511e-10, 
    1.274924e-10, 1.280576e-10, 1.281187e-10, 1.284542e-10, 1.279046e-10, 
    1.284324e-10, 1.264411e-10, 1.273291e-10, 1.248995e-10, 1.254888e-10, 
    1.252175e-10, 1.249203e-10, 1.258387e-10, 1.268207e-10, 1.268417e-10, 
    1.271574e-10, 1.280489e-10, 1.265182e-10, 1.312856e-10, 1.283313e-10, 
    1.239819e-10, 1.24869e-10, 1.24996e-10, 1.246518e-10, 1.269967e-10, 
    1.261446e-10, 1.28446e-10, 1.27822e-10, 1.288451e-10, 1.283362e-10, 
    1.282615e-10, 1.276095e-10, 1.272044e-10, 1.261836e-10, 1.253561e-10, 
    1.247017e-10, 1.248538e-10, 1.25573e-10, 1.268809e-10, 1.281242e-10, 
    1.278513e-10, 1.287672e-10, 1.263499e-10, 1.273608e-10, 1.269696e-10, 
    1.279909e-10, 1.257583e-10, 1.276581e-10, 1.252749e-10, 1.25483e-10, 
    1.261278e-10, 1.274295e-10, 1.277184e-10, 1.280272e-10, 1.278366e-10, 
    1.269142e-10, 1.267634e-10, 1.261121e-10, 1.259325e-10, 1.254377e-10, 
    1.250287e-10, 1.254023e-10, 1.257953e-10, 1.269146e-10, 1.279273e-10, 
    1.290359e-10, 1.29308e-10, 1.306103e-10, 1.295496e-10, 1.313022e-10, 
    1.298114e-10, 1.323973e-10, 1.277687e-10, 1.297677e-10, 1.261572e-10, 
    1.265438e-10, 1.272445e-10, 1.288587e-10, 1.279861e-10, 1.290069e-10, 
    1.267575e-10, 1.255979e-10, 1.252987e-10, 1.247415e-10, 1.253115e-10, 
    1.252651e-10, 1.258116e-10, 1.256359e-10, 1.269518e-10, 1.262441e-10, 
    1.282596e-10, 1.289989e-10, 1.310978e-10, 1.323926e-10, 1.337169e-10, 
    1.343036e-10, 1.344824e-10, 1.345572e-10,
  1.315679e-10, 1.327967e-10, 1.325573e-10, 1.335522e-10, 1.329998e-10, 
    1.33652e-10, 1.318165e-10, 1.328456e-10, 1.321881e-10, 1.316783e-10, 
    1.354951e-10, 1.335966e-10, 1.374835e-10, 1.362606e-10, 1.393445e-10, 
    1.372928e-10, 1.397603e-10, 1.39285e-10, 1.407184e-10, 1.403068e-10, 
    1.421496e-10, 1.409085e-10, 1.431103e-10, 1.418526e-10, 1.42049e-10, 
    1.408677e-10, 1.339774e-10, 1.352579e-10, 1.339018e-10, 1.340839e-10, 
    1.340021e-10, 1.330112e-10, 1.325134e-10, 1.314743e-10, 1.316626e-10, 
    1.324259e-10, 1.341658e-10, 1.335737e-10, 1.350688e-10, 1.350349e-10, 
    1.367105e-10, 1.359536e-10, 1.387878e-10, 1.379788e-10, 1.40324e-10, 
    1.39732e-10, 1.402962e-10, 1.40125e-10, 1.402984e-10, 1.394308e-10, 
    1.398022e-10, 1.390401e-10, 1.360951e-10, 1.369569e-10, 1.343961e-10, 
    1.328699e-10, 1.318615e-10, 1.311487e-10, 1.312494e-10, 1.314414e-10, 
    1.324304e-10, 1.333641e-10, 1.340783e-10, 1.345572e-10, 1.350301e-10, 
    1.364673e-10, 1.372315e-10, 1.389517e-10, 1.386403e-10, 1.39168e-10, 
    1.396732e-10, 1.405239e-10, 1.403836e-10, 1.407592e-10, 1.391541e-10, 
    1.402196e-10, 1.384631e-10, 1.389423e-10, 1.351589e-10, 1.337333e-10, 
    1.331301e-10, 1.326033e-10, 1.313268e-10, 1.322076e-10, 1.3186e-10, 
    1.326878e-10, 1.332154e-10, 1.329543e-10, 1.345703e-10, 1.339407e-10, 
    1.372769e-10, 1.358341e-10, 1.396143e-10, 1.387042e-10, 1.398329e-10, 
    1.392563e-10, 1.402451e-10, 1.39355e-10, 1.40899e-10, 1.412366e-10, 
    1.410059e-10, 1.418933e-10, 1.393057e-10, 1.402962e-10, 1.32947e-10, 
    1.329895e-10, 1.331879e-10, 1.323172e-10, 1.32264e-10, 1.314691e-10, 
    1.321763e-10, 1.324781e-10, 1.33246e-10, 1.337014e-10, 1.341352e-10, 
    1.350917e-10, 1.361647e-10, 1.376733e-10, 1.387631e-10, 1.394964e-10, 
    1.390465e-10, 1.394436e-10, 1.389997e-10, 1.387919e-10, 1.411101e-10, 
    1.398056e-10, 1.417655e-10, 1.416566e-10, 1.407681e-10, 1.416689e-10, 
    1.330194e-10, 1.327746e-10, 1.319266e-10, 1.325899e-10, 1.313827e-10, 
    1.320577e-10, 1.324467e-10, 1.339539e-10, 1.342863e-10, 1.34595e-10, 
    1.352059e-10, 1.359922e-10, 1.373781e-10, 1.385905e-10, 1.397027e-10, 
    1.39621e-10, 1.396497e-10, 1.398989e-10, 1.392823e-10, 1.400002e-10, 
    1.40121e-10, 1.398055e-10, 1.41642e-10, 1.411159e-10, 1.416543e-10, 
    1.413116e-10, 1.328541e-10, 1.332664e-10, 1.330435e-10, 1.334628e-10, 
    1.331674e-10, 1.34484e-10, 1.348802e-10, 1.367431e-10, 1.359768e-10, 
    1.371976e-10, 1.361005e-10, 1.362945e-10, 1.372376e-10, 1.361596e-10, 
    1.385235e-10, 1.369183e-10, 1.399085e-10, 1.382964e-10, 1.400099e-10, 
    1.396978e-10, 1.402148e-10, 1.406787e-10, 1.412637e-10, 1.423467e-10, 
    1.420954e-10, 1.430039e-10, 1.338824e-10, 1.344196e-10, 1.343722e-10, 
    1.349357e-10, 1.353533e-10, 1.362609e-10, 1.37724e-10, 1.371727e-10, 
    1.381857e-10, 1.383896e-10, 1.36851e-10, 1.377945e-10, 1.347799e-10, 
    1.352643e-10, 1.349758e-10, 1.339247e-10, 1.372997e-10, 1.355616e-10, 
    1.387811e-10, 1.378321e-10, 1.406125e-10, 1.392257e-10, 1.419573e-10, 
    1.431345e-10, 1.442476e-10, 1.455549e-10, 1.347133e-10, 1.343477e-10, 
    1.350028e-10, 1.359122e-10, 1.367591e-10, 1.378898e-10, 1.380058e-10, 
    1.382184e-10, 1.387697e-10, 1.392343e-10, 1.382856e-10, 1.393509e-10, 
    1.353769e-10, 1.374511e-10, 1.342096e-10, 1.35181e-10, 1.358585e-10, 
    1.355611e-10, 1.371098e-10, 1.374763e-10, 1.389716e-10, 1.381974e-10, 
    1.428434e-10, 1.407769e-10, 1.465548e-10, 1.449264e-10, 1.342201e-10, 
    1.347121e-10, 1.364325e-10, 1.356124e-10, 1.379655e-10, 1.385483e-10, 
    1.390232e-10, 1.396316e-10, 1.396973e-10, 1.400586e-10, 1.394669e-10, 
    1.400352e-10, 1.378923e-10, 1.388475e-10, 1.362352e-10, 1.368684e-10, 
    1.365769e-10, 1.362576e-10, 1.372445e-10, 1.383005e-10, 1.383231e-10, 
    1.386628e-10, 1.396226e-10, 1.379751e-10, 1.431115e-10, 1.399266e-10, 
    1.352498e-10, 1.362026e-10, 1.36339e-10, 1.359692e-10, 1.384898e-10, 
    1.375734e-10, 1.400498e-10, 1.39378e-10, 1.404797e-10, 1.399316e-10, 
    1.398511e-10, 1.391492e-10, 1.387132e-10, 1.376154e-10, 1.367258e-10, 
    1.360228e-10, 1.361861e-10, 1.36959e-10, 1.383653e-10, 1.397033e-10, 
    1.394096e-10, 1.403958e-10, 1.377941e-10, 1.388816e-10, 1.384607e-10, 
    1.395598e-10, 1.371581e-10, 1.392018e-10, 1.366385e-10, 1.368622e-10, 
    1.375553e-10, 1.389556e-10, 1.392665e-10, 1.395989e-10, 1.393937e-10, 
    1.384011e-10, 1.382388e-10, 1.375384e-10, 1.373454e-10, 1.368135e-10, 
    1.36374e-10, 1.367755e-10, 1.371979e-10, 1.384015e-10, 1.394914e-10, 
    1.406853e-10, 1.409784e-10, 1.423828e-10, 1.41239e-10, 1.431294e-10, 
    1.415214e-10, 1.443117e-10, 1.393208e-10, 1.414742e-10, 1.375868e-10, 
    1.380026e-10, 1.387565e-10, 1.404945e-10, 1.395546e-10, 1.406541e-10, 
    1.382325e-10, 1.369857e-10, 1.366642e-10, 1.360655e-10, 1.366779e-10, 
    1.36628e-10, 1.372154e-10, 1.370264e-10, 1.384415e-10, 1.376804e-10, 
    1.398491e-10, 1.406454e-10, 1.429086e-10, 1.443064e-10, 1.457375e-10, 
    1.46372e-10, 1.465654e-10, 1.466463e-10,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GC_HEAT1 =
  24573.48, 24593.75, 24589.78, 24606.36, 24597.13, 24608.04, 24577.56, 
    24594.57, 24583.67, 24575.29, 24639.27, 24607.11, 24673.71, 24652.42, 
    24706.31, 24670.37, 24713.7, 24705.26, 24730.89, 24723.48, 24757.06, 
    24734.34, 24774.97, 24751.58, 24755.21, 24733.6, 24613.51, 24635.23, 
    24612.24, 24615.31, 24613.93, 24597.32, 24589.05, 24571.95, 24575.03, 
    24587.6, 24616.69, 24606.72, 24632, 24631.43, 24660.21, 24647.13, 
    24696.49, 24682.36, 24723.79, 24713.19, 24723.29, 24720.21, 24723.32, 
    24707.84, 24714.44, 24700.93, 24649.57, 24664.5, 24620.59, 24594.97, 
    24578.3, 24566.63, 24568.27, 24571.41, 24587.68, 24603.21, 24615.21, 
    24623.32, 24631.34, 24656, 24669.29, 24699.38, 24693.9, 24703.19, 
    24712.15, 24727.38, 24724.86, 24731.63, 24702.94, 24721.91, 24690.8, 
    24699.21, 24633.54, 24609.4, 24599.31, 24590.54, 24569.54, 24584, 
    24578.27, 24591.94, 24600.73, 24596.38, 24623.54, 24612.89, 24670.09, 
    24645.08, 24711.1, 24695.02, 24714.99, 24704.75, 24722.37, 24706.5, 
    24734.17, 24740.3, 24736.1, 24752.33, 24705.62, 24723.29, 24596.25, 
    24596.96, 24600.27, 24585.81, 24584.93, 24571.86, 24583.48, 24588.47, 
    24601.24, 24608.87, 24616.17, 24632.39, 24650.77, 24677.04, 24696.06, 
    24709, 24701.04, 24708.07, 24700.22, 24696.56, 24738, 24714.51, 24749.98, 
    24747.98, 24731.79, 24748.21, 24597.46, 24593.38, 24579.37, 24590.32, 
    24570.45, 24581.53, 24587.95, 24613.12, 24618.73, 24623.96, 24634.33, 
    24647.79, 24671.86, 24693.03, 24712.67, 24711.22, 24711.73, 24716.17, 
    24705.21, 24717.98, 24720.14, 24714.5, 24747.71, 24738.1, 24747.94, 
    24741.67, 24594.71, 24601.58, 24597.86, 24604.87, 24599.93, 24622.08, 
    24628.8, 24660.78, 24647.53, 24668.7, 24649.66, 24653.01, 24669.4, 
    24650.68, 24691.86, 24663.83, 24716.34, 24687.89, 24718.15, 24712.58, 
    24721.82, 24730.18, 24740.79, 24760.71, 24756.06, 24772.97, 24611.91, 
    24620.99, 24620.18, 24629.74, 24636.85, 24652.43, 24677.93, 24668.26, 
    24685.96, 24689.52, 24662.66, 24679.17, 24627.1, 24635.33, 24630.42, 
    24612.62, 24670.48, 24640.41, 24696.37, 24679.82, 24728.98, 24704.21, 
    24753.51, 24775.42, 24796.51, 24821.57, 24625.97, 24619.77, 24630.88, 
    24646.42, 24661.06, 24680.82, 24682.83, 24686.53, 24696.17, 24704.36, 
    24687.7, 24706.42, 24637.25, 24673.14, 24617.43, 24633.91, 24645.5, 
    24640.4, 24667.17, 24673.58, 24699.72, 24686.16, 24769.97, 24731.96, 
    24840.86, 24809.54, 24617.61, 24625.95, 24655.39, 24641.28, 24682.13, 
    24692.29, 24700.63, 24711.41, 24712.57, 24719.03, 24708.48, 24718.61, 
    24680.86, 24697.54, 24651.98, 24662.96, 24657.89, 24652.37, 24669.52, 
    24687.96, 24688.35, 24694.3, 24711.25, 24682.3, 24775, 24716.67, 
    24635.08, 24651.42, 24653.78, 24647.4, 24691.27, 24675.28, 24718.87, 
    24706.9, 24726.59, 24716.75, 24715.32, 24702.86, 24695.18, 24676.02, 
    24660.48, 24648.32, 24651.13, 24664.54, 24689.09, 24712.68, 24707.46, 
    24725.08, 24679.16, 24698.14, 24690.76, 24710.13, 24668.01, 24703.79, 
    24658.96, 24662.85, 24674.96, 24699.44, 24704.93, 24710.82, 24707.18, 
    24689.72, 24686.88, 24674.67, 24671.28, 24662, 24654.38, 24661.34, 
    24668.71, 24689.72, 24708.91, 24730.3, 24735.61, 24761.39, 24740.35, 
    24775.33, 24745.51, 24797.74, 24705.89, 24744.64, 24675.52, 24682.77, 
    24695.94, 24726.86, 24710.04, 24729.73, 24686.77, 24665, 24659.41, 
    24649.05, 24659.65, 24658.78, 24669.01, 24665.71, 24690.42, 24677.16, 
    24715.28, 24729.58, 24771.18, 24797.64, 24825.07, 24837.31, 24841.06, 
    24842.64 ;

 GC_ICE1 =
  17682.08, 17714.56, 17708.19, 17734.75, 17719.97, 17737.43, 17688.61, 
    17715.86, 17698.41, 17684.98, 17787.43, 17735.94, 17842.51, 17808.46, 
    17894.55, 17837.17, 17906.34, 17892.87, 17933.77, 17921.94, 17975.51, 
    17939.26, 18004.06, 17966.77, 17972.55, 17938.08, 17746.2, 17780.96, 
    17744.16, 17749.07, 17746.86, 17720.27, 17707.03, 17679.62, 17684.56, 
    17704.71, 17751.29, 17735.33, 17775.8, 17774.88, 17820.93, 17800, 
    17878.88, 17856.34, 17922.43, 17905.53, 17921.63, 17916.73, 17921.7, 
    17896.99, 17907.53, 17885.97, 17803.9, 17827.79, 17757.53, 17716.51, 
    17689.8, 17671.11, 17673.74, 17678.76, 17704.83, 17729.71, 17748.92, 
    17761.9, 17774.74, 17814.19, 17835.45, 17883.48, 17874.75, 17889.57, 
    17903.86, 17928.17, 17924.14, 17934.95, 17889.18, 17919.44, 17869.8, 
    17883.22, 17778.26, 17739.62, 17723.45, 17709.41, 17675.77, 17698.93, 
    17689.76, 17711.66, 17725.72, 17718.75, 17762.26, 17745.21, 17836.72, 
    17796.71, 17902.19, 17876.54, 17908.4, 17892.06, 17920.17, 17894.85, 
    17938.99, 17948.78, 17942.08, 17967.97, 17893.46, 17921.63, 17718.56, 
    17719.7, 17724.99, 17701.83, 17700.42, 17679.49, 17698.1, 17706.09, 
    17726.54, 17738.76, 17750.46, 17776.42, 17805.82, 17847.84, 17878.19, 
    17898.85, 17886.15, 17897.35, 17884.83, 17879, 17945.1, 17907.63, 
    17964.21, 17961.03, 17935.21, 17961.38, 17720.49, 17713.97, 17691.51, 
    17709.06, 17677.23, 17694.97, 17705.26, 17745.56, 17754.55, 17762.93, 
    17779.53, 17801.06, 17839.55, 17873.36, 17904.7, 17902.38, 17903.2, 
    17910.28, 17892.79, 17913.17, 17916.62, 17907.62, 17960.6, 17945.27, 
    17960.96, 17950.96, 17716.08, 17727.09, 17721.13, 17732.35, 17724.44, 
    17759.92, 17770.68, 17821.84, 17800.64, 17834.5, 17804.04, 17809.4, 
    17835.62, 17805.67, 17871.49, 17826.72, 17910.55, 17865.16, 17913.45, 
    17904.56, 17919.3, 17932.63, 17949.56, 17981.33, 17973.91, 18000.88, 
    17743.63, 17758.17, 17756.88, 17772.18, 17783.55, 17808.47, 17849.26, 
    17833.81, 17862.08, 17867.75, 17824.84, 17851.24, 17767.96, 17781.12, 
    17773.27, 17744.77, 17837.36, 17789.24, 17878.7, 17852.28, 17930.72, 
    17891.2, 17969.85, 18004.79, 18038.41, 18078.31, 17766.15, 17756.21, 
    17774, 17798.86, 17822.29, 17853.88, 17857.09, 17862.99, 17878.38, 
    17891.44, 17864.86, 17894.73, 17784.2, 17841.6, 17752.47, 17778.86, 
    17797.39, 17789.23, 17832.05, 17842.3, 17884.04, 17862.4, 17996.09, 
    17935.46, 18108.97, 18059.19, 17752.75, 17766.12, 17813.22, 17790.63, 
    17855.97, 17872.18, 17885.49, 17902.68, 17904.55, 17914.84, 17898.01, 
    17914.17, 17853.94, 17880.56, 17807.76, 17825.33, 17817.22, 17808.38, 
    17835.81, 17865.28, 17865.9, 17875.38, 17902.44, 17856.23, 18004.11, 
    17911.08, 17780.72, 17806.87, 17810.63, 17800.43, 17870.55, 17845.03, 
    17914.58, 17895.5, 17926.9, 17911.21, 17908.92, 17889.04, 17876.79, 
    17846.21, 17821.36, 17801.9, 17806.4, 17827.85, 17867.08, 17904.72, 
    17896.39, 17924.49, 17851.23, 17881.52, 17869.74, 17900.64, 17833.4, 
    17890.53, 17818.93, 17825.15, 17844.52, 17883.6, 17892.35, 17901.75, 
    17895.94, 17868.08, 17863.56, 17844.04, 17838.63, 17823.79, 17811.6, 
    17822.74, 17834.51, 17868.09, 17898.71, 17932.82, 17941.29, 17982.4, 
    17948.85, 18004.64, 17957.09, 18040.37, 17893.88, 17955.7, 17845.4, 
    17857, 17878.01, 17927.33, 17900.5, 17931.92, 17863.38, 17828.59, 
    17819.64, 17803.08, 17820.02, 17818.64, 17835, 17829.72, 17869.2, 
    17848.03, 17908.86, 17931.67, 17998.03, 18040.21, 18083.88, 18103.33, 
    18109.29, 18111.79 ;

 GC_LIQ1 =
  5232.649, 5234.678, 5234.28, 5235.941, 5235.016, 5236.109, 5233.057, 
    5234.759, 5233.669, 5232.83, 5239.249, 5236.016, 5242.728, 5240.577, 
    5246.078, 5242.39, 5246.839, 5245.969, 5248.612, 5247.847, 5251.313, 
    5248.967, 5253.162, 5250.747, 5251.121, 5248.891, 5236.657, 5238.841, 
    5236.53, 5236.837, 5236.699, 5235.035, 5234.207, 5232.496, 5232.804, 
    5234.062, 5236.976, 5235.977, 5238.515, 5238.457, 5241.364, 5240.042, 
    5245.065, 5243.61, 5247.879, 5246.787, 5247.827, 5247.51, 5247.832, 
    5246.235, 5246.916, 5245.523, 5240.288, 5241.797, 5237.367, 5234.8, 
    5233.131, 5231.964, 5232.128, 5232.442, 5234.07, 5235.625, 5236.828, 
    5237.641, 5238.449, 5240.938, 5242.282, 5245.362, 5244.799, 5245.756, 
    5246.679, 5248.25, 5247.989, 5248.688, 5245.73, 5247.686, 5244.479, 
    5245.345, 5238.67, 5236.246, 5235.234, 5234.356, 5232.255, 5233.701, 
    5233.128, 5234.497, 5235.376, 5234.94, 5237.663, 5236.595, 5242.362, 
    5239.835, 5246.571, 5244.914, 5246.972, 5245.916, 5247.733, 5246.096, 
    5248.949, 5249.583, 5249.149, 5250.824, 5246.006, 5247.827, 5234.928, 
    5234.999, 5235.33, 5233.882, 5233.794, 5232.487, 5233.649, 5234.148, 
    5235.427, 5236.192, 5236.924, 5238.555, 5240.41, 5243.065, 5245.021, 
    5246.354, 5245.534, 5246.258, 5245.45, 5245.073, 5249.345, 5246.922, 
    5250.582, 5250.375, 5248.705, 5250.398, 5235.049, 5234.641, 5233.238, 
    5234.334, 5232.346, 5233.454, 5234.097, 5236.618, 5237.181, 5237.706, 
    5238.75, 5240.109, 5242.541, 5244.709, 5246.733, 5246.583, 5246.636, 
    5247.093, 5245.964, 5247.28, 5247.503, 5246.921, 5250.348, 5249.356, 
    5250.371, 5249.724, 5234.773, 5235.461, 5235.089, 5235.791, 5235.296, 
    5237.517, 5238.192, 5241.421, 5240.083, 5242.222, 5240.297, 5240.636, 
    5242.292, 5240.4, 5244.588, 5241.729, 5247.111, 5244.18, 5247.298, 
    5246.724, 5247.676, 5248.538, 5249.633, 5251.689, 5251.209, 5252.956, 
    5236.497, 5237.407, 5237.326, 5238.287, 5239.004, 5240.577, 5243.155, 
    5242.178, 5243.98, 5244.347, 5241.61, 5243.281, 5238.021, 5238.852, 
    5238.356, 5236.568, 5242.402, 5239.364, 5245.053, 5243.348, 5248.415, 
    5245.861, 5250.946, 5253.209, 5255.39, 5258.008, 5237.907, 5237.285, 
    5238.402, 5239.971, 5241.449, 5243.451, 5243.659, 5244.039, 5245.033, 
    5245.876, 5244.16, 5246.089, 5239.045, 5242.67, 5237.05, 5238.708, 
    5239.877, 5239.362, 5242.066, 5242.715, 5245.398, 5244.001, 5252.646, 
    5248.721, 5260.053, 5256.742, 5237.068, 5237.905, 5240.877, 5239.451, 
    5243.586, 5244.633, 5245.492, 5246.603, 5246.723, 5247.388, 5246.301, 
    5247.345, 5243.456, 5245.173, 5240.532, 5241.641, 5241.129, 5240.571, 
    5242.304, 5244.187, 5244.228, 5244.839, 5246.586, 5243.604, 5253.165, 
    5247.145, 5238.826, 5240.476, 5240.713, 5240.069, 5244.527, 5242.888, 
    5247.372, 5246.138, 5248.167, 5247.154, 5247.005, 5245.721, 5244.931, 
    5242.962, 5241.391, 5240.163, 5240.446, 5241.8, 5244.303, 5246.734, 
    5246.196, 5248.012, 5243.28, 5245.235, 5244.475, 5246.471, 5242.152, 
    5245.818, 5241.237, 5241.63, 5242.855, 5245.37, 5245.935, 5246.542, 
    5246.167, 5244.368, 5244.076, 5242.825, 5242.483, 5241.544, 5240.774, 
    5241.478, 5242.222, 5244.368, 5246.346, 5248.55, 5249.098, 5251.759, 
    5249.587, 5253.199, 5250.12, 5255.518, 5246.034, 5250.031, 5242.911, 
    5243.653, 5245.009, 5248.195, 5246.461, 5248.492, 5244.064, 5241.848, 
    5241.282, 5240.237, 5241.306, 5241.219, 5242.253, 5241.919, 5244.44, 
    5243.078, 5247.002, 5248.476, 5252.771, 5255.507, 5258.378, 5259.676, 
    5260.075, 5260.242 ;

 GPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 GROSS_NMIN =
  8.721962e-09, 8.760422e-09, 8.752946e-09, 8.783966e-09, 8.766759e-09, 
    8.787071e-09, 8.72976e-09, 8.761948e-09, 8.7414e-09, 8.725426e-09, 
    8.844167e-09, 8.785351e-09, 8.905277e-09, 8.867761e-09, 8.962011e-09, 
    8.899439e-09, 8.974629e-09, 8.960209e-09, 9.003618e-09, 8.991182e-09, 
    9.046705e-09, 9.009359e-09, 9.075491e-09, 9.037787e-09, 9.043684e-09, 
    9.008126e-09, 8.797189e-09, 8.836844e-09, 8.794839e-09, 8.800494e-09, 
    8.797957e-09, 8.767114e-09, 8.75157e-09, 8.719024e-09, 8.724933e-09, 
    8.748838e-09, 8.803037e-09, 8.78464e-09, 8.83101e-09, 8.829963e-09, 
    8.881588e-09, 8.858311e-09, 8.945088e-09, 8.920424e-09, 8.991701e-09, 
    8.973775e-09, 8.990859e-09, 8.985679e-09, 8.990926e-09, 8.964635e-09, 
    8.975899e-09, 8.952767e-09, 8.86267e-09, 8.889146e-09, 8.810181e-09, 
    8.762701e-09, 8.731171e-09, 8.708796e-09, 8.71196e-09, 8.717989e-09, 
    8.748978e-09, 8.778116e-09, 8.800321e-09, 8.815175e-09, 8.829812e-09, 
    8.874111e-09, 8.897564e-09, 8.950074e-09, 8.9406e-09, 8.956653e-09, 
    8.971992e-09, 8.997742e-09, 8.993504e-09, 9.004849e-09, 8.95623e-09, 
    8.988541e-09, 8.935203e-09, 8.94979e-09, 8.833783e-09, 8.789603e-09, 
    8.770819e-09, 8.754382e-09, 8.714392e-09, 8.742008e-09, 8.731121e-09, 
    8.757023e-09, 8.773481e-09, 8.765341e-09, 8.815582e-09, 8.796049e-09, 
    8.898954e-09, 8.854627e-09, 8.970202e-09, 8.942544e-09, 8.976832e-09, 
    8.959336e-09, 8.989314e-09, 8.962334e-09, 9.009072e-09, 9.019248e-09, 
    9.012294e-09, 9.039011e-09, 8.960838e-09, 8.990858e-09, 8.765113e-09, 
    8.766441e-09, 8.772626e-09, 8.745437e-09, 8.743775e-09, 8.718861e-09, 
    8.741029e-09, 8.750469e-09, 8.774436e-09, 8.788612e-09, 8.802087e-09, 
    8.831718e-09, 8.864809e-09, 8.911087e-09, 8.944338e-09, 8.966627e-09, 
    8.952959e-09, 8.965025e-09, 8.951537e-09, 8.945215e-09, 9.015435e-09, 
    8.976004e-09, 9.035169e-09, 9.031895e-09, 9.005118e-09, 9.032264e-09, 
    8.767373e-09, 8.759733e-09, 8.733209e-09, 8.753966e-09, 8.716149e-09, 
    8.737316e-09, 8.749487e-09, 8.796456e-09, 8.806778e-09, 8.816346e-09, 
    8.835246e-09, 8.859502e-09, 8.902054e-09, 8.939081e-09, 8.972885e-09, 
    8.970408e-09, 8.97128e-09, 8.97883e-09, 8.960125e-09, 8.981901e-09, 
    8.985555e-09, 8.976e-09, 9.031456e-09, 9.015613e-09, 9.031825e-09, 
    9.02151e-09, 8.762217e-09, 8.775071e-09, 8.768126e-09, 8.781187e-09, 
    8.771985e-09, 8.812903e-09, 8.825173e-09, 8.882585e-09, 8.859024e-09, 
    8.896524e-09, 8.862834e-09, 8.868803e-09, 8.897745e-09, 8.864655e-09, 
    8.937038e-09, 8.887961e-09, 8.979124e-09, 8.93011e-09, 8.982195e-09, 
    8.972738e-09, 8.988397e-09, 9.002421e-09, 9.020066e-09, 9.052621e-09, 
    9.045082e-09, 9.07231e-09, 8.794236e-09, 8.810909e-09, 8.809443e-09, 
    8.826892e-09, 8.839797e-09, 8.867771e-09, 8.912638e-09, 8.895766e-09, 
    8.926742e-09, 8.93296e-09, 8.885901e-09, 8.914792e-09, 8.822069e-09, 
    8.837048e-09, 8.82813e-09, 8.795551e-09, 8.899652e-09, 8.846224e-09, 
    8.944887e-09, 8.915942e-09, 9.000421e-09, 8.958406e-09, 9.040932e-09, 
    9.076211e-09, 9.109422e-09, 9.148227e-09, 8.82001e-09, 8.808681e-09, 
    8.828968e-09, 8.857034e-09, 8.88308e-09, 8.917707e-09, 8.92125e-09, 
    8.927737e-09, 8.944541e-09, 8.958669e-09, 8.929787e-09, 8.962211e-09, 
    8.840519e-09, 8.904291e-09, 8.804397e-09, 8.834474e-09, 8.85538e-09, 
    8.846211e-09, 8.893839e-09, 8.905063e-09, 8.95068e-09, 8.927099e-09, 
    9.067502e-09, 9.005381e-09, 9.177779e-09, 9.129597e-09, 8.804722e-09, 
    8.819972e-09, 8.873046e-09, 8.847794e-09, 8.920019e-09, 8.937797e-09, 
    8.952251e-09, 8.970726e-09, 8.972722e-09, 8.983669e-09, 8.965731e-09, 
    8.982961e-09, 8.91778e-09, 8.946908e-09, 8.866982e-09, 8.886434e-09, 
    8.877485e-09, 8.867669e-09, 8.897965e-09, 8.930241e-09, 8.930932e-09, 
    8.941282e-09, 8.970442e-09, 8.920312e-09, 9.075516e-09, 8.979659e-09, 
    8.836602e-09, 8.865973e-09, 8.870171e-09, 8.858793e-09, 8.936015e-09, 
    8.908033e-09, 8.983402e-09, 8.963033e-09, 8.996409e-09, 8.979824e-09, 
    8.977383e-09, 8.956082e-09, 8.94282e-09, 8.909316e-09, 8.882057e-09, 
    8.860443e-09, 8.865469e-09, 8.889211e-09, 8.932216e-09, 8.972902e-09, 
    8.96399e-09, 8.993872e-09, 8.914782e-09, 8.947944e-09, 8.935126e-09, 
    8.968549e-09, 8.895317e-09, 8.957672e-09, 8.879379e-09, 8.886244e-09, 
    8.907478e-09, 8.950192e-09, 8.959645e-09, 8.969735e-09, 8.96351e-09, 
    8.933308e-09, 8.928361e-09, 8.906962e-09, 8.901053e-09, 8.884749e-09, 
    8.87125e-09, 8.883584e-09, 8.896535e-09, 8.933322e-09, 8.966474e-09, 
    9.00262e-09, 9.011467e-09, 9.053698e-09, 9.019318e-09, 9.07605e-09, 
    9.027812e-09, 9.11132e-09, 8.961289e-09, 9.026397e-09, 8.908445e-09, 
    8.921152e-09, 8.944133e-09, 8.99685e-09, 8.968392e-09, 9.001675e-09, 
    8.928168e-09, 8.89003e-09, 8.880165e-09, 8.861757e-09, 8.880586e-09, 
    8.879055e-09, 8.897072e-09, 8.891282e-09, 8.934543e-09, 8.911305e-09, 
    8.977321e-09, 9.001413e-09, 9.069456e-09, 9.11117e-09, 9.153638e-09, 
    9.172386e-09, 9.178093e-09, 9.180479e-09 ;

 H2OCAN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSNO_TOP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 H2OSOI =
  6.171655, 6.200645, 6.195002, 6.218437, 6.205429, 6.220785, 6.177525, 
    6.201798, 6.186295, 6.174261, 6.264087, 6.219483, 6.310639, 6.282028, 
    6.354062, 6.306181, 6.363744, 6.352676, 6.386025, 6.376459, 6.419241, 
    6.390443, 6.441489, 6.412355, 6.416908, 6.389494, 6.228442, 6.258523, 
    6.226663, 6.230945, 6.229023, 6.205698, 6.193966, 6.169443, 6.17389, 
    6.191904, 6.232872, 6.218944, 6.254083, 6.253288, 6.292562, 6.274834, 
    6.341086, 6.322209, 6.376858, 6.363086, 6.376211, 6.372229, 6.376263, 
    6.356072, 6.364718, 6.34697, 6.278152, 6.298326, 6.238285, 6.202369, 
    6.178588, 6.161751, 6.16413, 6.168665, 6.192009, 6.214011, 6.230813, 
    6.24207, 6.253174, 6.286869, 6.304749, 6.344909, 6.337648, 6.349951, 
    6.361717, 6.381505, 6.378245, 6.386973, 6.349625, 6.374431, 6.333515, 
    6.344689, 6.256199, 6.222699, 6.2085, 6.196086, 6.165959, 6.186754, 
    6.178551, 6.198078, 6.210508, 6.204358, 6.242378, 6.227578, 6.30581, 
    6.272033, 6.360344, 6.339138, 6.365433, 6.352006, 6.375024, 6.354306, 
    6.390223, 6.398062, 6.392704, 6.413299, 6.353158, 6.376212, 6.204186, 
    6.205189, 6.209861, 6.18934, 6.188086, 6.169321, 6.186015, 6.193134, 
    6.211228, 6.221949, 6.232151, 6.254622, 6.279781, 6.315075, 6.340511, 
    6.357599, 6.347117, 6.35637, 6.346027, 6.341182, 6.395124, 6.364799, 
    6.410334, 6.407809, 6.387181, 6.408093, 6.205893, 6.200123, 6.180123, 
    6.195771, 6.16728, 6.183218, 6.192395, 6.227888, 6.235704, 6.242958, 
    6.257301, 6.275741, 6.308176, 6.336486, 6.362401, 6.3605, 6.36117, 
    6.366968, 6.352612, 6.369327, 6.372136, 6.364795, 6.40747, 6.395259, 
    6.407755, 6.399802, 6.201998, 6.211709, 6.206461, 6.216333, 6.209377, 
    6.24035, 6.249656, 6.293324, 6.275377, 6.303955, 6.278276, 6.282821, 
    6.30489, 6.279662, 6.334923, 6.297424, 6.367194, 6.329623, 6.369553, 
    6.362289, 6.374318, 6.385104, 6.39869, 6.423807, 6.417985, 6.439026, 
    6.226206, 6.238837, 6.237723, 6.250958, 6.260759, 6.282034, 6.316259, 
    6.303374, 6.327041, 6.331799, 6.295849, 6.317906, 6.2473, 6.258672, 
    6.251899, 6.227202, 6.306343, 6.265645, 6.340932, 6.318783, 6.383566, 
    6.351295, 6.414782, 6.442049, 6.467774, 6.497926, 6.245737, 6.237146, 
    6.252533, 6.273865, 6.293699, 6.320133, 6.322841, 6.327803, 6.340666, 
    6.351495, 6.329373, 6.354211, 6.261313, 6.309884, 6.233901, 6.256718, 
    6.272606, 6.265632, 6.301903, 6.310472, 6.345372, 6.327314, 6.435313, 
    6.387385, 6.520941, 6.483441, 6.234147, 6.245707, 6.286054, 6.266835, 
    6.321899, 6.335503, 6.346574, 6.360747, 6.362278, 6.370686, 6.356912, 
    6.370141, 6.320189, 6.34248, 6.281433, 6.296256, 6.289433, 6.281956, 
    6.305052, 6.329721, 6.330247, 6.338171, 6.360538, 6.322123, 6.441518, 
    6.367613, 6.258329, 6.280669, 6.283863, 6.2752, 6.334138, 6.312741, 
    6.370481, 6.354842, 6.380479, 6.367731, 6.365857, 6.349511, 6.339349, 
    6.313721, 6.292919, 6.276456, 6.280281, 6.298375, 6.331232, 6.362417, 
    6.355577, 6.378528, 6.317896, 6.343275, 6.333458, 6.359075, 6.303032, 
    6.350739, 6.290877, 6.29611, 6.312316, 6.344999, 6.352243, 6.359986, 
    6.355207, 6.332067, 6.32828, 6.311922, 6.307411, 6.294971, 6.284684, 
    6.294082, 6.303962, 6.332076, 6.357483, 6.385258, 6.392066, 6.424644, 
    6.398118, 6.441931, 6.404673, 6.469255, 6.353509, 6.403576, 6.313054, 
    6.322765, 6.340357, 6.380822, 6.358954, 6.384533, 6.328132, 6.299, 
    6.291476, 6.277456, 6.291797, 6.29063, 6.304371, 6.299953, 6.333011, 
    6.315239, 6.36581, 6.38433, 6.43682, 6.469134, 6.502132, 6.516735, 
    6.521183, 6.523044,
  3.963831, 3.983115, 3.979361, 3.994949, 3.986296, 3.996511, 3.967734, 
    3.983883, 3.973569, 3.965563, 4.025311, 3.995645, 4.056252, 4.037231, 
    4.085108, 4.05329, 4.091541, 4.084184, 4.10634, 4.099986, 4.128411, 
    4.109275, 4.143185, 4.123834, 4.126859, 4.108646, 4.001601, 4.021612, 
    4.000418, 4.003267, 4.001988, 3.986476, 3.978675, 3.962357, 3.965316, 
    3.977301, 4.004549, 3.995284, 4.018651, 4.018122, 4.044233, 4.032447, 
    4.076483, 4.063938, 4.100251, 4.091101, 4.099822, 4.097176, 4.099856, 
    4.086441, 4.092185, 4.080392, 4.034654, 4.048065, 4.008148, 3.984266, 
    3.968443, 3.95724, 3.958823, 3.961841, 3.977371, 3.992003, 4.003177, 
    4.010663, 4.018046, 4.040455, 4.052337, 4.079025, 4.074197, 4.082375, 
    4.090191, 4.103339, 4.101172, 4.106972, 4.082157, 4.09864, 4.07145, 
    4.078876, 4.020068, 3.997782, 3.988343, 3.980083, 3.96004, 3.973875, 
    3.968418, 3.981406, 3.989674, 3.985583, 4.010868, 4.001027, 4.053042, 
    4.030587, 4.089279, 4.075188, 4.09266, 4.083738, 4.099034, 4.085267, 
    4.10913, 4.114339, 4.110779, 4.124459, 4.084504, 4.099823, 3.985469, 
    3.986136, 3.989243, 3.975595, 3.974761, 3.962276, 3.973383, 3.978119, 
    3.990152, 3.997283, 4.004068, 4.01901, 4.035739, 4.059198, 4.0761, 
    4.087454, 4.080489, 4.086638, 4.079765, 4.076546, 4.112388, 4.09224, 
    4.122489, 4.120812, 4.10711, 4.121001, 3.986604, 3.982766, 3.969463, 
    3.979872, 3.960918, 3.971522, 3.977628, 4.001235, 4.00643, 4.011254, 
    4.020791, 4.03305, 4.054612, 4.073427, 4.090646, 4.089382, 4.089827, 
    4.09368, 4.084141, 4.095248, 4.097115, 4.092236, 4.120587, 4.112475, 
    4.120776, 4.115493, 3.984013, 3.990473, 3.986982, 3.993549, 3.988923, 
    4.009522, 4.015711, 4.044743, 4.032809, 4.051807, 4.034736, 4.037758, 
    4.052433, 4.035656, 4.072391, 4.047469, 4.09383, 4.068871, 4.095397, 
    4.090571, 4.098563, 4.10573, 4.114754, 4.131441, 4.127573, 4.141548, 
    4.000113, 4.008515, 4.007772, 4.016573, 4.02309, 4.037234, 4.059984, 
    4.051419, 4.067148, 4.070311, 4.046417, 4.06108, 4.014142, 4.021706, 
    4.0172, 4.000777, 4.053395, 4.026341, 4.076381, 4.061661, 4.104708, 
    4.083269, 4.125445, 4.143559, 4.160269, 4.179707, 4.013102, 4.007389, 
    4.01762, 4.031806, 4.044989, 4.062558, 4.064357, 4.067655, 4.076203, 
    4.083399, 4.068701, 4.085204, 4.023466, 4.055748, 4.005232, 4.020407, 
    4.030968, 4.02633, 4.05044, 4.056136, 4.079332, 4.06733, 4.139086, 
    4.107248, 4.194534, 4.17037, 4.005394, 4.013081, 4.039908, 4.02713, 
    4.063732, 4.072773, 4.080129, 4.089548, 4.090564, 4.096151, 4.086998, 
    4.095788, 4.062596, 4.077408, 4.036833, 4.046688, 4.042152, 4.037181, 
    4.052534, 4.068933, 4.069279, 4.074547, 4.08942, 4.06388, 4.143214, 
    4.094119, 4.021474, 4.03633, 4.03845, 4.03269, 4.071866, 4.057645, 
    4.096014, 4.085622, 4.102656, 4.094187, 4.092942, 4.08208, 4.075328, 
    4.058297, 4.044471, 4.033525, 4.036068, 4.048098, 4.069936, 4.090657, 
    4.086113, 4.10136, 4.061071, 4.077939, 4.071415, 4.088436, 4.051193, 
    4.082907, 4.043111, 4.04659, 4.057363, 4.079087, 4.083896, 4.089042, 
    4.085865, 4.070491, 4.067973, 4.0571, 4.054103, 4.045832, 4.038994, 
    4.045243, 4.051812, 4.070496, 4.087379, 4.105833, 4.110354, 4.132002, 
    4.11438, 4.143489, 4.118742, 4.161234, 4.084743, 4.118008, 4.057852, 
    4.064307, 4.076001, 4.102889, 4.088356, 4.105353, 4.067874, 4.048515, 
    4.04351, 4.03419, 4.043723, 4.042947, 4.052081, 4.049144, 4.071116, 
    4.059305, 4.092912, 4.105217, 4.140083, 4.16115, 4.182412, 4.191823, 
    4.194689, 4.195888,
  3.282615, 3.29986, 3.296503, 3.310447, 3.302706, 3.311845, 3.286105, 
    3.300548, 3.291322, 3.284163, 3.337622, 3.31107, 3.365334, 3.348295, 
    3.391198, 3.362681, 3.396966, 3.39037, 3.41024, 3.40454, 3.430043, 
    3.412873, 3.443305, 3.425935, 3.42865, 3.412308, 3.316399, 3.33431, 
    3.315341, 3.31789, 3.316745, 3.302867, 3.29589, 3.281297, 3.283943, 
    3.294661, 3.319037, 3.310747, 3.331659, 3.331186, 3.354567, 3.344012, 
    3.383466, 3.372221, 3.404777, 3.396571, 3.404392, 3.402019, 3.404423, 
    3.392393, 3.397544, 3.38697, 3.345988, 3.358, 3.322258, 3.30089, 
    3.286739, 3.276723, 3.278138, 3.280837, 3.294724, 3.307812, 3.31781, 
    3.324509, 3.331118, 3.351183, 3.361827, 3.385744, 3.381417, 3.388747, 
    3.395756, 3.407547, 3.405604, 3.410806, 3.388552, 3.403332, 3.378954, 
    3.385611, 3.332927, 3.312982, 3.304537, 3.297148, 3.279226, 3.291597, 
    3.286717, 3.298332, 3.305727, 3.302068, 3.324692, 3.315885, 3.362458, 
    3.342346, 3.394938, 3.382304, 3.39797, 3.38997, 3.403686, 3.39134, 
    3.412742, 3.417415, 3.414222, 3.426496, 3.390657, 3.404393, 3.301966, 
    3.302563, 3.305342, 3.293135, 3.292388, 3.281226, 3.291156, 3.295392, 
    3.306156, 3.312535, 3.318606, 3.33198, 3.346959, 3.367975, 3.383123, 
    3.393302, 3.387057, 3.39257, 3.386408, 3.383522, 3.415665, 3.397593, 
    3.424729, 3.423223, 3.41093, 3.423393, 3.302981, 3.299548, 3.287651, 
    3.296959, 3.280011, 3.289493, 3.294953, 3.316071, 3.32072, 3.325038, 
    3.333575, 3.344552, 3.363865, 3.380726, 3.396163, 3.39503, 3.395429, 
    3.398885, 3.390331, 3.40029, 3.401965, 3.397589, 3.423022, 3.415743, 
    3.423191, 3.418451, 3.300664, 3.306442, 3.303319, 3.309194, 3.305056, 
    3.323488, 3.329027, 3.355024, 3.344336, 3.361352, 3.346061, 3.348768, 
    3.361913, 3.346885, 3.379797, 3.357466, 3.399019, 3.376642, 3.400425, 
    3.396096, 3.403263, 3.409692, 3.417788, 3.432762, 3.42929, 3.441835, 
    3.315068, 3.322587, 3.321922, 3.329799, 3.335634, 3.348298, 3.368678, 
    3.361005, 3.375098, 3.377933, 3.356523, 3.36966, 3.327623, 3.334394, 
    3.33036, 3.315662, 3.362775, 3.338544, 3.383374, 3.370181, 3.408775, 
    3.389549, 3.427381, 3.443641, 3.458978, 3.476969, 3.326692, 3.321579, 
    3.330736, 3.343438, 3.355244, 3.370985, 3.372597, 3.375553, 3.383214, 
    3.389665, 3.37649, 3.391284, 3.33597, 3.364882, 3.319649, 3.333231, 
    3.342687, 3.338535, 3.360128, 3.365231, 3.38602, 3.375262, 3.439625, 
    3.411054, 3.490699, 3.468326, 3.319793, 3.326674, 3.350693, 3.339251, 
    3.372037, 3.380139, 3.386734, 3.395179, 3.39609, 3.4011, 3.392892, 
    3.400775, 3.371019, 3.384295, 3.347939, 3.356766, 3.352703, 3.348251, 
    3.362003, 3.376698, 3.377009, 3.38173, 3.395064, 3.37217, 3.443331, 
    3.399278, 3.334187, 3.347489, 3.349387, 3.344229, 3.379327, 3.366583, 
    3.400978, 3.391659, 3.406935, 3.399339, 3.398222, 3.388484, 3.38243, 
    3.367167, 3.35478, 3.344976, 3.347254, 3.358029, 3.377597, 3.396174, 
    3.392099, 3.405772, 3.369653, 3.38477, 3.378923, 3.394182, 3.360801, 
    3.389224, 3.353562, 3.356679, 3.36633, 3.3858, 3.390111, 3.394726, 
    3.391877, 3.378094, 3.375838, 3.366095, 3.363409, 3.356, 3.349875, 
    3.355472, 3.361356, 3.378098, 3.393234, 3.409784, 3.413841, 3.433266, 
    3.417453, 3.443578, 3.421366, 3.45987, 3.390871, 3.420707, 3.366769, 
    3.372552, 3.383034, 3.407143, 3.39411, 3.409354, 3.375749, 3.358403, 
    3.35392, 3.345572, 3.35411, 3.353415, 3.361598, 3.358967, 3.378655, 
    3.36807, 3.398195, 3.409232, 3.44052, 3.459792, 3.479474, 3.488188, 
    3.490842, 3.491953,
  2.997048, 3.013985, 3.010687, 3.024135, 3.016772, 3.025464, 3.000475, 
    3.01466, 3.005599, 2.998569, 3.049998, 3.024727, 3.076403, 3.060166, 
    3.101074, 3.073874, 3.106579, 3.100284, 3.119254, 3.113811, 3.138175, 
    3.121769, 3.150856, 3.134249, 3.136844, 3.121229, 3.029798, 3.046844, 
    3.02879, 3.031216, 3.030127, 3.016925, 3.010084, 2.995755, 2.998352, 
    3.008877, 3.032307, 3.02442, 3.044322, 3.043871, 3.066141, 3.056085, 
    3.093696, 3.082971, 3.114038, 3.106203, 3.11367, 3.111404, 3.113699, 
    3.102215, 3.107132, 3.09704, 3.057967, 3.069413, 3.035372, 3.014996, 
    3.001097, 2.991264, 2.992653, 2.995302, 3.008939, 3.021628, 3.03114, 
    3.037515, 3.043806, 3.062916, 3.07306, 3.09587, 3.091742, 3.098736, 
    3.105424, 3.116682, 3.114827, 3.119795, 3.098549, 3.112658, 3.089393, 
    3.095743, 3.045527, 3.026546, 3.018512, 3.011321, 2.993721, 3.005868, 
    3.001076, 3.012484, 3.019646, 3.016155, 3.03769, 3.029308, 3.073662, 
    3.054498, 3.104644, 3.092588, 3.107538, 3.099903, 3.112995, 3.10121, 
    3.121644, 3.126108, 3.123057, 3.134785, 3.100558, 3.113671, 3.016054, 
    3.016636, 3.019279, 3.007379, 3.006645, 2.995684, 3.005435, 3.009595, 
    3.020053, 3.026121, 3.031898, 3.044627, 3.058892, 3.078921, 3.093369, 
    3.103082, 3.097123, 3.102384, 3.096503, 3.09375, 3.124436, 3.107178, 
    3.133096, 3.131658, 3.119913, 3.13182, 3.017034, 3.013679, 3.001993, 
    3.011136, 2.994492, 3.003801, 3.009164, 3.029485, 3.03391, 3.038019, 
    3.046145, 3.056599, 3.075004, 3.091082, 3.105814, 3.104732, 3.105113, 
    3.108412, 3.100247, 3.109753, 3.111352, 3.107175, 3.131465, 3.124511, 
    3.131627, 3.127098, 3.014775, 3.020326, 3.017355, 3.022943, 3.019006, 
    3.036543, 3.041816, 3.066576, 3.056394, 3.072608, 3.058037, 3.060616, 
    3.073142, 3.058823, 3.090196, 3.068903, 3.10854, 3.087186, 3.109882, 
    3.10575, 3.112592, 3.118731, 3.126465, 3.140775, 3.137456, 3.14945, 
    3.028531, 3.035685, 3.035053, 3.042551, 3.048106, 3.060169, 3.079592, 
    3.072277, 3.085715, 3.088419, 3.068006, 3.080529, 3.040479, 3.046925, 
    3.043085, 3.029096, 3.073964, 3.050877, 3.093609, 3.081026, 3.117855, 
    3.0995, 3.135631, 3.151177, 3.165851, 3.183075, 3.039593, 3.034726, 
    3.043443, 3.055538, 3.066787, 3.081792, 3.08333, 3.086149, 3.093457, 
    3.099612, 3.087042, 3.101156, 3.048425, 3.075973, 3.032889, 3.045817, 
    3.054823, 3.050869, 3.071441, 3.076306, 3.096133, 3.085871, 3.147336, 
    3.120031, 3.19623, 3.174799, 3.033028, 3.039576, 3.06245, 3.05155, 
    3.082795, 3.090523, 3.096814, 3.104874, 3.105743, 3.110527, 3.102692, 
    3.110216, 3.081824, 3.094488, 3.059827, 3.068238, 3.064366, 3.060124, 
    3.073229, 3.08724, 3.087537, 3.09204, 3.104762, 3.082922, 3.150878, 
    3.108785, 3.046728, 3.059397, 3.061206, 3.056292, 3.089748, 3.077595, 
    3.110409, 3.101515, 3.116098, 3.108845, 3.107779, 3.098484, 3.092708, 
    3.078152, 3.066344, 3.057004, 3.059174, 3.069441, 3.088098, 3.105823, 
    3.101934, 3.114988, 3.080522, 3.094941, 3.089363, 3.103922, 3.072083, 
    3.099189, 3.065185, 3.068154, 3.077354, 3.095922, 3.100038, 3.104441, 
    3.101723, 3.088572, 3.08642, 3.077129, 3.074569, 3.067507, 3.061671, 
    3.067004, 3.072612, 3.088576, 3.103018, 3.118819, 3.122694, 3.141255, 
    3.126143, 3.151114, 3.12988, 3.166703, 3.100761, 3.129252, 3.077772, 
    3.083287, 3.093283, 3.116296, 3.103853, 3.118407, 3.086336, 3.069797, 
    3.065525, 3.057572, 3.065707, 3.065044, 3.072842, 3.070335, 3.089107, 
    3.079013, 3.107753, 3.118292, 3.148193, 3.16663, 3.185476, 3.193824, 
    3.196368, 3.197431,
  2.977271, 2.993924, 2.990679, 3.004162, 2.996675, 3.005514, 2.980639, 
    2.994588, 2.985676, 2.978765, 3.030494, 3.004765, 3.057168, 3.040863, 
    3.081575, 3.054667, 3.087028, 3.080793, 3.099591, 3.094194, 3.118366, 
    3.102085, 3.130966, 3.114469, 3.117045, 3.10155, 3.009924, 3.027281, 
    3.008899, 3.011368, 3.010259, 2.99683, 2.990086, 2.976, 2.978552, 
    2.988899, 3.012478, 3.004453, 3.024713, 3.024254, 3.046959, 3.036702, 
    3.074272, 3.063662, 3.094419, 3.086656, 3.094055, 3.091809, 3.094084, 
    3.082706, 3.087576, 3.077581, 3.038621, 3.05026, 3.015598, 2.994917, 
    2.98125, 2.971588, 2.972953, 2.975555, 2.98896, 3.001613, 3.01129, 
    3.017781, 3.024188, 3.043667, 3.053864, 3.076423, 3.072338, 3.07926, 
    3.085885, 3.097041, 3.095202, 3.100127, 3.079076, 3.093051, 3.070014, 
    3.076298, 3.025939, 3.006616, 2.998444, 2.991303, 2.974002, 2.98594, 
    2.981229, 2.992447, 2.999597, 2.996058, 3.017958, 3.009427, 3.054458, 
    3.035084, 3.085111, 3.073176, 3.087979, 3.080416, 3.093386, 3.081711, 
    3.101962, 3.106389, 3.103363, 3.115002, 3.081065, 3.094055, 2.99596, 
    2.996536, 2.999225, 2.987426, 2.986705, 2.97593, 2.985515, 2.989606, 
    3.000011, 3.006184, 3.012062, 3.025024, 3.039564, 3.059657, 3.073948, 
    3.083565, 3.077664, 3.082873, 3.077051, 3.074325, 3.10473, 3.087622, 
    3.113325, 3.111897, 3.100245, 3.112058, 2.996942, 2.993623, 2.982131, 
    2.991121, 2.974759, 2.983908, 2.989181, 3.009606, 3.01411, 3.018293, 
    3.026571, 3.037226, 3.055784, 3.071685, 3.08627, 3.085199, 3.085576, 
    3.088844, 3.080757, 3.090173, 3.091757, 3.087619, 3.111706, 3.104805, 
    3.111867, 3.107372, 2.994701, 3.000288, 2.997268, 3.00295, 2.998947, 
    3.01679, 3.022159, 3.047402, 3.037016, 3.053417, 3.038692, 3.041322, 
    3.053944, 3.039494, 3.070807, 3.049756, 3.088971, 3.06783, 3.090301, 
    3.086207, 3.092987, 3.099072, 3.106743, 3.120949, 3.117654, 3.129569, 
    3.008636, 3.015917, 3.015274, 3.022909, 3.028568, 3.040866, 3.060321, 
    3.05309, 3.066375, 3.06905, 3.048862, 3.061246, 3.020798, 3.027364, 
    3.023452, 3.00921, 3.054757, 3.031392, 3.074185, 3.061738, 3.098204, 
    3.080017, 3.115841, 3.131284, 3.145882, 3.163034, 3.019897, 3.014941, 
    3.023818, 3.036143, 3.047617, 3.062496, 3.064016, 3.066804, 3.074035, 
    3.080128, 3.067687, 3.081657, 3.028892, 3.056743, 3.013071, 3.026236, 
    3.035415, 3.031384, 3.052265, 3.057072, 3.076683, 3.066529, 3.127467, 
    3.100361, 3.176151, 3.154789, 3.013212, 3.019879, 3.043193, 3.032079, 
    3.063488, 3.071132, 3.077359, 3.085339, 3.0862, 3.09094, 3.083178, 
    3.090632, 3.062527, 3.075055, 3.040518, 3.049098, 3.045147, 3.040821, 
    3.054031, 3.067883, 3.068177, 3.072633, 3.085226, 3.063613, 3.130987, 
    3.089212, 3.027165, 3.040078, 3.041924, 3.036913, 3.070365, 3.058346, 
    3.090824, 3.082012, 3.096462, 3.089273, 3.088217, 3.079011, 3.073294, 
    3.058896, 3.047166, 3.037639, 3.039852, 3.050288, 3.068732, 3.08628, 
    3.082428, 3.095361, 3.061239, 3.075503, 3.069983, 3.084397, 3.052899, 
    3.079707, 3.045983, 3.049013, 3.058108, 3.076475, 3.080549, 3.08491, 
    3.082218, 3.069201, 3.067073, 3.057886, 3.055355, 3.048353, 3.042399, 
    3.047839, 3.053421, 3.069206, 3.0835, 3.099159, 3.103002, 3.121426, 
    3.106423, 3.131222, 3.11013, 3.146727, 3.081265, 3.109508, 3.058521, 
    3.063974, 3.073863, 3.096658, 3.084329, 3.098751, 3.066989, 3.050639, 
    3.04633, 3.038218, 3.046516, 3.04584, 3.053649, 3.051171, 3.069731, 
    3.059748, 3.088191, 3.098636, 3.128319, 3.146656, 3.165427, 3.173751, 
    3.176289, 3.17735,
  2.975963, 2.994363, 2.990775, 3.005696, 2.997407, 3.007194, 2.979681, 
    2.995097, 2.985244, 2.977613, 3.034918, 3.006363, 3.064926, 3.046454, 
    3.09312, 3.062044, 3.099434, 3.092216, 3.113999, 3.107739, 3.135817, 
    3.116894, 3.150495, 3.131283, 3.13428, 3.116272, 3.012081, 3.031345, 
    3.010945, 3.013681, 3.012453, 2.997578, 2.990118, 2.974561, 2.977378, 
    2.988806, 3.014913, 3.006018, 3.028493, 3.027983, 3.053245, 3.041823, 
    3.084674, 3.072418, 3.108, 3.099003, 3.107577, 3.104974, 3.107611, 
    3.094429, 3.100068, 3.0885, 3.043958, 3.056966, 3.018374, 2.995461, 
    2.980356, 2.969662, 2.971199, 2.97407, 2.988873, 3.002873, 3.013596, 
    3.020796, 3.02791, 3.049576, 3.061117, 3.08716, 3.082438, 3.090442, 
    3.09811, 3.11104, 3.108907, 3.114621, 3.090229, 3.106414, 3.079753, 
    3.087016, 3.029854, 3.008414, 2.999364, 2.991464, 2.972356, 2.985536, 
    2.980332, 2.992729, 3.000641, 2.996725, 3.020993, 3.011529, 3.061803, 
    3.040022, 3.097214, 3.083407, 3.100535, 3.091779, 3.106801, 3.093278, 
    3.11675, 3.121892, 3.118377, 3.131903, 3.09253, 3.107578, 2.996615, 
    2.997253, 3.000229, 2.987178, 2.986381, 2.974484, 2.985067, 2.989588, 
    3.0011, 3.007936, 3.014451, 3.028838, 3.045008, 3.067797, 3.084299, 
    3.095424, 3.088596, 3.094623, 3.087887, 3.084735, 3.119964, 3.100121, 
    3.129953, 3.128293, 3.114757, 3.128479, 2.997702, 2.99403, 2.981328, 
    2.991263, 2.973192, 2.983292, 2.989119, 3.011728, 3.016722, 3.021364, 
    3.030557, 3.042406, 3.063332, 3.081684, 3.098557, 3.097316, 3.097753, 
    3.101537, 3.092174, 3.103078, 3.104913, 3.100118, 3.12807, 3.120052, 
    3.128257, 3.123033, 2.995223, 3.001406, 2.998063, 3.004354, 2.999921, 
    3.019696, 3.025656, 3.053738, 3.042173, 3.060603, 3.044038, 3.046965, 
    3.061209, 3.04493, 3.08067, 3.056385, 3.101685, 3.077229, 3.103225, 
    3.098483, 3.106339, 3.113397, 3.122303, 3.138824, 3.134988, 3.148867, 
    3.010653, 3.018728, 3.018014, 3.026489, 3.032777, 3.046458, 3.068563, 
    3.060227, 3.075551, 3.078639, 3.055366, 3.069631, 3.024145, 3.031439, 
    3.027093, 3.01129, 3.062147, 3.035916, 3.084573, 3.070198, 3.112389, 
    3.091318, 3.132879, 3.150866, 3.167812, 3.187246, 3.023144, 3.017645, 
    3.027499, 3.041201, 3.053979, 3.071072, 3.072827, 3.076046, 3.0844, 
    3.091447, 3.077065, 3.093216, 3.033136, 3.064437, 3.01557, 3.030185, 
    3.04039, 3.035907, 3.059275, 3.064816, 3.087461, 3.075728, 3.146416, 
    3.114892, 3.202144, 3.177897, 3.015727, 3.023124, 3.049049, 3.03668, 
    3.072217, 3.081045, 3.088243, 3.097478, 3.098476, 3.103966, 3.094976, 
    3.103609, 3.071109, 3.08558, 3.04607, 3.055629, 3.051226, 3.046407, 
    3.061311, 3.077291, 3.077632, 3.082779, 3.097346, 3.072362, 3.150518, 
    3.101963, 3.031217, 3.04558, 3.047636, 3.042058, 3.080158, 3.066285, 
    3.103831, 3.093627, 3.110368, 3.102035, 3.100812, 3.090155, 3.083544, 
    3.06692, 3.053476, 3.042866, 3.045329, 3.056998, 3.078272, 3.098567, 
    3.094107, 3.109092, 3.069623, 3.086097, 3.079718, 3.096387, 3.060006, 
    3.090959, 3.052157, 3.055534, 3.06601, 3.08722, 3.091934, 3.096981, 
    3.093865, 3.078814, 3.076356, 3.065755, 3.062837, 3.054799, 3.048165, 
    3.054226, 3.060607, 3.07882, 3.095349, 3.113497, 3.117958, 3.139378, 
    3.12193, 3.150792, 3.126237, 3.168768, 3.092761, 3.125515, 3.066487, 
    3.072778, 3.0842, 3.110595, 3.096308, 3.113024, 3.076259, 3.057402, 
    3.052544, 3.04351, 3.052751, 3.051998, 3.060871, 3.058016, 3.079426, 
    3.067902, 3.100781, 3.112891, 3.147409, 3.168687, 3.189962, 3.199416, 
    3.202301, 3.203508,
  3.255175, 3.278651, 3.274064, 3.293171, 3.282547, 3.295094, 3.25991, 
    3.279591, 3.267002, 3.257275, 3.330354, 3.294028, 3.368128, 3.344837, 
    3.403923, 3.364486, 3.41198, 3.402771, 3.430626, 3.422602, 3.458712, 
    3.434342, 3.477714, 3.452861, 3.456727, 3.433544, 3.301373, 3.325879, 
    3.299912, 3.30343, 3.30185, 3.282766, 3.273225, 3.253391, 3.256976, 
    3.271549, 3.305014, 3.293585, 3.32231, 3.321672, 3.353385, 3.339017, 
    3.393168, 3.377611, 3.422936, 3.41143, 3.422395, 3.419063, 3.422438, 
    3.405593, 3.412791, 3.398038, 3.3417, 3.358076, 3.309469, 3.280057, 
    3.260769, 3.247204, 3.249116, 3.252766, 3.271635, 3.28955, 3.30332, 
    3.312589, 3.32158, 3.348765, 3.363315, 3.396332, 3.390326, 3.40051, 
    3.41029, 3.426831, 3.424098, 3.431424, 3.400239, 3.420905, 3.386915, 
    3.396148, 3.324013, 3.296661, 3.285053, 3.274945, 3.250587, 3.267375, 
    3.260739, 3.276563, 3.286689, 3.281673, 3.312843, 3.300663, 3.364182, 
    3.336756, 3.409146, 3.391557, 3.413387, 3.402214, 3.421402, 3.404124, 
    3.434157, 3.440765, 3.436247, 3.45366, 3.403171, 3.422395, 3.281533, 
    3.282351, 3.286161, 3.26947, 3.268453, 3.253294, 3.266776, 3.272547, 
    3.287277, 3.296046, 3.304421, 3.322742, 3.343019, 3.371759, 3.392692, 
    3.406861, 3.398159, 3.40584, 3.397256, 3.393247, 3.438287, 3.412859, 
    3.451145, 3.449005, 3.431599, 3.449246, 3.282924, 3.278226, 3.262009, 
    3.274688, 3.25165, 3.264512, 3.271948, 3.300919, 3.307343, 3.313323, 
    3.324893, 3.33975, 3.366113, 3.389368, 3.41086, 3.409276, 3.409833, 
    3.414668, 3.402717, 3.416637, 3.418985, 3.412855, 3.448719, 3.4384, 
    3.44896, 3.442233, 3.279752, 3.28767, 3.283387, 3.29145, 3.285767, 
    3.311172, 3.318763, 3.354007, 3.339457, 3.362666, 3.3418, 3.34548, 
    3.363432, 3.342921, 3.388079, 3.357343, 3.414856, 3.383712, 3.416826, 
    3.410766, 3.42081, 3.429853, 3.441294, 3.462598, 3.457642, 3.475602, 
    3.299537, 3.309925, 3.309006, 3.319804, 3.327672, 3.344842, 3.372729, 
    3.362191, 3.381582, 3.385501, 3.356058, 3.37408, 3.316874, 3.325996, 
    3.320558, 3.300355, 3.364616, 3.331606, 3.39304, 3.374799, 3.428561, 
    3.401626, 3.45492, 3.478196, 3.500371, 3.526644, 3.315617, 3.308531, 
    3.321067, 3.338236, 3.35431, 3.375906, 3.378129, 3.38221, 3.39282, 
    3.40179, 3.383503, 3.404046, 3.328121, 3.36751, 3.30586, 3.324426, 
    3.337219, 3.331594, 3.36099, 3.36799, 3.396715, 3.381808, 3.472425, 
    3.431772, 3.54653, 3.513984, 3.306062, 3.315592, 3.348101, 3.332563, 
    3.377356, 3.388556, 3.39771, 3.409482, 3.410757, 3.417773, 3.40629, 
    3.417317, 3.375952, 3.39432, 3.344355, 3.35639, 3.350843, 3.344779, 
    3.36356, 3.38379, 3.384223, 3.39076, 3.409314, 3.37754, 3.477744, 
    3.415212, 3.325719, 3.343738, 3.346324, 3.339313, 3.38743, 3.369847, 
    3.417601, 3.404569, 3.425971, 3.415304, 3.413741, 3.400144, 3.391732, 
    3.37065, 3.353676, 3.340328, 3.343422, 3.358116, 3.385035, 3.410873, 
    3.405182, 3.424335, 3.374071, 3.394979, 3.38687, 3.40809, 3.361912, 
    3.401168, 3.352015, 3.356271, 3.369499, 3.396408, 3.402411, 3.408849, 
    3.404873, 3.385723, 3.382603, 3.369176, 3.365488, 3.355343, 3.346989, 
    3.354621, 3.362672, 3.38573, 3.406766, 3.429983, 3.435709, 3.463314, 
    3.440814, 3.478099, 3.446357, 3.501659, 3.403466, 3.445426, 3.370103, 
    3.378067, 3.392566, 3.426261, 3.40799, 3.429375, 3.382481, 3.358626, 
    3.352502, 3.341137, 3.352763, 3.351814, 3.363004, 3.359401, 3.3865, 
    3.371893, 3.413702, 3.429204, 3.473712, 3.50155, 3.53033, 3.542928, 
    3.546737, 3.548332,
  3.812404, 3.852935, 3.844963, 3.878335, 3.859724, 3.881718, 3.820526, 
    3.85457, 3.832741, 3.816003, 3.945439, 3.879842, 4.016918, 3.9726, 
    4.084901, 4.009933, 4.100402, 4.082692, 4.136672, 4.120995, 4.192386, 
    4.143967, 4.230846, 4.180668, 4.188405, 4.142399, 3.892797, 3.937107, 
    3.890216, 3.896439, 3.893642, 3.860107, 3.843508, 3.809351, 3.81549, 
    3.840605, 3.899246, 3.879063, 3.930481, 3.929299, 3.988772, 3.961649, 
    4.064366, 4.034974, 4.121646, 4.09934, 4.120591, 4.114113, 4.120676, 
    4.088104, 4.101967, 4.073641, 3.966691, 3.997692, 3.907158, 3.855382, 
    3.822003, 3.79879, 3.802049, 3.808282, 3.840753, 3.871976, 3.896244, 
    3.912714, 3.929129, 3.980018, 4.007694, 4.070388, 4.058969, 4.078364, 
    4.097141, 4.129246, 4.12391, 4.138237, 4.077846, 4.117693, 4.052508, 
    4.070038, 3.93364, 3.884479, 3.864102, 3.846492, 3.804559, 3.833384, 
    3.821951, 3.849302, 3.866964, 3.8582, 3.913167, 3.891543, 4.009351, 
    3.957408, 4.094938, 4.061305, 4.103119, 4.081626, 4.118659, 4.085286, 
    4.143604, 4.156631, 4.147717, 4.182266, 4.083459, 4.120593, 3.857956, 
    3.859382, 3.86604, 3.837005, 3.835248, 3.809184, 3.83235, 3.842334, 
    3.867993, 3.883395, 3.898193, 3.931283, 3.969174, 4.0239, 4.063461, 
    4.090542, 4.073873, 4.088579, 4.07215, 4.064516, 4.151737, 4.102098, 
    4.177245, 4.17298, 4.13858, 4.17346, 3.860383, 3.852195, 3.824135, 
    3.846047, 3.806375, 3.828445, 3.841295, 3.891995, 3.903378, 3.914021, 
    3.935274, 3.963025, 4.013051, 4.057152, 4.09824, 4.095188, 4.096262, 
    4.105596, 4.08259, 4.109409, 4.113963, 4.102091, 4.17241, 4.15196, 
    4.172889, 4.159536, 3.854851, 3.868681, 3.861192, 3.87531, 3.86535, 
    3.910189, 3.923914, 3.989952, 3.962475, 4.006453, 3.966879, 3.973813, 
    4.007917, 3.968989, 4.054711, 3.996297, 4.10596, 4.046457, 4.109775, 
    4.09806, 4.117507, 4.135158, 4.157678, 4.200199, 4.190238, 4.22654, 
    3.889553, 3.907968, 3.906334, 3.925841, 3.940442, 3.972609, 4.025767, 
    4.005544, 4.042443, 4.049835, 3.993851, 4.028355, 3.920425, 3.937325, 
    3.927237, 3.890998, 4.010183, 3.947774, 4.064123, 4.0297, 4.132628, 
    4.080499, 4.184785, 4.23183, 4.277549, 4.332258, 3.918117, 3.905489, 
    3.928178, 3.960184, 3.990528, 4.031776, 4.035948, 4.043625, 4.063704, 
    4.080814, 4.046064, 4.085135, 3.941279, 4.01573, 3.900746, 3.934408, 
    3.958276, 3.947753, 4.00325, 4.016651, 4.071118, 4.042867, 4.220077, 
    4.138919, 4.374618, 4.306069, 3.901104, 3.918072, 3.978763, 3.949563, 
    4.034496, 4.055614, 4.073015, 4.095585, 4.098041, 4.11161, 4.089443, 
    4.110727, 4.031862, 4.066557, 3.97169, 3.994482, 3.983951, 3.972489, 
    4.008162, 4.046605, 4.047421, 4.059792, 4.095261, 4.034841, 4.230908, 
    4.106648, 3.93681, 3.970529, 3.975405, 3.962204, 4.053482, 4.020219, 
    4.111277, 4.08614, 4.127563, 4.106827, 4.103803, 4.077665, 4.061636, 
    4.021764, 3.989324, 3.96411, 3.969933, 3.997768, 4.048954, 4.098266, 
    4.087316, 4.124372, 4.028337, 4.067811, 4.052423, 4.092905, 4.005012, 
    4.079624, 3.986172, 3.994256, 4.019552, 4.070532, 4.082003, 4.094365, 
    4.086723, 4.050254, 4.044367, 4.01893, 4.011853, 3.992491, 3.97666, 
    3.991119, 4.006463, 4.050267, 4.090358, 4.135411, 4.146657, 4.201643, 
    4.15673, 4.231632, 4.167714, 4.280233, 4.084023, 4.165866, 4.020712, 
    4.035832, 4.063222, 4.128131, 4.092711, 4.134221, 4.044136, 3.998741, 
    3.987096, 3.965631, 3.987591, 3.985792, 4.007099, 4.000217, 4.051724, 
    4.024157, 4.103728, 4.133887, 4.222694, 4.280007, 4.339907, 4.366786, 
    4.375068, 4.378545,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 6.889972, 
    6.889972, 6.889972,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HC =
  24856.02, 24876.84, 24872.76, 24889.8, 24880.32, 24891.52, 24860.21, 
    24877.68, 24866.49, 24857.88, 24923.61, 24890.56, 24958.98, 24937.12, 
    24992.49, 24955.55, 25000.08, 24991.4, 25017.75, 25010.13, 25044.64, 
    25021.29, 25063.04, 25039.01, 25042.73, 25020.53, 24897.14, 24919.45, 
    24895.83, 24898.99, 24897.57, 24880.51, 24872.02, 24854.44, 24857.61, 
    24870.53, 24900.41, 24890.17, 24916.14, 24915.55, 24945.12, 24931.68, 
    24982.4, 24967.88, 25010.44, 24999.56, 25009.93, 25006.77, 25009.97, 
    24994.06, 25000.84, 24986.96, 24934.18, 24949.53, 24904.41, 24878.1, 
    24860.97, 24848.98, 24850.67, 24853.89, 24870.6, 24886.56, 24898.89, 
    24907.22, 24915.46, 24940.79, 24954.45, 24985.36, 24979.74, 24989.28, 
    24998.48, 25014.14, 25011.54, 25018.51, 24989.03, 25008.52, 24976.55, 
    24985.19, 24917.72, 24892.92, 24882.55, 24873.54, 24851.97, 24866.82, 
    24860.94, 24874.98, 24884.01, 24879.54, 24907.45, 24896.51, 24955.27, 
    24929.57, 24997.41, 24980.89, 25001.41, 24990.88, 25008.99, 24992.68, 
    25021.11, 25027.42, 25023.1, 25039.78, 24991.78, 25009.93, 24879.41, 
    24880.14, 24883.54, 24868.68, 24867.78, 24854.36, 24866.29, 24871.41, 
    24884.53, 24892.37, 24899.88, 24916.54, 24935.42, 24962.41, 24981.95, 
    24995.25, 24987.07, 24994.29, 24986.23, 24982.47, 25025.05, 25000.91, 
    25037.36, 25035.31, 25018.67, 25035.54, 24880.65, 24876.47, 24862.06, 
    24873.32, 24852.9, 24864.28, 24870.88, 24896.73, 24902.5, 24907.88, 
    24918.54, 24932.36, 24957.08, 24978.84, 24999.02, 24997.53, 24998.05, 
    25002.62, 24991.35, 25004.48, 25006.7, 25000.9, 25035.03, 25025.16, 
    25035.26, 25028.82, 24877.82, 24884.88, 24881.06, 24888.26, 24883.19, 
    24905.94, 24912.85, 24945.71, 24932.09, 24953.84, 24934.28, 24937.72, 
    24954.56, 24935.32, 24977.64, 24948.84, 25002.79, 24973.56, 25004.66, 
    24998.93, 25008.43, 25017.01, 25027.92, 25048.39, 25043.61, 25060.98, 
    24895.5, 24904.82, 24904, 24913.82, 24921.12, 24937.12, 24963.32, 
    24953.39, 24971.57, 24975.23, 24947.63, 24964.59, 24911.1, 24919.56, 
    24914.52, 24896.23, 24955.68, 24924.77, 24982.28, 24965.26, 25015.79, 
    24990.33, 25040.99, 25063.51, 25085.18, 25110.93, 24909.95, 24903.57, 
    24914.99, 24930.95, 24945.99, 24966.29, 24968.36, 24972.16, 24982.07, 
    24990.48, 24973.37, 24992.6, 24921.53, 24958.4, 24901.17, 24918.1, 24930, 
    24924.76, 24952.26, 24958.85, 24985.72, 24971.78, 25057.9, 25018.84, 
    25130.76, 25098.57, 24901.35, 24909.92, 24940.17, 24925.66, 24967.64, 
    24978.08, 24986.65, 24997.72, 24998.92, 25005.55, 24994.71, 25005.12, 
    24966.33, 24983.47, 24936.66, 24947.95, 24942.74, 24937.06, 24954.68, 
    24973.63, 24974.04, 24980.14, 24997.56, 24967.81, 25063.07, 25003.13, 
    24919.3, 24936.09, 24938.51, 24931.96, 24977.03, 24960.6, 25005.39, 
    24993.1, 25013.32, 25003.22, 25001.74, 24988.94, 24981.05, 24961.36, 
    24945.4, 24932.9, 24935.79, 24949.56, 24974.79, 24999.04, 24993.67, 
    25011.77, 24964.59, 24984.09, 24976.51, 24996.41, 24953.13, 24989.9, 
    24943.84, 24947.83, 24960.28, 24985.43, 24991.07, 24997.12, 24993.38, 
    24975.44, 24972.53, 24959.97, 24956.5, 24946.96, 24939.13, 24946.28, 
    24953.85, 24975.44, 24995.16, 25017.14, 25022.59, 25049.08, 25027.46, 
    25063.41, 25032.77, 25086.44, 24992.06, 25031.88, 24960.84, 24968.3, 
    24981.83, 25013.6, 24996.32, 25016.56, 24972.41, 24950.04, 24944.29, 
    24933.66, 24944.54, 24943.65, 24954.16, 24950.77, 24976.16, 24962.53, 
    25001.71, 25016.4, 25059.15, 25086.33, 25114.53, 25127.11, 25130.97, 
    25132.58 ;

 HCSOI =
  24856.02, 24876.84, 24872.76, 24889.8, 24880.32, 24891.52, 24860.21, 
    24877.68, 24866.49, 24857.88, 24923.61, 24890.56, 24958.98, 24937.12, 
    24992.49, 24955.55, 25000.08, 24991.4, 25017.75, 25010.13, 25044.64, 
    25021.29, 25063.04, 25039.01, 25042.73, 25020.53, 24897.14, 24919.45, 
    24895.83, 24898.99, 24897.57, 24880.51, 24872.02, 24854.44, 24857.61, 
    24870.53, 24900.41, 24890.17, 24916.14, 24915.55, 24945.12, 24931.68, 
    24982.4, 24967.88, 25010.44, 24999.56, 25009.93, 25006.77, 25009.97, 
    24994.06, 25000.84, 24986.96, 24934.18, 24949.53, 24904.41, 24878.1, 
    24860.97, 24848.98, 24850.67, 24853.89, 24870.6, 24886.56, 24898.89, 
    24907.22, 24915.46, 24940.79, 24954.45, 24985.36, 24979.74, 24989.28, 
    24998.48, 25014.14, 25011.54, 25018.51, 24989.03, 25008.52, 24976.55, 
    24985.19, 24917.72, 24892.92, 24882.55, 24873.54, 24851.97, 24866.82, 
    24860.94, 24874.98, 24884.01, 24879.54, 24907.45, 24896.51, 24955.27, 
    24929.57, 24997.41, 24980.89, 25001.41, 24990.88, 25008.99, 24992.68, 
    25021.11, 25027.42, 25023.1, 25039.78, 24991.78, 25009.93, 24879.41, 
    24880.14, 24883.54, 24868.68, 24867.78, 24854.36, 24866.29, 24871.41, 
    24884.53, 24892.37, 24899.88, 24916.54, 24935.42, 24962.41, 24981.95, 
    24995.25, 24987.07, 24994.29, 24986.23, 24982.47, 25025.05, 25000.91, 
    25037.36, 25035.31, 25018.67, 25035.54, 24880.65, 24876.47, 24862.06, 
    24873.32, 24852.9, 24864.28, 24870.88, 24896.73, 24902.5, 24907.88, 
    24918.54, 24932.36, 24957.08, 24978.84, 24999.02, 24997.53, 24998.05, 
    25002.62, 24991.35, 25004.48, 25006.7, 25000.9, 25035.03, 25025.16, 
    25035.26, 25028.82, 24877.82, 24884.88, 24881.06, 24888.26, 24883.19, 
    24905.94, 24912.85, 24945.71, 24932.09, 24953.84, 24934.28, 24937.72, 
    24954.56, 24935.32, 24977.64, 24948.84, 25002.79, 24973.56, 25004.66, 
    24998.93, 25008.43, 25017.01, 25027.92, 25048.39, 25043.61, 25060.98, 
    24895.5, 24904.82, 24904, 24913.82, 24921.12, 24937.12, 24963.32, 
    24953.39, 24971.57, 24975.23, 24947.63, 24964.59, 24911.1, 24919.56, 
    24914.52, 24896.23, 24955.68, 24924.77, 24982.28, 24965.26, 25015.79, 
    24990.33, 25040.99, 25063.51, 25085.18, 25110.93, 24909.95, 24903.57, 
    24914.99, 24930.95, 24945.99, 24966.29, 24968.36, 24972.16, 24982.07, 
    24990.48, 24973.37, 24992.6, 24921.53, 24958.4, 24901.17, 24918.1, 24930, 
    24924.76, 24952.26, 24958.85, 24985.72, 24971.78, 25057.9, 25018.84, 
    25130.76, 25098.57, 24901.35, 24909.92, 24940.17, 24925.66, 24967.64, 
    24978.08, 24986.65, 24997.72, 24998.92, 25005.55, 24994.71, 25005.12, 
    24966.33, 24983.47, 24936.66, 24947.95, 24942.74, 24937.06, 24954.68, 
    24973.63, 24974.04, 24980.14, 24997.56, 24967.81, 25063.07, 25003.13, 
    24919.3, 24936.09, 24938.51, 24931.96, 24977.03, 24960.6, 25005.39, 
    24993.1, 25013.32, 25003.22, 25001.74, 24988.94, 24981.05, 24961.36, 
    24945.4, 24932.9, 24935.79, 24949.56, 24974.79, 24999.04, 24993.67, 
    25011.77, 24964.59, 24984.09, 24976.51, 24996.41, 24953.13, 24989.9, 
    24943.84, 24947.83, 24960.28, 24985.43, 24991.07, 24997.12, 24993.38, 
    24975.44, 24972.53, 24959.97, 24956.5, 24946.96, 24939.13, 24946.28, 
    24953.85, 24975.44, 24995.16, 25017.14, 25022.59, 25049.08, 25027.46, 
    25063.41, 25032.77, 25086.44, 24992.06, 25031.88, 24960.84, 24968.3, 
    24981.83, 25013.6, 24996.32, 25016.56, 24972.41, 24950.04, 24944.29, 
    24933.66, 24944.54, 24943.65, 24954.16, 24950.77, 24976.16, 24962.53, 
    25001.71, 25016.4, 25059.15, 25086.33, 25114.53, 25127.11, 25130.97, 
    25132.58 ;

 HEAT_FROM_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HR =
  6.191209e-08, 6.218511e-08, 6.213204e-08, 6.235225e-08, 6.22301e-08, 
    6.237429e-08, 6.196745e-08, 6.219594e-08, 6.205008e-08, 6.193667e-08, 
    6.277961e-08, 6.236208e-08, 6.321343e-08, 6.29471e-08, 6.361618e-08, 
    6.317198e-08, 6.370576e-08, 6.360339e-08, 6.391155e-08, 6.382326e-08, 
    6.421742e-08, 6.39523e-08, 6.442178e-08, 6.415411e-08, 6.419598e-08, 
    6.394355e-08, 6.244612e-08, 6.272763e-08, 6.242944e-08, 6.246958e-08, 
    6.245157e-08, 6.223262e-08, 6.212228e-08, 6.189123e-08, 6.193318e-08, 
    6.210288e-08, 6.248763e-08, 6.235703e-08, 6.26862e-08, 6.267877e-08, 
    6.304526e-08, 6.288002e-08, 6.349605e-08, 6.332096e-08, 6.382695e-08, 
    6.369969e-08, 6.382097e-08, 6.37842e-08, 6.382145e-08, 6.363481e-08, 
    6.371478e-08, 6.355055e-08, 6.291096e-08, 6.309892e-08, 6.253835e-08, 
    6.220129e-08, 6.197747e-08, 6.181863e-08, 6.184109e-08, 6.188389e-08, 
    6.210387e-08, 6.231072e-08, 6.246836e-08, 6.25738e-08, 6.267771e-08, 
    6.299219e-08, 6.315867e-08, 6.353144e-08, 6.346419e-08, 6.357814e-08, 
    6.368703e-08, 6.386984e-08, 6.383975e-08, 6.392029e-08, 6.357515e-08, 
    6.380452e-08, 6.342587e-08, 6.352943e-08, 6.27059e-08, 6.239227e-08, 
    6.225892e-08, 6.214224e-08, 6.185834e-08, 6.205439e-08, 6.19771e-08, 
    6.216099e-08, 6.227782e-08, 6.222004e-08, 6.257669e-08, 6.243803e-08, 
    6.316854e-08, 6.285387e-08, 6.367434e-08, 6.347799e-08, 6.372139e-08, 
    6.359719e-08, 6.381001e-08, 6.361848e-08, 6.395027e-08, 6.402251e-08, 
    6.397314e-08, 6.41628e-08, 6.360786e-08, 6.382096e-08, 6.221842e-08, 
    6.222784e-08, 6.227175e-08, 6.207874e-08, 6.206693e-08, 6.189008e-08, 
    6.204745e-08, 6.211446e-08, 6.22846e-08, 6.238523e-08, 6.248089e-08, 
    6.269123e-08, 6.292615e-08, 6.325467e-08, 6.349072e-08, 6.364895e-08, 
    6.355192e-08, 6.363758e-08, 6.354183e-08, 6.349695e-08, 6.399544e-08, 
    6.371552e-08, 6.413553e-08, 6.411229e-08, 6.39222e-08, 6.411491e-08, 
    6.223446e-08, 6.218023e-08, 6.199193e-08, 6.213929e-08, 6.187082e-08, 
    6.202109e-08, 6.210749e-08, 6.244091e-08, 6.251418e-08, 6.258211e-08, 
    6.271628e-08, 6.288847e-08, 6.319055e-08, 6.34534e-08, 6.369337e-08, 
    6.367579e-08, 6.368198e-08, 6.373558e-08, 6.36028e-08, 6.375738e-08, 
    6.378333e-08, 6.371549e-08, 6.410917e-08, 6.39967e-08, 6.411179e-08, 
    6.403856e-08, 6.219786e-08, 6.228911e-08, 6.22398e-08, 6.233252e-08, 
    6.22672e-08, 6.255767e-08, 6.264477e-08, 6.305234e-08, 6.288508e-08, 
    6.315129e-08, 6.291213e-08, 6.29545e-08, 6.315996e-08, 6.292505e-08, 
    6.34389e-08, 6.30905e-08, 6.373767e-08, 6.338972e-08, 6.375947e-08, 
    6.369233e-08, 6.38035e-08, 6.390305e-08, 6.402831e-08, 6.425942e-08, 
    6.420591e-08, 6.43992e-08, 6.242516e-08, 6.254352e-08, 6.25331e-08, 
    6.265698e-08, 6.27486e-08, 6.294718e-08, 6.326568e-08, 6.314591e-08, 
    6.33658e-08, 6.340995e-08, 6.307588e-08, 6.328098e-08, 6.262274e-08, 
    6.272907e-08, 6.266577e-08, 6.243449e-08, 6.317349e-08, 6.279422e-08, 
    6.349462e-08, 6.328914e-08, 6.388886e-08, 6.359058e-08, 6.417645e-08, 
    6.442689e-08, 6.466265e-08, 6.493813e-08, 6.260812e-08, 6.25277e-08, 
    6.267172e-08, 6.287096e-08, 6.305586e-08, 6.330166e-08, 6.332682e-08, 
    6.337287e-08, 6.349217e-08, 6.359246e-08, 6.338743e-08, 6.361761e-08, 
    6.275372e-08, 6.320642e-08, 6.249729e-08, 6.27108e-08, 6.285921e-08, 
    6.279412e-08, 6.313223e-08, 6.321191e-08, 6.353574e-08, 6.336835e-08, 
    6.436507e-08, 6.392407e-08, 6.514793e-08, 6.480587e-08, 6.249959e-08, 
    6.260785e-08, 6.298463e-08, 6.280536e-08, 6.331808e-08, 6.344429e-08, 
    6.35469e-08, 6.367805e-08, 6.369222e-08, 6.376993e-08, 6.364259e-08, 
    6.376491e-08, 6.330219e-08, 6.350896e-08, 6.294157e-08, 6.307966e-08, 
    6.301614e-08, 6.294646e-08, 6.316152e-08, 6.339064e-08, 6.339556e-08, 
    6.346902e-08, 6.367603e-08, 6.332016e-08, 6.442196e-08, 6.374147e-08, 
    6.27259e-08, 6.293441e-08, 6.296421e-08, 6.288344e-08, 6.343164e-08, 
    6.3233e-08, 6.376804e-08, 6.362344e-08, 6.386038e-08, 6.374263e-08, 
    6.372531e-08, 6.357409e-08, 6.347994e-08, 6.32421e-08, 6.304859e-08, 
    6.289515e-08, 6.293084e-08, 6.309938e-08, 6.340467e-08, 6.36935e-08, 
    6.363022e-08, 6.384236e-08, 6.32809e-08, 6.351632e-08, 6.342533e-08, 
    6.36626e-08, 6.314273e-08, 6.358538e-08, 6.302958e-08, 6.307831e-08, 
    6.322905e-08, 6.353228e-08, 6.359939e-08, 6.367102e-08, 6.362682e-08, 
    6.341242e-08, 6.33773e-08, 6.322539e-08, 6.318344e-08, 6.30677e-08, 
    6.297188e-08, 6.305942e-08, 6.315137e-08, 6.341251e-08, 6.364786e-08, 
    6.390447e-08, 6.396727e-08, 6.426707e-08, 6.4023e-08, 6.442575e-08, 
    6.40833e-08, 6.467612e-08, 6.361105e-08, 6.407326e-08, 6.323592e-08, 
    6.332613e-08, 6.348927e-08, 6.386351e-08, 6.366148e-08, 6.389776e-08, 
    6.337593e-08, 6.310519e-08, 6.303516e-08, 6.290448e-08, 6.303815e-08, 
    6.302728e-08, 6.315518e-08, 6.311409e-08, 6.342119e-08, 6.325622e-08, 
    6.372487e-08, 6.38959e-08, 6.437893e-08, 6.467506e-08, 6.497654e-08, 
    6.510964e-08, 6.515015e-08, 6.516709e-08 ;

 HR_vr =
  2.673865e-07, 2.681188e-07, 2.679765e-07, 2.685667e-07, 2.682395e-07, 
    2.686258e-07, 2.675351e-07, 2.681477e-07, 2.677568e-07, 2.674526e-07, 
    2.697106e-07, 2.685931e-07, 2.708713e-07, 2.701594e-07, 2.719471e-07, 
    2.707604e-07, 2.721862e-07, 2.719132e-07, 2.727355e-07, 2.725e-07, 
    2.735503e-07, 2.728441e-07, 2.740947e-07, 2.733819e-07, 2.734933e-07, 
    2.728208e-07, 2.688184e-07, 2.695715e-07, 2.687736e-07, 2.688811e-07, 
    2.688329e-07, 2.682461e-07, 2.679501e-07, 2.673307e-07, 2.674432e-07, 
    2.678983e-07, 2.689294e-07, 2.685797e-07, 2.694614e-07, 2.694415e-07, 
    2.70422e-07, 2.6998e-07, 2.716266e-07, 2.71159e-07, 2.725099e-07, 
    2.721703e-07, 2.724938e-07, 2.723958e-07, 2.724951e-07, 2.719971e-07, 
    2.722105e-07, 2.717722e-07, 2.700627e-07, 2.705654e-07, 2.690653e-07, 
    2.681618e-07, 2.675619e-07, 2.671358e-07, 2.671961e-07, 2.673109e-07, 
    2.679009e-07, 2.684556e-07, 2.68878e-07, 2.691604e-07, 2.694386e-07, 
    2.702795e-07, 2.707249e-07, 2.71721e-07, 2.715416e-07, 2.718457e-07, 
    2.721365e-07, 2.726242e-07, 2.72544e-07, 2.727587e-07, 2.718378e-07, 
    2.724499e-07, 2.714393e-07, 2.717158e-07, 2.695133e-07, 2.686741e-07, 
    2.683163e-07, 2.680038e-07, 2.672424e-07, 2.677682e-07, 2.675609e-07, 
    2.680542e-07, 2.683674e-07, 2.682126e-07, 2.691681e-07, 2.687967e-07, 
    2.707513e-07, 2.699099e-07, 2.721026e-07, 2.715784e-07, 2.722282e-07, 
    2.718967e-07, 2.724645e-07, 2.719536e-07, 2.728387e-07, 2.730312e-07, 
    2.728996e-07, 2.734052e-07, 2.719252e-07, 2.724938e-07, 2.682082e-07, 
    2.682334e-07, 2.683512e-07, 2.678335e-07, 2.678019e-07, 2.673276e-07, 
    2.677497e-07, 2.679294e-07, 2.683856e-07, 2.686552e-07, 2.689115e-07, 
    2.694748e-07, 2.701032e-07, 2.709817e-07, 2.716124e-07, 2.720349e-07, 
    2.717759e-07, 2.720045e-07, 2.717489e-07, 2.716291e-07, 2.72959e-07, 
    2.722124e-07, 2.733325e-07, 2.732706e-07, 2.727637e-07, 2.732776e-07, 
    2.682512e-07, 2.681058e-07, 2.676008e-07, 2.679961e-07, 2.672759e-07, 
    2.67679e-07, 2.679106e-07, 2.688043e-07, 2.690007e-07, 2.691826e-07, 
    2.695419e-07, 2.700026e-07, 2.708103e-07, 2.715126e-07, 2.721534e-07, 
    2.721065e-07, 2.72123e-07, 2.72266e-07, 2.719117e-07, 2.723242e-07, 
    2.723933e-07, 2.722124e-07, 2.732623e-07, 2.729625e-07, 2.732693e-07, 
    2.730741e-07, 2.681531e-07, 2.683977e-07, 2.682655e-07, 2.68514e-07, 
    2.683389e-07, 2.69117e-07, 2.693501e-07, 2.704407e-07, 2.699935e-07, 
    2.707054e-07, 2.700659e-07, 2.701792e-07, 2.707282e-07, 2.701005e-07, 
    2.714737e-07, 2.705426e-07, 2.722716e-07, 2.713422e-07, 2.723298e-07, 
    2.721507e-07, 2.724473e-07, 2.727127e-07, 2.730468e-07, 2.736624e-07, 
    2.7352e-07, 2.740347e-07, 2.687622e-07, 2.690792e-07, 2.690514e-07, 
    2.693831e-07, 2.696283e-07, 2.701597e-07, 2.710112e-07, 2.706911e-07, 
    2.712788e-07, 2.713967e-07, 2.70504e-07, 2.71052e-07, 2.692913e-07, 
    2.695758e-07, 2.694066e-07, 2.687871e-07, 2.707647e-07, 2.697502e-07, 
    2.716228e-07, 2.710739e-07, 2.726749e-07, 2.718789e-07, 2.734415e-07, 
    2.741081e-07, 2.747359e-07, 2.754679e-07, 2.692523e-07, 2.690369e-07, 
    2.694226e-07, 2.699556e-07, 2.704503e-07, 2.711074e-07, 2.711747e-07, 
    2.712976e-07, 2.716163e-07, 2.718841e-07, 2.713363e-07, 2.719512e-07, 
    2.696414e-07, 2.708528e-07, 2.689554e-07, 2.695269e-07, 2.699242e-07, 
    2.697501e-07, 2.706546e-07, 2.708676e-07, 2.717325e-07, 2.712856e-07, 
    2.739434e-07, 2.727685e-07, 2.760254e-07, 2.751165e-07, 2.689617e-07, 
    2.692516e-07, 2.702597e-07, 2.697802e-07, 2.711513e-07, 2.714884e-07, 
    2.717625e-07, 2.721124e-07, 2.721503e-07, 2.723577e-07, 2.720179e-07, 
    2.723443e-07, 2.711087e-07, 2.716612e-07, 2.701448e-07, 2.70514e-07, 
    2.703442e-07, 2.701578e-07, 2.707329e-07, 2.713449e-07, 2.713583e-07, 
    2.715544e-07, 2.721062e-07, 2.711569e-07, 2.740944e-07, 2.722809e-07, 
    2.695676e-07, 2.701253e-07, 2.702052e-07, 2.699892e-07, 2.714546e-07, 
    2.709239e-07, 2.723527e-07, 2.719668e-07, 2.72599e-07, 2.722849e-07, 
    2.722386e-07, 2.718351e-07, 2.715836e-07, 2.709482e-07, 2.704309e-07, 
    2.700206e-07, 2.70116e-07, 2.705667e-07, 2.713824e-07, 2.721536e-07, 
    2.719847e-07, 2.72551e-07, 2.71052e-07, 2.716807e-07, 2.714376e-07, 
    2.720713e-07, 2.706826e-07, 2.718644e-07, 2.703802e-07, 2.705104e-07, 
    2.709133e-07, 2.717231e-07, 2.719026e-07, 2.720937e-07, 2.719758e-07, 
    2.714032e-07, 2.713094e-07, 2.709036e-07, 2.707914e-07, 2.704821e-07, 
    2.702258e-07, 2.704599e-07, 2.707056e-07, 2.714035e-07, 2.720319e-07, 
    2.727165e-07, 2.728841e-07, 2.736824e-07, 2.730322e-07, 2.741044e-07, 
    2.731923e-07, 2.74771e-07, 2.719332e-07, 2.73166e-07, 2.709318e-07, 
    2.711728e-07, 2.716083e-07, 2.72607e-07, 2.720683e-07, 2.726984e-07, 
    2.713058e-07, 2.70582e-07, 2.70395e-07, 2.700455e-07, 2.704031e-07, 
    2.70374e-07, 2.70716e-07, 2.706061e-07, 2.714267e-07, 2.70986e-07, 
    2.722374e-07, 2.726935e-07, 2.739807e-07, 2.747686e-07, 2.755703e-07, 
    2.759238e-07, 2.760314e-07, 2.760764e-07,
  2.332964e-07, 2.341776e-07, 2.340064e-07, 2.347166e-07, 2.343228e-07, 
    2.347877e-07, 2.334752e-07, 2.342125e-07, 2.33742e-07, 2.333759e-07, 
    2.360931e-07, 2.347483e-07, 2.374888e-07, 2.366325e-07, 2.387822e-07, 
    2.373555e-07, 2.390697e-07, 2.387413e-07, 2.397297e-07, 2.394467e-07, 
    2.407094e-07, 2.398604e-07, 2.413635e-07, 2.405068e-07, 2.406408e-07, 
    2.398323e-07, 2.350193e-07, 2.359258e-07, 2.349655e-07, 2.350949e-07, 
    2.350369e-07, 2.343309e-07, 2.339748e-07, 2.332291e-07, 2.333646e-07, 
    2.339123e-07, 2.35153e-07, 2.347321e-07, 2.357928e-07, 2.357689e-07, 
    2.369482e-07, 2.364167e-07, 2.383967e-07, 2.378344e-07, 2.394585e-07, 
    2.390503e-07, 2.394393e-07, 2.393214e-07, 2.394408e-07, 2.388421e-07, 
    2.390987e-07, 2.385717e-07, 2.365162e-07, 2.371207e-07, 2.353165e-07, 
    2.342296e-07, 2.335075e-07, 2.329946e-07, 2.330672e-07, 2.332054e-07, 
    2.339155e-07, 2.345828e-07, 2.35091e-07, 2.354308e-07, 2.357654e-07, 
    2.367773e-07, 2.373127e-07, 2.385103e-07, 2.382945e-07, 2.386602e-07, 
    2.390097e-07, 2.39596e-07, 2.394995e-07, 2.397577e-07, 2.386507e-07, 
    2.393865e-07, 2.381715e-07, 2.385039e-07, 2.358558e-07, 2.348457e-07, 
    2.344156e-07, 2.340393e-07, 2.331229e-07, 2.337558e-07, 2.335064e-07, 
    2.340999e-07, 2.344767e-07, 2.342904e-07, 2.354401e-07, 2.349932e-07, 
    2.373445e-07, 2.363325e-07, 2.389689e-07, 2.383388e-07, 2.391199e-07, 
    2.387214e-07, 2.394041e-07, 2.387897e-07, 2.398538e-07, 2.400852e-07, 
    2.399271e-07, 2.405347e-07, 2.387557e-07, 2.394392e-07, 2.342851e-07, 
    2.343155e-07, 2.344572e-07, 2.338344e-07, 2.337963e-07, 2.332254e-07, 
    2.337335e-07, 2.339497e-07, 2.344986e-07, 2.34823e-07, 2.351314e-07, 
    2.35809e-07, 2.36565e-07, 2.376214e-07, 2.383796e-07, 2.388875e-07, 
    2.385762e-07, 2.38851e-07, 2.385437e-07, 2.383997e-07, 2.399985e-07, 
    2.39101e-07, 2.404473e-07, 2.403729e-07, 2.397638e-07, 2.403813e-07, 
    2.343369e-07, 2.34162e-07, 2.335542e-07, 2.340299e-07, 2.331632e-07, 
    2.336484e-07, 2.339271e-07, 2.350024e-07, 2.352387e-07, 2.354575e-07, 
    2.358896e-07, 2.364439e-07, 2.374153e-07, 2.382598e-07, 2.390301e-07, 
    2.389737e-07, 2.389935e-07, 2.391654e-07, 2.387394e-07, 2.392354e-07, 
    2.393185e-07, 2.39101e-07, 2.40363e-07, 2.400026e-07, 2.403713e-07, 
    2.401368e-07, 2.342188e-07, 2.345131e-07, 2.343541e-07, 2.346531e-07, 
    2.344424e-07, 2.353787e-07, 2.356592e-07, 2.369709e-07, 2.364329e-07, 
    2.372891e-07, 2.3652e-07, 2.366563e-07, 2.373167e-07, 2.365616e-07, 
    2.382131e-07, 2.370935e-07, 2.391721e-07, 2.380551e-07, 2.392421e-07, 
    2.390267e-07, 2.393833e-07, 2.397024e-07, 2.401039e-07, 2.40844e-07, 
    2.406727e-07, 2.412914e-07, 2.349518e-07, 2.353331e-07, 2.352997e-07, 
    2.356987e-07, 2.359936e-07, 2.366328e-07, 2.376568e-07, 2.372719e-07, 
    2.379785e-07, 2.381203e-07, 2.370467e-07, 2.377059e-07, 2.355883e-07, 
    2.359307e-07, 2.35727e-07, 2.349818e-07, 2.373604e-07, 2.361404e-07, 
    2.383921e-07, 2.377322e-07, 2.396569e-07, 2.387001e-07, 2.405783e-07, 
    2.413798e-07, 2.421339e-07, 2.430137e-07, 2.355413e-07, 2.352822e-07, 
    2.357462e-07, 2.363874e-07, 2.369823e-07, 2.377724e-07, 2.378533e-07, 
    2.380012e-07, 2.383843e-07, 2.387063e-07, 2.380478e-07, 2.38787e-07, 
    2.360098e-07, 2.374663e-07, 2.351842e-07, 2.358718e-07, 2.363497e-07, 
    2.361402e-07, 2.372279e-07, 2.374841e-07, 2.385241e-07, 2.379867e-07, 
    2.411819e-07, 2.397697e-07, 2.436833e-07, 2.425913e-07, 2.351917e-07, 
    2.355405e-07, 2.367532e-07, 2.361764e-07, 2.378252e-07, 2.382306e-07, 
    2.3856e-07, 2.389808e-07, 2.390263e-07, 2.392756e-07, 2.388671e-07, 
    2.392595e-07, 2.377741e-07, 2.384382e-07, 2.366148e-07, 2.370588e-07, 
    2.368546e-07, 2.366305e-07, 2.373221e-07, 2.380582e-07, 2.380741e-07, 
    2.383099e-07, 2.389739e-07, 2.378319e-07, 2.413637e-07, 2.391839e-07, 
    2.359206e-07, 2.365915e-07, 2.366876e-07, 2.364277e-07, 2.381899e-07, 
    2.375518e-07, 2.392696e-07, 2.388057e-07, 2.395657e-07, 2.391881e-07, 
    2.391325e-07, 2.386473e-07, 2.383451e-07, 2.37581e-07, 2.369589e-07, 
    2.364654e-07, 2.365802e-07, 2.371222e-07, 2.381032e-07, 2.390304e-07, 
    2.388273e-07, 2.395079e-07, 2.377057e-07, 2.384618e-07, 2.381696e-07, 
    2.389313e-07, 2.372616e-07, 2.386831e-07, 2.368979e-07, 2.370546e-07, 
    2.375391e-07, 2.385129e-07, 2.387285e-07, 2.389583e-07, 2.388165e-07, 
    2.381281e-07, 2.380154e-07, 2.375274e-07, 2.373925e-07, 2.370205e-07, 
    2.367123e-07, 2.369938e-07, 2.372894e-07, 2.381285e-07, 2.38884e-07, 
    2.397069e-07, 2.399083e-07, 2.408682e-07, 2.400866e-07, 2.413757e-07, 
    2.402795e-07, 2.421765e-07, 2.387657e-07, 2.402476e-07, 2.375612e-07, 
    2.378511e-07, 2.383749e-07, 2.395755e-07, 2.389277e-07, 2.396854e-07, 
    2.38011e-07, 2.371408e-07, 2.369158e-07, 2.364954e-07, 2.369254e-07, 
    2.368905e-07, 2.373017e-07, 2.371696e-07, 2.381564e-07, 2.376265e-07, 
    2.391311e-07, 2.396794e-07, 2.412265e-07, 2.421734e-07, 2.431365e-07, 
    2.435612e-07, 2.436905e-07, 2.437445e-07,
  2.190337e-07, 2.200033e-07, 2.198149e-07, 2.205965e-07, 2.20163e-07, 
    2.206747e-07, 2.192303e-07, 2.200417e-07, 2.195238e-07, 2.19121e-07, 
    2.221121e-07, 2.206314e-07, 2.236492e-07, 2.227059e-07, 2.250745e-07, 
    2.235024e-07, 2.253914e-07, 2.250293e-07, 2.26119e-07, 2.258069e-07, 
    2.271995e-07, 2.26263e-07, 2.27921e-07, 2.269759e-07, 2.271238e-07, 
    2.262321e-07, 2.209296e-07, 2.219278e-07, 2.208704e-07, 2.210128e-07, 
    2.209489e-07, 2.201719e-07, 2.197801e-07, 2.189596e-07, 2.191086e-07, 
    2.197113e-07, 2.210768e-07, 2.206135e-07, 2.217811e-07, 2.217548e-07, 
    2.230536e-07, 2.224682e-07, 2.246496e-07, 2.240299e-07, 2.258199e-07, 
    2.2537e-07, 2.257988e-07, 2.256688e-07, 2.258005e-07, 2.251405e-07, 
    2.254233e-07, 2.248425e-07, 2.225778e-07, 2.232437e-07, 2.212568e-07, 
    2.200606e-07, 2.192659e-07, 2.187016e-07, 2.187814e-07, 2.189335e-07, 
    2.197148e-07, 2.204492e-07, 2.210085e-07, 2.213825e-07, 2.21751e-07, 
    2.228655e-07, 2.234553e-07, 2.247748e-07, 2.245369e-07, 2.2494e-07, 
    2.253252e-07, 2.259715e-07, 2.258652e-07, 2.261498e-07, 2.249295e-07, 
    2.257406e-07, 2.244013e-07, 2.247677e-07, 2.218508e-07, 2.207385e-07, 
    2.202652e-07, 2.198511e-07, 2.188428e-07, 2.195391e-07, 2.192646e-07, 
    2.199176e-07, 2.203324e-07, 2.201273e-07, 2.213928e-07, 2.209009e-07, 
    2.234902e-07, 2.223755e-07, 2.252803e-07, 2.245857e-07, 2.254467e-07, 
    2.250075e-07, 2.2576e-07, 2.250827e-07, 2.262558e-07, 2.26511e-07, 
    2.263366e-07, 2.270067e-07, 2.250452e-07, 2.257987e-07, 2.201215e-07, 
    2.20155e-07, 2.203108e-07, 2.196256e-07, 2.195837e-07, 2.189555e-07, 
    2.195145e-07, 2.197524e-07, 2.203564e-07, 2.207135e-07, 2.21053e-07, 
    2.217989e-07, 2.226316e-07, 2.237952e-07, 2.246307e-07, 2.251905e-07, 
    2.248473e-07, 2.251503e-07, 2.248116e-07, 2.246528e-07, 2.264154e-07, 
    2.254259e-07, 2.269103e-07, 2.268282e-07, 2.261566e-07, 2.268375e-07, 
    2.201785e-07, 2.19986e-07, 2.193173e-07, 2.198406e-07, 2.188871e-07, 
    2.194208e-07, 2.197277e-07, 2.209111e-07, 2.211711e-07, 2.21412e-07, 
    2.218878e-07, 2.224981e-07, 2.235682e-07, 2.244987e-07, 2.253476e-07, 
    2.252854e-07, 2.253073e-07, 2.254969e-07, 2.250273e-07, 2.25574e-07, 
    2.256657e-07, 2.254258e-07, 2.268172e-07, 2.264199e-07, 2.268265e-07, 
    2.265678e-07, 2.200485e-07, 2.203725e-07, 2.201974e-07, 2.205265e-07, 
    2.202947e-07, 2.213253e-07, 2.216342e-07, 2.230787e-07, 2.224861e-07, 
    2.234292e-07, 2.225819e-07, 2.227321e-07, 2.234598e-07, 2.226278e-07, 
    2.244473e-07, 2.232138e-07, 2.255042e-07, 2.242732e-07, 2.255813e-07, 
    2.253439e-07, 2.25737e-07, 2.260889e-07, 2.265316e-07, 2.273478e-07, 
    2.271589e-07, 2.278413e-07, 2.208552e-07, 2.212751e-07, 2.212382e-07, 
    2.216775e-07, 2.220023e-07, 2.227062e-07, 2.238342e-07, 2.234102e-07, 
    2.241887e-07, 2.243449e-07, 2.231621e-07, 2.238884e-07, 2.215561e-07, 
    2.219331e-07, 2.217087e-07, 2.208883e-07, 2.235078e-07, 2.22164e-07, 
    2.246445e-07, 2.239173e-07, 2.260387e-07, 2.24984e-07, 2.270548e-07, 
    2.279389e-07, 2.287709e-07, 2.29742e-07, 2.215043e-07, 2.21219e-07, 
    2.217298e-07, 2.22436e-07, 2.230912e-07, 2.239616e-07, 2.240507e-07, 
    2.242137e-07, 2.246359e-07, 2.249907e-07, 2.242652e-07, 2.250796e-07, 
    2.220203e-07, 2.236244e-07, 2.211111e-07, 2.218683e-07, 2.223944e-07, 
    2.221637e-07, 2.233617e-07, 2.236439e-07, 2.2479e-07, 2.241977e-07, 
    2.277207e-07, 2.261631e-07, 2.304812e-07, 2.292758e-07, 2.211193e-07, 
    2.215033e-07, 2.228388e-07, 2.222035e-07, 2.240198e-07, 2.244664e-07, 
    2.248295e-07, 2.252934e-07, 2.253435e-07, 2.256183e-07, 2.25168e-07, 
    2.256006e-07, 2.239635e-07, 2.246953e-07, 2.226863e-07, 2.231755e-07, 
    2.229505e-07, 2.227036e-07, 2.234654e-07, 2.242766e-07, 2.24294e-07, 
    2.24554e-07, 2.252861e-07, 2.240271e-07, 2.279214e-07, 2.255175e-07, 
    2.219219e-07, 2.226609e-07, 2.227665e-07, 2.224803e-07, 2.244217e-07, 
    2.237185e-07, 2.256116e-07, 2.251003e-07, 2.259381e-07, 2.255218e-07, 
    2.254605e-07, 2.249257e-07, 2.245926e-07, 2.237507e-07, 2.230654e-07, 
    2.225218e-07, 2.226483e-07, 2.232453e-07, 2.243262e-07, 2.25348e-07, 
    2.251242e-07, 2.258744e-07, 2.238882e-07, 2.247213e-07, 2.243993e-07, 
    2.252388e-07, 2.233989e-07, 2.249654e-07, 2.229981e-07, 2.231707e-07, 
    2.237046e-07, 2.247777e-07, 2.250152e-07, 2.252685e-07, 2.251122e-07, 
    2.243536e-07, 2.242294e-07, 2.236916e-07, 2.235431e-07, 2.231332e-07, 
    2.227937e-07, 2.231038e-07, 2.234295e-07, 2.24354e-07, 2.251866e-07, 
    2.260939e-07, 2.263159e-07, 2.273747e-07, 2.265127e-07, 2.279348e-07, 
    2.267256e-07, 2.288182e-07, 2.250564e-07, 2.266902e-07, 2.237289e-07, 
    2.240482e-07, 2.246256e-07, 2.259491e-07, 2.252348e-07, 2.260701e-07, 
    2.242245e-07, 2.232659e-07, 2.230179e-07, 2.225549e-07, 2.230285e-07, 
    2.2299e-07, 2.23443e-07, 2.232974e-07, 2.243847e-07, 2.238008e-07, 
    2.25459e-07, 2.260636e-07, 2.277697e-07, 2.288146e-07, 2.298775e-07, 
    2.303464e-07, 2.304891e-07, 2.305487e-07,
  2.100142e-07, 2.110117e-07, 2.108178e-07, 2.116223e-07, 2.11176e-07, 
    2.117028e-07, 2.102165e-07, 2.110513e-07, 2.105184e-07, 2.10104e-07, 
    2.131831e-07, 2.116581e-07, 2.14767e-07, 2.137947e-07, 2.162371e-07, 
    2.146157e-07, 2.16564e-07, 2.161904e-07, 2.173149e-07, 2.169928e-07, 
    2.184308e-07, 2.174636e-07, 2.191762e-07, 2.181999e-07, 2.183526e-07, 
    2.174317e-07, 2.119651e-07, 2.129933e-07, 2.119042e-07, 2.120508e-07, 
    2.11985e-07, 2.111852e-07, 2.107821e-07, 2.09938e-07, 2.100912e-07, 
    2.107113e-07, 2.121167e-07, 2.116397e-07, 2.12842e-07, 2.128148e-07, 
    2.14153e-07, 2.135497e-07, 2.157986e-07, 2.151595e-07, 2.170062e-07, 
    2.165418e-07, 2.169844e-07, 2.168502e-07, 2.169861e-07, 2.163051e-07, 
    2.165969e-07, 2.159975e-07, 2.136627e-07, 2.143489e-07, 2.12302e-07, 
    2.110708e-07, 2.102531e-07, 2.096727e-07, 2.097547e-07, 2.099111e-07, 
    2.107149e-07, 2.114705e-07, 2.120463e-07, 2.124315e-07, 2.128109e-07, 
    2.139593e-07, 2.145671e-07, 2.159278e-07, 2.156823e-07, 2.160982e-07, 
    2.164956e-07, 2.171627e-07, 2.170529e-07, 2.173468e-07, 2.160873e-07, 
    2.169244e-07, 2.155425e-07, 2.159204e-07, 2.129139e-07, 2.117684e-07, 
    2.112813e-07, 2.108551e-07, 2.098178e-07, 2.105341e-07, 2.102518e-07, 
    2.109235e-07, 2.113504e-07, 2.111393e-07, 2.12442e-07, 2.119355e-07, 
    2.146031e-07, 2.134542e-07, 2.164493e-07, 2.157327e-07, 2.16621e-07, 
    2.161678e-07, 2.169444e-07, 2.162454e-07, 2.174562e-07, 2.177198e-07, 
    2.175396e-07, 2.182316e-07, 2.162067e-07, 2.169844e-07, 2.111334e-07, 
    2.111678e-07, 2.113282e-07, 2.106231e-07, 2.105799e-07, 2.099338e-07, 
    2.105088e-07, 2.107536e-07, 2.113751e-07, 2.117427e-07, 2.120921e-07, 
    2.128603e-07, 2.137182e-07, 2.149176e-07, 2.157792e-07, 2.163566e-07, 
    2.160025e-07, 2.163152e-07, 2.159657e-07, 2.158019e-07, 2.17621e-07, 
    2.165996e-07, 2.181321e-07, 2.180473e-07, 2.173538e-07, 2.180568e-07, 
    2.111919e-07, 2.109938e-07, 2.103059e-07, 2.108443e-07, 2.098634e-07, 
    2.104125e-07, 2.107281e-07, 2.119461e-07, 2.122137e-07, 2.124618e-07, 
    2.129518e-07, 2.135806e-07, 2.146835e-07, 2.156429e-07, 2.165188e-07, 
    2.164546e-07, 2.164772e-07, 2.166728e-07, 2.161882e-07, 2.167523e-07, 
    2.16847e-07, 2.165995e-07, 2.180359e-07, 2.176256e-07, 2.180455e-07, 
    2.177783e-07, 2.110582e-07, 2.113916e-07, 2.112115e-07, 2.115502e-07, 
    2.113115e-07, 2.123726e-07, 2.126907e-07, 2.141789e-07, 2.135682e-07, 
    2.145402e-07, 2.136669e-07, 2.138217e-07, 2.145718e-07, 2.137141e-07, 
    2.1559e-07, 2.143182e-07, 2.166804e-07, 2.154105e-07, 2.1676e-07, 
    2.16515e-07, 2.169206e-07, 2.172839e-07, 2.177409e-07, 2.18584e-07, 
    2.183888e-07, 2.190939e-07, 2.118885e-07, 2.123209e-07, 2.122828e-07, 
    2.127352e-07, 2.130698e-07, 2.137949e-07, 2.149577e-07, 2.145205e-07, 
    2.153232e-07, 2.154843e-07, 2.142648e-07, 2.150136e-07, 2.126102e-07, 
    2.129985e-07, 2.127673e-07, 2.119226e-07, 2.146212e-07, 2.132364e-07, 
    2.157934e-07, 2.150434e-07, 2.172321e-07, 2.161437e-07, 2.182813e-07, 
    2.191949e-07, 2.200547e-07, 2.210592e-07, 2.125568e-07, 2.122631e-07, 
    2.12789e-07, 2.135166e-07, 2.141917e-07, 2.150891e-07, 2.151809e-07, 
    2.15349e-07, 2.157844e-07, 2.161505e-07, 2.154021e-07, 2.162422e-07, 
    2.130885e-07, 2.147414e-07, 2.12152e-07, 2.129318e-07, 2.134738e-07, 
    2.13236e-07, 2.144705e-07, 2.147615e-07, 2.159435e-07, 2.153325e-07, 
    2.189694e-07, 2.173606e-07, 2.21824e-07, 2.20577e-07, 2.121604e-07, 
    2.125558e-07, 2.139317e-07, 2.132771e-07, 2.15149e-07, 2.156097e-07, 
    2.159842e-07, 2.164629e-07, 2.165146e-07, 2.167981e-07, 2.163334e-07, 
    2.167798e-07, 2.15091e-07, 2.158457e-07, 2.137744e-07, 2.142786e-07, 
    2.140467e-07, 2.137923e-07, 2.145775e-07, 2.154139e-07, 2.154318e-07, 
    2.157e-07, 2.164555e-07, 2.151566e-07, 2.191769e-07, 2.166943e-07, 
    2.129869e-07, 2.137483e-07, 2.138571e-07, 2.135622e-07, 2.155635e-07, 
    2.148384e-07, 2.167912e-07, 2.162635e-07, 2.171282e-07, 2.166985e-07, 
    2.166353e-07, 2.160834e-07, 2.157398e-07, 2.148717e-07, 2.141652e-07, 
    2.13605e-07, 2.137352e-07, 2.143506e-07, 2.154651e-07, 2.165192e-07, 
    2.162883e-07, 2.170624e-07, 2.150133e-07, 2.158726e-07, 2.155405e-07, 
    2.164064e-07, 2.145089e-07, 2.161247e-07, 2.140958e-07, 2.142737e-07, 
    2.14824e-07, 2.159309e-07, 2.161758e-07, 2.164372e-07, 2.162759e-07, 
    2.154934e-07, 2.153652e-07, 2.148107e-07, 2.146575e-07, 2.14235e-07, 
    2.138851e-07, 2.142048e-07, 2.145404e-07, 2.154937e-07, 2.163527e-07, 
    2.17289e-07, 2.175182e-07, 2.186119e-07, 2.177215e-07, 2.191908e-07, 
    2.179416e-07, 2.201039e-07, 2.162184e-07, 2.179049e-07, 2.148491e-07, 
    2.151784e-07, 2.157739e-07, 2.171396e-07, 2.164024e-07, 2.172646e-07, 
    2.153602e-07, 2.143719e-07, 2.141162e-07, 2.13639e-07, 2.141271e-07, 
    2.140874e-07, 2.145544e-07, 2.144043e-07, 2.155254e-07, 2.149232e-07, 
    2.166337e-07, 2.172578e-07, 2.1902e-07, 2.201e-07, 2.211992e-07, 
    2.216844e-07, 2.218321e-07, 2.218938e-07,
  2.030062e-07, 2.03953e-07, 2.037689e-07, 2.045329e-07, 2.04109e-07, 
    2.046094e-07, 2.03198e-07, 2.039906e-07, 2.034846e-07, 2.030913e-07, 
    2.060171e-07, 2.04567e-07, 2.075249e-07, 2.065989e-07, 2.089264e-07, 
    2.073808e-07, 2.092382e-07, 2.088817e-07, 2.09955e-07, 2.096474e-07, 
    2.110213e-07, 2.10097e-07, 2.11734e-07, 2.108005e-07, 2.109465e-07, 
    2.100665e-07, 2.048587e-07, 2.058365e-07, 2.048008e-07, 2.049402e-07, 
    2.048776e-07, 2.041178e-07, 2.037351e-07, 2.029338e-07, 2.030792e-07, 
    2.036677e-07, 2.050028e-07, 2.045495e-07, 2.056923e-07, 2.056665e-07, 
    2.069401e-07, 2.063657e-07, 2.085081e-07, 2.078988e-07, 2.096603e-07, 
    2.09217e-07, 2.096395e-07, 2.095113e-07, 2.096411e-07, 2.089912e-07, 
    2.092696e-07, 2.086978e-07, 2.064732e-07, 2.071266e-07, 2.051789e-07, 
    2.040092e-07, 2.032328e-07, 2.026821e-07, 2.0276e-07, 2.029084e-07, 
    2.036712e-07, 2.043888e-07, 2.049359e-07, 2.05302e-07, 2.056628e-07, 
    2.067557e-07, 2.073345e-07, 2.086313e-07, 2.083972e-07, 2.087939e-07, 
    2.09173e-07, 2.098097e-07, 2.097049e-07, 2.099855e-07, 2.087834e-07, 
    2.095822e-07, 2.082638e-07, 2.086243e-07, 2.05761e-07, 2.046718e-07, 
    2.042091e-07, 2.038042e-07, 2.028198e-07, 2.034996e-07, 2.032316e-07, 
    2.038692e-07, 2.042746e-07, 2.040741e-07, 2.05312e-07, 2.048306e-07, 
    2.073688e-07, 2.062749e-07, 2.091287e-07, 2.084452e-07, 2.092926e-07, 
    2.088602e-07, 2.096013e-07, 2.089343e-07, 2.100899e-07, 2.103417e-07, 
    2.101696e-07, 2.108307e-07, 2.088973e-07, 2.096395e-07, 2.040685e-07, 
    2.041012e-07, 2.042535e-07, 2.03584e-07, 2.035431e-07, 2.029298e-07, 
    2.034755e-07, 2.037079e-07, 2.042981e-07, 2.046473e-07, 2.049794e-07, 
    2.057098e-07, 2.065261e-07, 2.076683e-07, 2.084895e-07, 2.090403e-07, 
    2.087026e-07, 2.090008e-07, 2.086674e-07, 2.085112e-07, 2.102474e-07, 
    2.092722e-07, 2.107356e-07, 2.106546e-07, 2.099922e-07, 2.106637e-07, 
    2.041241e-07, 2.03936e-07, 2.03283e-07, 2.03794e-07, 2.02863e-07, 
    2.033841e-07, 2.036838e-07, 2.048407e-07, 2.05095e-07, 2.053309e-07, 
    2.057968e-07, 2.063951e-07, 2.074453e-07, 2.083597e-07, 2.09195e-07, 
    2.091338e-07, 2.091553e-07, 2.09342e-07, 2.088797e-07, 2.09418e-07, 
    2.095083e-07, 2.092721e-07, 2.106437e-07, 2.102517e-07, 2.106529e-07, 
    2.103976e-07, 2.039971e-07, 2.043138e-07, 2.041427e-07, 2.044644e-07, 
    2.042378e-07, 2.052461e-07, 2.055485e-07, 2.069647e-07, 2.063833e-07, 
    2.073088e-07, 2.064773e-07, 2.066246e-07, 2.07339e-07, 2.065222e-07, 
    2.083093e-07, 2.070975e-07, 2.093493e-07, 2.081382e-07, 2.094252e-07, 
    2.091914e-07, 2.095786e-07, 2.099254e-07, 2.103619e-07, 2.111677e-07, 
    2.10981e-07, 2.116552e-07, 2.047859e-07, 2.051969e-07, 2.051607e-07, 
    2.055909e-07, 2.059091e-07, 2.065991e-07, 2.077066e-07, 2.0729e-07, 
    2.080548e-07, 2.082084e-07, 2.070465e-07, 2.077598e-07, 2.05472e-07, 
    2.058413e-07, 2.056214e-07, 2.048183e-07, 2.07386e-07, 2.060677e-07, 
    2.085031e-07, 2.077881e-07, 2.098759e-07, 2.088372e-07, 2.108783e-07, 
    2.117519e-07, 2.125746e-07, 2.135369e-07, 2.054212e-07, 2.051419e-07, 
    2.05642e-07, 2.063343e-07, 2.069769e-07, 2.078317e-07, 2.079192e-07, 
    2.080794e-07, 2.084945e-07, 2.088437e-07, 2.081301e-07, 2.089312e-07, 
    2.059271e-07, 2.075005e-07, 2.050363e-07, 2.057779e-07, 2.062935e-07, 
    2.060672e-07, 2.072424e-07, 2.075195e-07, 2.086463e-07, 2.080637e-07, 
    2.115363e-07, 2.099987e-07, 2.1427e-07, 2.130748e-07, 2.050443e-07, 
    2.054202e-07, 2.067293e-07, 2.061063e-07, 2.078888e-07, 2.08328e-07, 
    2.086851e-07, 2.091417e-07, 2.09191e-07, 2.094617e-07, 2.090182e-07, 
    2.094442e-07, 2.078336e-07, 2.08553e-07, 2.065796e-07, 2.070596e-07, 
    2.068388e-07, 2.065966e-07, 2.073443e-07, 2.081414e-07, 2.081584e-07, 
    2.084141e-07, 2.09135e-07, 2.07896e-07, 2.117349e-07, 2.093628e-07, 
    2.058302e-07, 2.065548e-07, 2.066583e-07, 2.063776e-07, 2.082839e-07, 
    2.075929e-07, 2.094551e-07, 2.089515e-07, 2.097767e-07, 2.093666e-07, 
    2.093063e-07, 2.087797e-07, 2.084521e-07, 2.076246e-07, 2.069516e-07, 
    2.064183e-07, 2.065423e-07, 2.071282e-07, 2.081901e-07, 2.091955e-07, 
    2.089752e-07, 2.09714e-07, 2.077595e-07, 2.085787e-07, 2.08262e-07, 
    2.090879e-07, 2.072789e-07, 2.088193e-07, 2.068855e-07, 2.070549e-07, 
    2.075791e-07, 2.086343e-07, 2.088678e-07, 2.091172e-07, 2.089633e-07, 
    2.082171e-07, 2.080949e-07, 2.075664e-07, 2.074205e-07, 2.07018e-07, 
    2.066849e-07, 2.069893e-07, 2.07309e-07, 2.082174e-07, 2.090366e-07, 
    2.099303e-07, 2.101492e-07, 2.111945e-07, 2.103435e-07, 2.117481e-07, 
    2.105539e-07, 2.126219e-07, 2.089086e-07, 2.105187e-07, 2.07603e-07, 
    2.079168e-07, 2.084846e-07, 2.097877e-07, 2.09084e-07, 2.09907e-07, 
    2.080901e-07, 2.071485e-07, 2.069049e-07, 2.064507e-07, 2.069153e-07, 
    2.068775e-07, 2.073222e-07, 2.071793e-07, 2.082476e-07, 2.076736e-07, 
    2.093048e-07, 2.099005e-07, 2.115845e-07, 2.12618e-07, 2.13671e-07, 
    2.141361e-07, 2.142777e-07, 2.143369e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 HTOP =
  0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 0.2360823, 
    0.2360823, 0.2360823 ;

 INT_SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAISHA =
  0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503, 0.001095503, 0.001095503, 
    0.001095503, 0.001095503, 0.001095503 ;

 LAISUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LAKEICEFRAC =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAKEICETHICK =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 LAND_UPTAKE =
  6.191209e-08, 6.218511e-08, 6.213204e-08, 6.235225e-08, 6.22301e-08, 
    6.237429e-08, 6.196745e-08, 6.219594e-08, 6.205008e-08, 6.193667e-08, 
    6.277961e-08, 6.236208e-08, 6.321343e-08, 6.29471e-08, 6.361618e-08, 
    6.317198e-08, 6.370576e-08, 6.360339e-08, 6.391155e-08, 6.382326e-08, 
    6.421742e-08, 6.39523e-08, 6.442178e-08, 6.415411e-08, 6.419598e-08, 
    6.394355e-08, 6.244612e-08, 6.272763e-08, 6.242944e-08, 6.246958e-08, 
    6.245157e-08, 6.223262e-08, 6.212228e-08, 6.189123e-08, 6.193318e-08, 
    6.210288e-08, 6.248763e-08, 6.235703e-08, 6.26862e-08, 6.267877e-08, 
    6.304526e-08, 6.288002e-08, 6.349605e-08, 6.332096e-08, 6.382695e-08, 
    6.369969e-08, 6.382097e-08, 6.37842e-08, 6.382145e-08, 6.363481e-08, 
    6.371478e-08, 6.355055e-08, 6.291096e-08, 6.309892e-08, 6.253835e-08, 
    6.220129e-08, 6.197747e-08, 6.181863e-08, 6.184109e-08, 6.188389e-08, 
    6.210387e-08, 6.231072e-08, 6.246836e-08, 6.25738e-08, 6.267771e-08, 
    6.299219e-08, 6.315867e-08, 6.353144e-08, 6.346419e-08, 6.357814e-08, 
    6.368703e-08, 6.386984e-08, 6.383975e-08, 6.392029e-08, 6.357515e-08, 
    6.380452e-08, 6.342587e-08, 6.352943e-08, 6.27059e-08, 6.239227e-08, 
    6.225892e-08, 6.214224e-08, 6.185834e-08, 6.205439e-08, 6.19771e-08, 
    6.216099e-08, 6.227782e-08, 6.222004e-08, 6.257669e-08, 6.243803e-08, 
    6.316854e-08, 6.285387e-08, 6.367434e-08, 6.347799e-08, 6.372139e-08, 
    6.359719e-08, 6.381001e-08, 6.361848e-08, 6.395027e-08, 6.402251e-08, 
    6.397314e-08, 6.41628e-08, 6.360786e-08, 6.382096e-08, 6.221842e-08, 
    6.222784e-08, 6.227175e-08, 6.207874e-08, 6.206693e-08, 6.189008e-08, 
    6.204745e-08, 6.211446e-08, 6.22846e-08, 6.238523e-08, 6.248089e-08, 
    6.269123e-08, 6.292615e-08, 6.325467e-08, 6.349072e-08, 6.364895e-08, 
    6.355192e-08, 6.363758e-08, 6.354183e-08, 6.349695e-08, 6.399544e-08, 
    6.371552e-08, 6.413553e-08, 6.411229e-08, 6.39222e-08, 6.411491e-08, 
    6.223446e-08, 6.218023e-08, 6.199193e-08, 6.213929e-08, 6.187082e-08, 
    6.202109e-08, 6.210749e-08, 6.244091e-08, 6.251418e-08, 6.258211e-08, 
    6.271628e-08, 6.288847e-08, 6.319055e-08, 6.34534e-08, 6.369337e-08, 
    6.367579e-08, 6.368198e-08, 6.373558e-08, 6.36028e-08, 6.375738e-08, 
    6.378333e-08, 6.371549e-08, 6.410917e-08, 6.39967e-08, 6.411179e-08, 
    6.403856e-08, 6.219786e-08, 6.228911e-08, 6.22398e-08, 6.233252e-08, 
    6.22672e-08, 6.255767e-08, 6.264477e-08, 6.305234e-08, 6.288508e-08, 
    6.315129e-08, 6.291213e-08, 6.29545e-08, 6.315996e-08, 6.292505e-08, 
    6.34389e-08, 6.30905e-08, 6.373767e-08, 6.338972e-08, 6.375947e-08, 
    6.369233e-08, 6.38035e-08, 6.390305e-08, 6.402831e-08, 6.425942e-08, 
    6.420591e-08, 6.43992e-08, 6.242516e-08, 6.254352e-08, 6.25331e-08, 
    6.265698e-08, 6.27486e-08, 6.294718e-08, 6.326568e-08, 6.314591e-08, 
    6.33658e-08, 6.340995e-08, 6.307588e-08, 6.328098e-08, 6.262274e-08, 
    6.272907e-08, 6.266577e-08, 6.243449e-08, 6.317349e-08, 6.279422e-08, 
    6.349462e-08, 6.328914e-08, 6.388886e-08, 6.359058e-08, 6.417645e-08, 
    6.442689e-08, 6.466265e-08, 6.493813e-08, 6.260812e-08, 6.25277e-08, 
    6.267172e-08, 6.287096e-08, 6.305586e-08, 6.330166e-08, 6.332682e-08, 
    6.337287e-08, 6.349217e-08, 6.359246e-08, 6.338743e-08, 6.361761e-08, 
    6.275372e-08, 6.320642e-08, 6.249729e-08, 6.27108e-08, 6.285921e-08, 
    6.279412e-08, 6.313223e-08, 6.321191e-08, 6.353574e-08, 6.336835e-08, 
    6.436507e-08, 6.392407e-08, 6.514793e-08, 6.480587e-08, 6.249959e-08, 
    6.260785e-08, 6.298463e-08, 6.280536e-08, 6.331808e-08, 6.344429e-08, 
    6.35469e-08, 6.367805e-08, 6.369222e-08, 6.376993e-08, 6.364259e-08, 
    6.376491e-08, 6.330219e-08, 6.350896e-08, 6.294157e-08, 6.307966e-08, 
    6.301614e-08, 6.294646e-08, 6.316152e-08, 6.339064e-08, 6.339556e-08, 
    6.346902e-08, 6.367603e-08, 6.332016e-08, 6.442196e-08, 6.374147e-08, 
    6.27259e-08, 6.293441e-08, 6.296421e-08, 6.288344e-08, 6.343164e-08, 
    6.3233e-08, 6.376804e-08, 6.362344e-08, 6.386038e-08, 6.374263e-08, 
    6.372531e-08, 6.357409e-08, 6.347994e-08, 6.32421e-08, 6.304859e-08, 
    6.289515e-08, 6.293084e-08, 6.309938e-08, 6.340467e-08, 6.36935e-08, 
    6.363022e-08, 6.384236e-08, 6.32809e-08, 6.351632e-08, 6.342533e-08, 
    6.36626e-08, 6.314273e-08, 6.358538e-08, 6.302958e-08, 6.307831e-08, 
    6.322905e-08, 6.353228e-08, 6.359939e-08, 6.367102e-08, 6.362682e-08, 
    6.341242e-08, 6.33773e-08, 6.322539e-08, 6.318344e-08, 6.30677e-08, 
    6.297188e-08, 6.305942e-08, 6.315137e-08, 6.341251e-08, 6.364786e-08, 
    6.390447e-08, 6.396727e-08, 6.426707e-08, 6.4023e-08, 6.442575e-08, 
    6.40833e-08, 6.467612e-08, 6.361105e-08, 6.407326e-08, 6.323592e-08, 
    6.332613e-08, 6.348927e-08, 6.386351e-08, 6.366148e-08, 6.389776e-08, 
    6.337593e-08, 6.310519e-08, 6.303516e-08, 6.290448e-08, 6.303815e-08, 
    6.302728e-08, 6.315518e-08, 6.311409e-08, 6.342119e-08, 6.325622e-08, 
    6.372487e-08, 6.38959e-08, 6.437893e-08, 6.467506e-08, 6.497654e-08, 
    6.510964e-08, 6.515015e-08, 6.516709e-08 ;

 LAND_USE_FLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC =
  0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 0.1428203, 
    0.1428203, 0.1428203 ;

 LEAFC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LEAFC_LOSS =
  8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 8.453843e-10, 
    8.453843e-10, 8.453843e-10, 8.453843e-10 ;

 LEAFN =
  0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507, 0.003570507, 0.003570507, 
    0.003570507, 0.003570507, 0.003570507 ;

 LEAF_MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LFC2 =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LF_CONV_CFLUX =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITFALL =
  1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 1.322617e-09, 
    1.322617e-09, 1.322617e-09, 1.322617e-09 ;

 LITHR =
  9.581084e-13, 9.607331e-13, 9.602232e-13, 9.623386e-13, 9.611656e-13, 
    9.625504e-13, 9.58641e-13, 9.608369e-13, 9.594355e-13, 9.583453e-13, 
    9.664388e-13, 9.62433e-13, 9.705987e-13, 9.680471e-13, 9.744543e-13, 
    9.702012e-13, 9.753114e-13, 9.743327e-13, 9.772797e-13, 9.764358e-13, 
    9.802e-13, 9.776691e-13, 9.82151e-13, 9.795963e-13, 9.799957e-13, 
    9.775854e-13, 9.632404e-13, 9.659401e-13, 9.630803e-13, 9.634654e-13, 
    9.632928e-13, 9.611896e-13, 9.601286e-13, 9.579082e-13, 9.583117e-13, 
    9.599426e-13, 9.636387e-13, 9.623851e-13, 9.655452e-13, 9.65474e-13, 
    9.689881e-13, 9.674041e-13, 9.733056e-13, 9.716297e-13, 9.764711e-13, 
    9.752541e-13, 9.764137e-13, 9.760622e-13, 9.764183e-13, 9.746334e-13, 
    9.753981e-13, 9.738274e-13, 9.677006e-13, 9.695021e-13, 9.641258e-13, 
    9.608874e-13, 9.587372e-13, 9.572099e-13, 9.574259e-13, 9.578373e-13, 
    9.599522e-13, 9.619403e-13, 9.634543e-13, 9.644665e-13, 9.654637e-13, 
    9.684779e-13, 9.700742e-13, 9.736439e-13, 9.730008e-13, 9.740908e-13, 
    9.75133e-13, 9.768808e-13, 9.765933e-13, 9.773628e-13, 9.740626e-13, 
    9.762561e-13, 9.726342e-13, 9.736252e-13, 9.657315e-13, 9.627235e-13, 
    9.614413e-13, 9.603211e-13, 9.575918e-13, 9.594766e-13, 9.587336e-13, 
    9.605016e-13, 9.616241e-13, 9.610692e-13, 9.644942e-13, 9.631629e-13, 
    9.701687e-13, 9.671529e-13, 9.750114e-13, 9.731329e-13, 9.754617e-13, 
    9.742737e-13, 9.763087e-13, 9.744773e-13, 9.776495e-13, 9.783394e-13, 
    9.778679e-13, 9.796799e-13, 9.743756e-13, 9.764134e-13, 9.610535e-13, 
    9.611439e-13, 9.61566e-13, 9.597106e-13, 9.595973e-13, 9.578971e-13, 
    9.594102e-13, 9.600541e-13, 9.616895e-13, 9.626558e-13, 9.635744e-13, 
    9.655932e-13, 9.678459e-13, 9.709942e-13, 9.732547e-13, 9.747688e-13, 
    9.738407e-13, 9.7466e-13, 9.737439e-13, 9.733145e-13, 9.780807e-13, 
    9.754051e-13, 9.794193e-13, 9.791974e-13, 9.77381e-13, 9.792225e-13, 
    9.612076e-13, 9.606866e-13, 9.588764e-13, 9.602932e-13, 9.577119e-13, 
    9.591566e-13, 9.599868e-13, 9.6319e-13, 9.638942e-13, 9.64546e-13, 
    9.658337e-13, 9.674852e-13, 9.7038e-13, 9.728972e-13, 9.751938e-13, 
    9.750256e-13, 9.750848e-13, 9.755972e-13, 9.743272e-13, 9.758057e-13, 
    9.760535e-13, 9.754052e-13, 9.791677e-13, 9.780933e-13, 9.791927e-13, 
    9.784933e-13, 9.608561e-13, 9.617326e-13, 9.61259e-13, 9.621495e-13, 
    9.615219e-13, 9.643109e-13, 9.651466e-13, 9.690552e-13, 9.674525e-13, 
    9.700038e-13, 9.67712e-13, 9.681181e-13, 9.700857e-13, 9.678362e-13, 
    9.727578e-13, 9.694207e-13, 9.756172e-13, 9.722864e-13, 9.758256e-13, 
    9.751838e-13, 9.762469e-13, 9.771981e-13, 9.783952e-13, 9.806018e-13, 
    9.800911e-13, 9.819359e-13, 9.630393e-13, 9.641754e-13, 9.640759e-13, 
    9.652648e-13, 9.661435e-13, 9.680481e-13, 9.710999e-13, 9.69953e-13, 
    9.720591e-13, 9.724815e-13, 9.692819e-13, 9.712463e-13, 9.649358e-13, 
    9.659555e-13, 9.653489e-13, 9.631287e-13, 9.702164e-13, 9.665804e-13, 
    9.732919e-13, 9.713247e-13, 9.770625e-13, 9.742096e-13, 9.798098e-13, 
    9.821989e-13, 9.844485e-13, 9.870719e-13, 9.647957e-13, 9.64024e-13, 
    9.654062e-13, 9.673165e-13, 9.690897e-13, 9.714446e-13, 9.716858e-13, 
    9.721266e-13, 9.732687e-13, 9.742284e-13, 9.722653e-13, 9.74469e-13, 
    9.661908e-13, 9.705321e-13, 9.637317e-13, 9.657801e-13, 9.672042e-13, 
    9.665802e-13, 9.698219e-13, 9.705853e-13, 9.736852e-13, 9.720834e-13, 
    9.816089e-13, 9.773983e-13, 9.890697e-13, 9.858125e-13, 9.637543e-13, 
    9.647933e-13, 9.684067e-13, 9.666881e-13, 9.716021e-13, 9.728103e-13, 
    9.737926e-13, 9.750469e-13, 9.751826e-13, 9.759256e-13, 9.747079e-13, 
    9.758778e-13, 9.714496e-13, 9.734293e-13, 9.679946e-13, 9.693178e-13, 
    9.687094e-13, 9.680413e-13, 9.701026e-13, 9.72296e-13, 9.72344e-13, 
    9.730467e-13, 9.750247e-13, 9.71622e-13, 9.821501e-13, 9.756509e-13, 
    9.659261e-13, 9.679249e-13, 9.682114e-13, 9.674372e-13, 9.726891e-13, 
    9.70787e-13, 9.759076e-13, 9.745247e-13, 9.767905e-13, 9.756648e-13, 
    9.75499e-13, 9.740527e-13, 9.731516e-13, 9.708741e-13, 9.6902e-13, 
    9.675496e-13, 9.678916e-13, 9.695067e-13, 9.724305e-13, 9.751945e-13, 
    9.745891e-13, 9.766184e-13, 9.71246e-13, 9.734994e-13, 9.726283e-13, 
    9.748992e-13, 9.699222e-13, 9.741579e-13, 9.688383e-13, 9.693053e-13, 
    9.707492e-13, 9.736515e-13, 9.742946e-13, 9.749795e-13, 9.745571e-13, 
    9.725048e-13, 9.721689e-13, 9.707144e-13, 9.703122e-13, 9.692037e-13, 
    9.682851e-13, 9.691241e-13, 9.700048e-13, 9.72506e-13, 9.747579e-13, 
    9.772116e-13, 9.778121e-13, 9.806733e-13, 9.783431e-13, 9.821861e-13, 
    9.78917e-13, 9.845746e-13, 9.744047e-13, 9.788228e-13, 9.708152e-13, 
    9.716791e-13, 9.732402e-13, 9.768193e-13, 9.748886e-13, 9.77147e-13, 
    9.721557e-13, 9.695619e-13, 9.688916e-13, 9.676388e-13, 9.689203e-13, 
    9.688162e-13, 9.700419e-13, 9.696481e-13, 9.725891e-13, 9.710097e-13, 
    9.754946e-13, 9.771293e-13, 9.817422e-13, 9.845659e-13, 9.874389e-13, 
    9.887056e-13, 9.890913e-13, 9.892524e-13 ;

 LITR1C =
  3.066879e-05, 3.066867e-05, 3.06687e-05, 3.06686e-05, 3.066865e-05, 
    3.066859e-05, 3.066877e-05, 3.066867e-05, 3.066873e-05, 3.066878e-05, 
    3.066842e-05, 3.066859e-05, 3.066823e-05, 3.066834e-05, 3.066805e-05, 
    3.066825e-05, 3.066802e-05, 3.066806e-05, 3.066792e-05, 3.066796e-05, 
    3.066779e-05, 3.066791e-05, 3.066771e-05, 3.066782e-05, 3.06678e-05, 
    3.066791e-05, 3.066856e-05, 3.066844e-05, 3.066857e-05, 3.066855e-05, 
    3.066856e-05, 3.066865e-05, 3.06687e-05, 3.06688e-05, 3.066878e-05, 
    3.066871e-05, 3.066854e-05, 3.06686e-05, 3.066846e-05, 3.066846e-05, 
    3.06683e-05, 3.066837e-05, 3.066811e-05, 3.066818e-05, 3.066796e-05, 
    3.066802e-05, 3.066796e-05, 3.066798e-05, 3.066796e-05, 3.066804e-05, 
    3.066801e-05, 3.066808e-05, 3.066836e-05, 3.066828e-05, 3.066852e-05, 
    3.066867e-05, 3.066876e-05, 3.066883e-05, 3.066882e-05, 3.066881e-05, 
    3.066871e-05, 3.066862e-05, 3.066855e-05, 3.06685e-05, 3.066846e-05, 
    3.066832e-05, 3.066825e-05, 3.066809e-05, 3.066812e-05, 3.066807e-05, 
    3.066802e-05, 3.066794e-05, 3.066796e-05, 3.066792e-05, 3.066807e-05, 
    3.066797e-05, 3.066814e-05, 3.066809e-05, 3.066845e-05, 3.066858e-05, 
    3.066864e-05, 3.066869e-05, 3.066882e-05, 3.066873e-05, 3.066876e-05, 
    3.066868e-05, 3.066863e-05, 3.066866e-05, 3.06685e-05, 3.066856e-05, 
    3.066825e-05, 3.066838e-05, 3.066803e-05, 3.066811e-05, 3.066801e-05, 
    3.066806e-05, 3.066797e-05, 3.066805e-05, 3.066791e-05, 3.066788e-05, 
    3.06679e-05, 3.066782e-05, 3.066806e-05, 3.066796e-05, 3.066866e-05, 
    3.066865e-05, 3.066863e-05, 3.066872e-05, 3.066873e-05, 3.06688e-05, 
    3.066873e-05, 3.06687e-05, 3.066863e-05, 3.066859e-05, 3.066854e-05, 
    3.066845e-05, 3.066835e-05, 3.066821e-05, 3.066811e-05, 3.066804e-05, 
    3.066808e-05, 3.066804e-05, 3.066808e-05, 3.06681e-05, 3.066789e-05, 
    3.066801e-05, 3.066783e-05, 3.066784e-05, 3.066792e-05, 3.066784e-05, 
    3.066865e-05, 3.066867e-05, 3.066876e-05, 3.066869e-05, 3.066881e-05, 
    3.066874e-05, 3.066871e-05, 3.066856e-05, 3.066853e-05, 3.06685e-05, 
    3.066844e-05, 3.066837e-05, 3.066824e-05, 3.066812e-05, 3.066802e-05, 
    3.066803e-05, 3.066802e-05, 3.0668e-05, 3.066806e-05, 3.066799e-05, 
    3.066798e-05, 3.066801e-05, 3.066784e-05, 3.066789e-05, 3.066784e-05, 
    3.066787e-05, 3.066867e-05, 3.066863e-05, 3.066865e-05, 3.066861e-05, 
    3.066864e-05, 3.066851e-05, 3.066847e-05, 3.06683e-05, 3.066837e-05, 
    3.066826e-05, 3.066836e-05, 3.066834e-05, 3.066825e-05, 3.066835e-05, 
    3.066813e-05, 3.066828e-05, 3.0668e-05, 3.066815e-05, 3.066799e-05, 
    3.066802e-05, 3.066797e-05, 3.066793e-05, 3.066787e-05, 3.066778e-05, 
    3.06678e-05, 3.066771e-05, 3.066857e-05, 3.066852e-05, 3.066852e-05, 
    3.066847e-05, 3.066843e-05, 3.066834e-05, 3.06682e-05, 3.066826e-05, 
    3.066816e-05, 3.066814e-05, 3.066829e-05, 3.06682e-05, 3.066848e-05, 
    3.066844e-05, 3.066846e-05, 3.066857e-05, 3.066825e-05, 3.066841e-05, 
    3.066811e-05, 3.066819e-05, 3.066794e-05, 3.066806e-05, 3.066781e-05, 
    3.06677e-05, 3.06676e-05, 3.066748e-05, 3.066849e-05, 3.066853e-05, 
    3.066846e-05, 3.066838e-05, 3.06683e-05, 3.066819e-05, 3.066818e-05, 
    3.066816e-05, 3.066811e-05, 3.066806e-05, 3.066815e-05, 3.066805e-05, 
    3.066843e-05, 3.066823e-05, 3.066854e-05, 3.066845e-05, 3.066838e-05, 
    3.066841e-05, 3.066826e-05, 3.066823e-05, 3.066809e-05, 3.066816e-05, 
    3.066773e-05, 3.066792e-05, 3.066739e-05, 3.066754e-05, 3.066854e-05, 
    3.066849e-05, 3.066833e-05, 3.066841e-05, 3.066818e-05, 3.066813e-05, 
    3.066808e-05, 3.066803e-05, 3.066802e-05, 3.066799e-05, 3.066804e-05, 
    3.066799e-05, 3.066819e-05, 3.06681e-05, 3.066834e-05, 3.066829e-05, 
    3.066831e-05, 3.066834e-05, 3.066825e-05, 3.066815e-05, 3.066815e-05, 
    3.066812e-05, 3.066803e-05, 3.066818e-05, 3.066771e-05, 3.0668e-05, 
    3.066844e-05, 3.066835e-05, 3.066834e-05, 3.066837e-05, 3.066813e-05, 
    3.066822e-05, 3.066799e-05, 3.066805e-05, 3.066795e-05, 3.0668e-05, 
    3.0668e-05, 3.066807e-05, 3.066811e-05, 3.066822e-05, 3.06683e-05, 
    3.066837e-05, 3.066835e-05, 3.066828e-05, 3.066814e-05, 3.066802e-05, 
    3.066805e-05, 3.066795e-05, 3.06682e-05, 3.06681e-05, 3.066814e-05, 
    3.066803e-05, 3.066826e-05, 3.066807e-05, 3.066831e-05, 3.066829e-05, 
    3.066822e-05, 3.066809e-05, 3.066806e-05, 3.066803e-05, 3.066805e-05, 
    3.066814e-05, 3.066816e-05, 3.066822e-05, 3.066824e-05, 3.066829e-05, 
    3.066833e-05, 3.066829e-05, 3.066826e-05, 3.066814e-05, 3.066804e-05, 
    3.066793e-05, 3.06679e-05, 3.066777e-05, 3.066788e-05, 3.06677e-05, 
    3.066785e-05, 3.06676e-05, 3.066806e-05, 3.066786e-05, 3.066822e-05, 
    3.066818e-05, 3.066811e-05, 3.066795e-05, 3.066803e-05, 3.066793e-05, 
    3.066816e-05, 3.066827e-05, 3.06683e-05, 3.066836e-05, 3.06683e-05, 
    3.066831e-05, 3.066825e-05, 3.066827e-05, 3.066814e-05, 3.066821e-05, 
    3.0668e-05, 3.066793e-05, 3.066772e-05, 3.06676e-05, 3.066747e-05, 
    3.066741e-05, 3.066739e-05, 3.066739e-05 ;

 LITR1C_TO_SOIL1C =
  6.381433e-13, 6.398912e-13, 6.395517e-13, 6.409603e-13, 6.401793e-13, 
    6.411013e-13, 6.38498e-13, 6.399603e-13, 6.390271e-13, 6.383011e-13, 
    6.436908e-13, 6.410233e-13, 6.464609e-13, 6.447618e-13, 6.490284e-13, 
    6.461962e-13, 6.495991e-13, 6.489474e-13, 6.509099e-13, 6.503479e-13, 
    6.528546e-13, 6.511692e-13, 6.541537e-13, 6.524525e-13, 6.527185e-13, 
    6.511135e-13, 6.415609e-13, 6.433586e-13, 6.414542e-13, 6.417107e-13, 
    6.415958e-13, 6.401951e-13, 6.394886e-13, 6.380101e-13, 6.382787e-13, 
    6.393648e-13, 6.418261e-13, 6.409913e-13, 6.430957e-13, 6.430482e-13, 
    6.453884e-13, 6.443335e-13, 6.482635e-13, 6.471474e-13, 6.503714e-13, 
    6.49561e-13, 6.503332e-13, 6.500992e-13, 6.503362e-13, 6.491476e-13, 
    6.496569e-13, 6.486109e-13, 6.44531e-13, 6.457306e-13, 6.421504e-13, 
    6.39994e-13, 6.385621e-13, 6.37545e-13, 6.376888e-13, 6.379628e-13, 
    6.393712e-13, 6.406951e-13, 6.417033e-13, 6.423773e-13, 6.430414e-13, 
    6.450486e-13, 6.461116e-13, 6.484887e-13, 6.480605e-13, 6.487864e-13, 
    6.494804e-13, 6.506442e-13, 6.504528e-13, 6.509652e-13, 6.487676e-13, 
    6.502282e-13, 6.478164e-13, 6.484762e-13, 6.432197e-13, 6.412166e-13, 
    6.403628e-13, 6.396168e-13, 6.377993e-13, 6.390545e-13, 6.385597e-13, 
    6.397371e-13, 6.404846e-13, 6.40115e-13, 6.423958e-13, 6.415093e-13, 
    6.461746e-13, 6.441663e-13, 6.493994e-13, 6.481484e-13, 6.496992e-13, 
    6.489081e-13, 6.502633e-13, 6.490437e-13, 6.511561e-13, 6.516155e-13, 
    6.513015e-13, 6.525082e-13, 6.48976e-13, 6.50333e-13, 6.401046e-13, 
    6.401648e-13, 6.404458e-13, 6.392103e-13, 6.391348e-13, 6.380026e-13, 
    6.390103e-13, 6.394391e-13, 6.40528e-13, 6.411716e-13, 6.417833e-13, 
    6.431276e-13, 6.446277e-13, 6.467243e-13, 6.482295e-13, 6.492378e-13, 
    6.486198e-13, 6.491654e-13, 6.485553e-13, 6.482694e-13, 6.514433e-13, 
    6.496615e-13, 6.523347e-13, 6.521869e-13, 6.509774e-13, 6.522036e-13, 
    6.402072e-13, 6.398603e-13, 6.386548e-13, 6.395982e-13, 6.378793e-13, 
    6.388414e-13, 6.393942e-13, 6.415273e-13, 6.419962e-13, 6.424303e-13, 
    6.432878e-13, 6.443875e-13, 6.463152e-13, 6.479915e-13, 6.495208e-13, 
    6.494088e-13, 6.494482e-13, 6.497895e-13, 6.489437e-13, 6.499284e-13, 
    6.500933e-13, 6.496616e-13, 6.521671e-13, 6.514517e-13, 6.521838e-13, 
    6.51718e-13, 6.399731e-13, 6.405568e-13, 6.402414e-13, 6.408344e-13, 
    6.404165e-13, 6.422737e-13, 6.428302e-13, 6.454331e-13, 6.443658e-13, 
    6.460647e-13, 6.445386e-13, 6.44809e-13, 6.461192e-13, 6.446212e-13, 
    6.478987e-13, 6.456764e-13, 6.498027e-13, 6.475847e-13, 6.499416e-13, 
    6.495142e-13, 6.502221e-13, 6.508556e-13, 6.516527e-13, 6.531221e-13, 
    6.52782e-13, 6.540105e-13, 6.41427e-13, 6.421834e-13, 6.421172e-13, 
    6.429089e-13, 6.434941e-13, 6.447625e-13, 6.467947e-13, 6.460309e-13, 
    6.474334e-13, 6.477147e-13, 6.455841e-13, 6.468921e-13, 6.426898e-13, 
    6.433689e-13, 6.429649e-13, 6.414864e-13, 6.462063e-13, 6.437851e-13, 
    6.482543e-13, 6.469444e-13, 6.507652e-13, 6.488655e-13, 6.525947e-13, 
    6.541857e-13, 6.556837e-13, 6.574307e-13, 6.425966e-13, 6.420827e-13, 
    6.430031e-13, 6.442752e-13, 6.45456e-13, 6.470242e-13, 6.471848e-13, 
    6.474783e-13, 6.482389e-13, 6.48878e-13, 6.475707e-13, 6.490382e-13, 
    6.435255e-13, 6.464166e-13, 6.41888e-13, 6.432521e-13, 6.442005e-13, 
    6.437849e-13, 6.459436e-13, 6.46452e-13, 6.485162e-13, 6.474496e-13, 
    6.537928e-13, 6.509888e-13, 6.58761e-13, 6.56592e-13, 6.41903e-13, 
    6.42595e-13, 6.450011e-13, 6.438567e-13, 6.471291e-13, 6.479336e-13, 
    6.485877e-13, 6.49423e-13, 6.495134e-13, 6.500082e-13, 6.491973e-13, 
    6.499763e-13, 6.470275e-13, 6.483459e-13, 6.447267e-13, 6.456079e-13, 
    6.452027e-13, 6.447579e-13, 6.461305e-13, 6.475912e-13, 6.476231e-13, 
    6.480911e-13, 6.494083e-13, 6.471423e-13, 6.541532e-13, 6.498252e-13, 
    6.433493e-13, 6.446803e-13, 6.448711e-13, 6.443556e-13, 6.478529e-13, 
    6.465862e-13, 6.499962e-13, 6.490753e-13, 6.505841e-13, 6.498345e-13, 
    6.497241e-13, 6.487609e-13, 6.481609e-13, 6.466443e-13, 6.454096e-13, 
    6.444304e-13, 6.446582e-13, 6.457337e-13, 6.476807e-13, 6.495213e-13, 
    6.491182e-13, 6.504695e-13, 6.468919e-13, 6.483925e-13, 6.478124e-13, 
    6.493247e-13, 6.460104e-13, 6.48831e-13, 6.452886e-13, 6.455995e-13, 
    6.465611e-13, 6.484938e-13, 6.489221e-13, 6.493781e-13, 6.490969e-13, 
    6.477302e-13, 6.475065e-13, 6.465379e-13, 6.462701e-13, 6.455319e-13, 
    6.449202e-13, 6.454789e-13, 6.460654e-13, 6.477311e-13, 6.492306e-13, 
    6.508645e-13, 6.512644e-13, 6.531697e-13, 6.51618e-13, 6.541771e-13, 
    6.520002e-13, 6.557676e-13, 6.489953e-13, 6.519375e-13, 6.466051e-13, 
    6.471804e-13, 6.482198e-13, 6.506033e-13, 6.493176e-13, 6.508215e-13, 
    6.474978e-13, 6.457705e-13, 6.453241e-13, 6.444898e-13, 6.453432e-13, 
    6.452738e-13, 6.460901e-13, 6.458279e-13, 6.477863e-13, 6.467346e-13, 
    6.497212e-13, 6.508098e-13, 6.538816e-13, 6.557618e-13, 6.57675e-13, 
    6.585186e-13, 6.587753e-13, 6.588826e-13 ;

 LITR1C_vr =
  0.00175122, 0.001751213, 0.001751214, 0.001751209, 0.001751212, 
    0.001751208, 0.001751218, 0.001751213, 0.001751216, 0.001751219, 
    0.001751198, 0.001751209, 0.001751187, 0.001751194, 0.001751178, 
    0.001751189, 0.001751175, 0.001751178, 0.00175117, 0.001751172, 
    0.001751163, 0.001751169, 0.001751158, 0.001751164, 0.001751163, 
    0.001751169, 0.001751206, 0.001751199, 0.001751207, 0.001751206, 
    0.001751206, 0.001751212, 0.001751214, 0.00175122, 0.001751219, 
    0.001751215, 0.001751205, 0.001751209, 0.001751201, 0.001751201, 
    0.001751192, 0.001751196, 0.001751181, 0.001751185, 0.001751172, 
    0.001751175, 0.001751172, 0.001751173, 0.001751172, 0.001751177, 
    0.001751175, 0.001751179, 0.001751195, 0.00175119, 0.001751204, 
    0.001751213, 0.001751218, 0.001751222, 0.001751221, 0.00175122, 
    0.001751215, 0.00175121, 0.001751206, 0.001751203, 0.001751201, 
    0.001751193, 0.001751189, 0.00175118, 0.001751181, 0.001751179, 
    0.001751176, 0.001751171, 0.001751172, 0.00175117, 0.001751179, 
    0.001751173, 0.001751182, 0.00175118, 0.0017512, 0.001751208, 
    0.001751211, 0.001751214, 0.001751221, 0.001751216, 0.001751218, 
    0.001751213, 0.001751211, 0.001751212, 0.001751203, 0.001751207, 
    0.001751189, 0.001751196, 0.001751176, 0.001751181, 0.001751175, 
    0.001751178, 0.001751173, 0.001751177, 0.001751169, 0.001751167, 
    0.001751169, 0.001751164, 0.001751178, 0.001751172, 0.001751212, 
    0.001751212, 0.001751211, 0.001751216, 0.001751216, 0.00175122, 
    0.001751216, 0.001751215, 0.00175121, 0.001751208, 0.001751206, 
    0.0017512, 0.001751195, 0.001751186, 0.001751181, 0.001751177, 
    0.001751179, 0.001751177, 0.001751179, 0.001751181, 0.001751168, 
    0.001751175, 0.001751165, 0.001751165, 0.00175117, 0.001751165, 
    0.001751212, 0.001751213, 0.001751218, 0.001751214, 0.001751221, 
    0.001751217, 0.001751215, 0.001751207, 0.001751205, 0.001751203, 
    0.0017512, 0.001751196, 0.001751188, 0.001751182, 0.001751176, 
    0.001751176, 0.001751176, 0.001751175, 0.001751178, 0.001751174, 
    0.001751173, 0.001751175, 0.001751165, 0.001751168, 0.001751165, 
    0.001751167, 0.001751213, 0.00175121, 0.001751212, 0.001751209, 
    0.001751211, 0.001751204, 0.001751202, 0.001751191, 0.001751196, 
    0.001751189, 0.001751195, 0.001751194, 0.001751189, 0.001751195, 
    0.001751182, 0.001751191, 0.001751175, 0.001751183, 0.001751174, 
    0.001751176, 0.001751173, 0.00175117, 0.001751167, 0.001751162, 
    0.001751163, 0.001751158, 0.001751207, 0.001751204, 0.001751204, 
    0.001751201, 0.001751199, 0.001751194, 0.001751186, 0.001751189, 
    0.001751184, 0.001751183, 0.001751191, 0.001751186, 0.001751202, 
    0.001751199, 0.001751201, 0.001751207, 0.001751188, 0.001751198, 
    0.001751181, 0.001751186, 0.001751171, 0.001751178, 0.001751164, 
    0.001751158, 0.001751152, 0.001751145, 0.001751202, 0.001751204, 
    0.001751201, 0.001751196, 0.001751191, 0.001751185, 0.001751185, 
    0.001751184, 0.001751181, 0.001751178, 0.001751183, 0.001751177, 
    0.001751199, 0.001751188, 0.001751205, 0.0017512, 0.001751196, 
    0.001751198, 0.001751189, 0.001751187, 0.00175118, 0.001751184, 
    0.001751159, 0.00175117, 0.00175114, 0.001751148, 0.001751205, 
    0.001751202, 0.001751193, 0.001751198, 0.001751185, 0.001751182, 
    0.001751179, 0.001751176, 0.001751176, 0.001751174, 0.001751177, 
    0.001751174, 0.001751185, 0.00175118, 0.001751194, 0.001751191, 
    0.001751192, 0.001751194, 0.001751189, 0.001751183, 0.001751183, 
    0.001751181, 0.001751176, 0.001751185, 0.001751158, 0.001751174, 
    0.001751199, 0.001751194, 0.001751194, 0.001751196, 0.001751182, 
    0.001751187, 0.001751174, 0.001751177, 0.001751172, 0.001751174, 
    0.001751175, 0.001751179, 0.001751181, 0.001751187, 0.001751192, 
    0.001751195, 0.001751194, 0.00175119, 0.001751183, 0.001751176, 
    0.001751177, 0.001751172, 0.001751186, 0.00175118, 0.001751182, 
    0.001751176, 0.001751189, 0.001751178, 0.001751192, 0.001751191, 
    0.001751187, 0.00175118, 0.001751178, 0.001751176, 0.001751177, 
    0.001751183, 0.001751183, 0.001751187, 0.001751188, 0.001751191, 
    0.001751193, 0.001751191, 0.001751189, 0.001751183, 0.001751177, 
    0.00175117, 0.001751169, 0.001751162, 0.001751167, 0.001751158, 
    0.001751166, 0.001751151, 0.001751178, 0.001751166, 0.001751187, 
    0.001751185, 0.001751181, 0.001751171, 0.001751176, 0.001751171, 
    0.001751183, 0.00175119, 0.001751192, 0.001751195, 0.001751192, 
    0.001751192, 0.001751189, 0.00175119, 0.001751182, 0.001751186, 
    0.001751175, 0.001751171, 0.001751159, 0.001751152, 0.001751144, 
    0.001751141, 0.00175114, 0.001751139,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N =
  9.733135e-07, 9.733097e-07, 9.733105e-07, 9.733075e-07, 9.733092e-07, 
    9.733071e-07, 9.733127e-07, 9.733096e-07, 9.733116e-07, 9.733131e-07, 
    9.733016e-07, 9.733074e-07, 9.732956e-07, 9.732993e-07, 9.732901e-07, 
    9.732962e-07, 9.732888e-07, 9.732903e-07, 9.732861e-07, 9.732872e-07, 
    9.732819e-07, 9.732855e-07, 9.73279e-07, 9.732827e-07, 9.732821e-07, 
    9.732856e-07, 9.733062e-07, 9.733022e-07, 9.733064e-07, 9.733059e-07, 
    9.733061e-07, 9.733091e-07, 9.733106e-07, 9.733138e-07, 9.733133e-07, 
    9.733109e-07, 9.733055e-07, 9.733074e-07, 9.733028e-07, 9.733029e-07, 
    9.732979e-07, 9.733002e-07, 9.732918e-07, 9.732942e-07, 9.732872e-07, 
    9.732889e-07, 9.732872e-07, 9.732878e-07, 9.732872e-07, 9.732898e-07, 
    9.732887e-07, 9.73291e-07, 9.732997e-07, 9.732972e-07, 9.733049e-07, 
    9.733095e-07, 9.733126e-07, 9.733147e-07, 9.733145e-07, 9.733139e-07, 
    9.733109e-07, 9.73308e-07, 9.733059e-07, 9.733044e-07, 9.733029e-07, 
    9.732987e-07, 9.732963e-07, 9.732912e-07, 9.732921e-07, 9.732906e-07, 
    9.732892e-07, 9.732867e-07, 9.73287e-07, 9.73286e-07, 9.732906e-07, 
    9.732875e-07, 9.732927e-07, 9.732913e-07, 9.733026e-07, 9.733069e-07, 
    9.733087e-07, 9.733103e-07, 9.733143e-07, 9.733116e-07, 9.733126e-07, 
    9.733101e-07, 9.733085e-07, 9.733093e-07, 9.733044e-07, 9.733062e-07, 
    9.732962e-07, 9.733005e-07, 9.732893e-07, 9.73292e-07, 9.732886e-07, 
    9.732903e-07, 9.732875e-07, 9.732901e-07, 9.732855e-07, 9.732845e-07, 
    9.732852e-07, 9.732826e-07, 9.732902e-07, 9.732872e-07, 9.733093e-07, 
    9.733092e-07, 9.733086e-07, 9.733112e-07, 9.733113e-07, 9.733138e-07, 
    9.733117e-07, 9.733108e-07, 9.733084e-07, 9.73307e-07, 9.733056e-07, 
    9.733028e-07, 9.732995e-07, 9.732951e-07, 9.732918e-07, 9.732896e-07, 
    9.73291e-07, 9.732898e-07, 9.732911e-07, 9.732918e-07, 9.732848e-07, 
    9.732887e-07, 9.73283e-07, 9.732832e-07, 9.732859e-07, 9.732832e-07, 
    9.733091e-07, 9.733099e-07, 9.733125e-07, 9.733104e-07, 9.733141e-07, 
    9.73312e-07, 9.733109e-07, 9.733062e-07, 9.733052e-07, 9.733043e-07, 
    9.733025e-07, 9.733001e-07, 9.73296e-07, 9.732923e-07, 9.73289e-07, 
    9.732893e-07, 9.732892e-07, 9.732885e-07, 9.732903e-07, 9.732881e-07, 
    9.732878e-07, 9.732887e-07, 9.732834e-07, 9.732848e-07, 9.732832e-07, 
    9.732843e-07, 9.733096e-07, 9.733084e-07, 9.733089e-07, 9.733077e-07, 
    9.733086e-07, 9.733046e-07, 9.733034e-07, 9.732978e-07, 9.733001e-07, 
    9.732964e-07, 9.732997e-07, 9.732992e-07, 9.732963e-07, 9.732996e-07, 
    9.732926e-07, 9.732973e-07, 9.732885e-07, 9.732933e-07, 9.732881e-07, 
    9.73289e-07, 9.732876e-07, 9.732862e-07, 9.732845e-07, 9.732813e-07, 
    9.73282e-07, 9.732794e-07, 9.733064e-07, 9.733049e-07, 9.73305e-07, 
    9.733033e-07, 9.73302e-07, 9.732993e-07, 9.732948e-07, 9.732966e-07, 
    9.732935e-07, 9.732929e-07, 9.732975e-07, 9.732947e-07, 9.733037e-07, 
    9.733022e-07, 9.733031e-07, 9.733063e-07, 9.732962e-07, 9.733013e-07, 
    9.732918e-07, 9.732946e-07, 9.732863e-07, 9.732904e-07, 9.732825e-07, 
    9.73279e-07, 9.732757e-07, 9.73272e-07, 9.733039e-07, 9.733051e-07, 
    9.73303e-07, 9.733003e-07, 9.732978e-07, 9.732944e-07, 9.73294e-07, 
    9.732935e-07, 9.732918e-07, 9.732904e-07, 9.732933e-07, 9.732901e-07, 
    9.733019e-07, 9.732958e-07, 9.733054e-07, 9.733026e-07, 9.733005e-07, 
    9.733013e-07, 9.732968e-07, 9.732956e-07, 9.732912e-07, 9.732935e-07, 
    9.732798e-07, 9.732859e-07, 9.732692e-07, 9.732738e-07, 9.733054e-07, 
    9.733039e-07, 9.732987e-07, 9.733012e-07, 9.732942e-07, 9.732925e-07, 
    9.732911e-07, 9.732893e-07, 9.73289e-07, 9.73288e-07, 9.732897e-07, 
    9.73288e-07, 9.732944e-07, 9.732915e-07, 9.732994e-07, 9.732975e-07, 
    9.732984e-07, 9.732993e-07, 9.732963e-07, 9.732931e-07, 9.732931e-07, 
    9.732921e-07, 9.732893e-07, 9.732942e-07, 9.73279e-07, 9.732884e-07, 
    9.733023e-07, 9.732994e-07, 9.732991e-07, 9.733002e-07, 9.732926e-07, 
    9.732953e-07, 9.73288e-07, 9.7329e-07, 9.732868e-07, 9.732884e-07, 
    9.732886e-07, 9.732906e-07, 9.73292e-07, 9.732952e-07, 9.732979e-07, 
    9.733e-07, 9.732995e-07, 9.732972e-07, 9.73293e-07, 9.73289e-07, 
    9.732898e-07, 9.73287e-07, 9.732947e-07, 9.732914e-07, 9.732927e-07, 
    9.732895e-07, 9.732966e-07, 9.732905e-07, 9.732981e-07, 9.732975e-07, 
    9.732954e-07, 9.732912e-07, 9.732903e-07, 9.732894e-07, 9.7329e-07, 
    9.732929e-07, 9.732934e-07, 9.732954e-07, 9.73296e-07, 9.732976e-07, 
    9.732989e-07, 9.732977e-07, 9.732964e-07, 9.732929e-07, 9.732896e-07, 
    9.732861e-07, 9.732853e-07, 9.732812e-07, 9.732845e-07, 9.73279e-07, 
    9.732837e-07, 9.732756e-07, 9.732902e-07, 9.732838e-07, 9.732953e-07, 
    9.73294e-07, 9.732918e-07, 9.732867e-07, 9.732895e-07, 9.732862e-07, 
    9.732934e-07, 9.732971e-07, 9.73298e-07, 9.732998e-07, 9.73298e-07, 
    9.732981e-07, 9.732964e-07, 9.73297e-07, 9.732928e-07, 9.732951e-07, 
    9.732886e-07, 9.732862e-07, 9.732796e-07, 9.732756e-07, 9.732714e-07, 
    9.732697e-07, 9.732692e-07, 9.732689e-07 ;

 LITR1N_TNDNCY_VERT_TRANS =
  1.960724e-25, 4.901811e-26, 4.313593e-25, -6.862535e-26, 9.313441e-26, 
    -4.215557e-25, -1.960724e-26, 4.117521e-25, 3.725376e-25, 7.695843e-25, 
    3.431268e-25, 7.352717e-26, -1.176435e-25, -2.646978e-25, -3.62734e-25, 
    -9.999695e-25, 1.56858e-25, 1.323489e-25, -1.960724e-26, 1.960724e-25, 
    1.862688e-25, 2.548942e-25, -6.862535e-25, 2.352869e-25, -4.509666e-25, 
    6.274318e-25, 6.764499e-25, 2.401887e-25, -3.823413e-25, 3.529304e-25, 
    1.372507e-25, 1.666616e-25, 9.705585e-25, -2.745014e-25, 2.941087e-25, 
    1.078398e-25, 8.333079e-26, 9.656568e-25, 4.019485e-25, 6.862535e-25, 
    1.078398e-25, 4.803775e-25, 4.313593e-25, 9.803622e-26, 7.352717e-26, 
    6.122413e-41, -6.274318e-25, 2.058761e-25, 5.391992e-26, -3.137159e-25, 
    -1.56858e-25, -4.460648e-25, 1.176435e-25, 3.725376e-25, 2.352869e-25, 
    -4.901811e-27, 4.460648e-25, 5.588064e-25, 3.529304e-25, -1.764652e-25, 
    8.82326e-26, 3.921449e-25, 3.431268e-25, 2.156797e-25, -4.215557e-25, 
    3.725376e-25, 2.107779e-25, 1.274471e-25, -4.019485e-25, 1.81367e-25, 
    5.637083e-25, 1.323489e-25, 6.372354e-25, -1.196042e-24, -1.617598e-25, 
    4.901811e-26, -3.921449e-26, 3.039123e-25, -2.450906e-25, -3.431268e-26, 
    -1.56858e-25, 5.490028e-25, 9.803622e-27, -3.284213e-25, 9.313441e-26, 
    7.352717e-26, 4.803775e-25, -2.695996e-25, 5.784137e-25, 5.882173e-25, 0, 
    -3.186177e-25, 4.509666e-25, -2.254833e-25, -4.117521e-25, 5.19592e-25, 
    1.764652e-25, 1.127417e-25, -1.764652e-25, -8.82326e-26, 6.372354e-26, 
    -1.470543e-25, -4.509666e-25, -8.82326e-26, 2.254833e-25, -1.274471e-25, 
    9.705585e-25, -5.98021e-25, -2.009742e-25, 2.401887e-25, 3.823413e-25, 
    7.156644e-25, 8.725224e-25, 1.666616e-25, -8.235043e-25, -6.372354e-26, 
    -1.519561e-25, 3.823413e-25, 5.588064e-25, -1.176435e-25, 3.872431e-25, 
    4.901811e-25, 1.960724e-26, -2.156797e-25, 9.950677e-25, -2.941087e-25, 
    -2.352869e-25, 3.676358e-25, -2.107779e-25, 4.607703e-25, 4.852793e-25, 
    4.901811e-25, 7.205662e-25, -3.039123e-25, -4.019485e-25, 4.901811e-25, 
    7.842898e-25, 6.764499e-25, 1.200944e-24, 6.862535e-26, 1.666616e-25, 
    -1.56858e-25, 1.323489e-25, 2.450906e-25, -1.048988e-24, 2.59796e-25, 
    -4.117521e-25, 4.313593e-25, 5.882173e-26, 5.784137e-25, 2.892069e-25, 
    -4.705739e-25, 4.41163e-25, 1.715634e-25, 5.686101e-25, 1.715634e-25, 
    -2.646978e-25, -3.921449e-26, 2.794032e-25, 4.705739e-25, 4.509666e-25, 
    -3.578322e-25, 3.186177e-25, 2.548942e-25, 4.901811e-25, 2.548942e-25, 
    2.941087e-25, -2.941087e-26, 6.568427e-25, -1.019577e-24, -1.02938e-25, 
    -2.794032e-25, 5.882173e-26, -3.284213e-25, 4.754757e-25, -9.411477e-25, 
    2.745014e-25, 1.274471e-25, 3.431268e-25, 6.372354e-25, -2.352869e-25, 
    -4.41163e-25, -3.431268e-26, -2.941087e-26, -9.803622e-27, -5.293956e-25, 
    2.941087e-26, 1.323489e-25, 4.166539e-25, -4.068503e-25, -5.391992e-26, 
    -6.911554e-25, 4.313593e-25, 6.274318e-25, -5.342974e-25, -6.862535e-26, 
    1.225453e-25, -6.862535e-26, 8.725224e-25, 3.725376e-25, 3.62734e-25, 
    -2.794032e-25, 1.56858e-25, -2.450906e-25, 3.186177e-25, -6.176282e-25, 
    4.313593e-25, -5.588064e-25, 7.891916e-25, -2.107779e-25, 9.803622e-27, 
    -3.62734e-25, 3.431268e-25, -1.764652e-25, 2.548942e-25, 1.176435e-25, 
    -9.803622e-26, -1.960724e-26, 1.715634e-25, 2.548942e-25, -8.82326e-26, 
    2.941087e-26, 6.617445e-25, 3.235195e-25, -8.82326e-26, 9.803622e-26, 
    -8.82326e-26, -4.607703e-25, 4.852793e-25, 6.372354e-25, 7.450753e-25, 
    3.872431e-25, 5.146902e-25, -1.764652e-25, 7.891916e-25, 2.59796e-25, 
    -2.254833e-25, 2.254833e-25, 1.176435e-25, -7.352717e-25, 3.529304e-25, 
    8.03897e-25, 4.999847e-25, 4.754757e-25, 5.882173e-26, -6.122413e-41, 
    9.85264e-25, 3.921449e-26, -6.862535e-26, 4.999847e-25, 6.274318e-25, 
    4.901811e-25, 7.842898e-26, 2.990105e-25, -7.25468e-25, 8.82326e-25, 
    5.293956e-25, 4.068503e-25, -6.372354e-25, -5.391992e-26, -1.470543e-26, 
    6.960572e-25, 3.284213e-25, -3.725376e-25, 4.901811e-25, -6.568427e-25, 
    -3.137159e-25, -9.705585e-25, -8.03897e-25, -1.960724e-26, -4.607703e-25, 
    -3.431268e-25, 1.56858e-25, -1.078398e-25, -5.490028e-25, 3.62734e-25, 
    -3.921449e-26, -3.921449e-26, -2.646978e-25, 1.323489e-25, 6.960572e-25, 
    -1.323489e-25, 9.411477e-25, -4.901811e-26, -3.039123e-25, -1.862688e-25, 
    8.03897e-25, 0, 2.646978e-25, 4.215557e-25, 8.137007e-25, -3.921449e-26, 
    4.999847e-25, -3.333231e-25, 5.686101e-25, 2.156797e-25, -4.313593e-25, 
    1.02938e-24, 9.803622e-25, 2.794032e-25, 5.293956e-25, -6.862535e-26, 
    3.921449e-26, 8.725224e-25, 4.313593e-25, 2.499924e-25, -2.156797e-25, 
    6.862535e-25, -2.254833e-25, -4.215557e-25, -5.391992e-25, 2.156797e-25, 
    1.127417e-24, -5.784137e-25, -5.391992e-25, 1.81367e-25, -4.313593e-25, 
    5.490028e-25, 2.450906e-25, -3.921449e-25, 1.421525e-25, 5.882173e-26, 
    -1.617598e-25, 4.705739e-25, 1.323489e-25, 5.097883e-25, 3.578322e-25, 
    2.156797e-25, -2.303851e-25, 1.56858e-25, 7.842898e-26, -5.98021e-25, 
    3.284213e-25, 4.803775e-25, 3.529304e-25, -4.509666e-25, 9.754604e-25, 
    -7.79388e-25,
  9.436976e-32, 9.436938e-32, 9.436946e-32, 9.436915e-32, 9.436932e-32, 
    9.436912e-32, 9.436969e-32, 9.436937e-32, 9.436957e-32, 9.436973e-32, 
    9.436856e-32, 9.436914e-32, 9.436796e-32, 9.436833e-32, 9.436741e-32, 
    9.436802e-32, 9.436728e-32, 9.436742e-32, 9.4367e-32, 9.436712e-32, 
    9.436658e-32, 9.436695e-32, 9.43663e-32, 9.436666e-32, 9.436661e-32, 
    9.436696e-32, 9.436902e-32, 9.436863e-32, 9.436905e-32, 9.436899e-32, 
    9.436902e-32, 9.436932e-32, 9.436947e-32, 9.436979e-32, 9.436973e-32, 
    9.43695e-32, 9.436896e-32, 9.436914e-32, 9.436869e-32, 9.43687e-32, 
    9.436819e-32, 9.436842e-32, 9.436758e-32, 9.436782e-32, 9.436712e-32, 
    9.436729e-32, 9.436712e-32, 9.436718e-32, 9.436712e-32, 9.436738e-32, 
    9.436727e-32, 9.43675e-32, 9.436838e-32, 9.436812e-32, 9.436889e-32, 
    9.436936e-32, 9.436967e-32, 9.436989e-32, 9.436986e-32, 9.43698e-32, 
    9.43695e-32, 9.436921e-32, 9.436899e-32, 9.436885e-32, 9.43687e-32, 
    9.436827e-32, 9.436804e-32, 9.436752e-32, 9.436762e-32, 9.436746e-32, 
    9.436731e-32, 9.436706e-32, 9.43671e-32, 9.436699e-32, 9.436746e-32, 
    9.436715e-32, 9.436767e-32, 9.436753e-32, 9.436866e-32, 9.43691e-32, 
    9.436928e-32, 9.436944e-32, 9.436983e-32, 9.436956e-32, 9.436967e-32, 
    9.436942e-32, 9.436926e-32, 9.436933e-32, 9.436884e-32, 9.436903e-32, 
    9.436802e-32, 9.436846e-32, 9.436733e-32, 9.43676e-32, 9.436726e-32, 
    9.436743e-32, 9.436714e-32, 9.436741e-32, 9.436695e-32, 9.436685e-32, 
    9.436692e-32, 9.436665e-32, 9.436742e-32, 9.436712e-32, 9.436934e-32, 
    9.436932e-32, 9.436926e-32, 9.436953e-32, 9.436954e-32, 9.436979e-32, 
    9.436957e-32, 9.436948e-32, 9.436924e-32, 9.43691e-32, 9.436897e-32, 
    9.436868e-32, 9.436836e-32, 9.43679e-32, 9.436758e-32, 9.436736e-32, 
    9.436749e-32, 9.436738e-32, 9.436751e-32, 9.436757e-32, 9.436689e-32, 
    9.436727e-32, 9.436669e-32, 9.436672e-32, 9.436699e-32, 9.436672e-32, 
    9.436932e-32, 9.436939e-32, 9.436965e-32, 9.436944e-32, 9.436981e-32, 
    9.436961e-32, 9.436949e-32, 9.436903e-32, 9.436893e-32, 9.436883e-32, 
    9.436865e-32, 9.436841e-32, 9.436799e-32, 9.436763e-32, 9.43673e-32, 
    9.436732e-32, 9.436732e-32, 9.436724e-32, 9.436743e-32, 9.436721e-32, 
    9.436718e-32, 9.436727e-32, 9.436673e-32, 9.436688e-32, 9.436672e-32, 
    9.436683e-32, 9.436936e-32, 9.436924e-32, 9.436931e-32, 9.436918e-32, 
    9.436927e-32, 9.436887e-32, 9.436875e-32, 9.436819e-32, 9.436842e-32, 
    9.436805e-32, 9.436838e-32, 9.436832e-32, 9.436803e-32, 9.436836e-32, 
    9.436765e-32, 9.436813e-32, 9.436724e-32, 9.436772e-32, 9.436721e-32, 
    9.436731e-32, 9.436715e-32, 9.436701e-32, 9.436684e-32, 9.436652e-32, 
    9.436659e-32, 9.436633e-32, 9.436905e-32, 9.436889e-32, 9.43689e-32, 
    9.436873e-32, 9.43686e-32, 9.436833e-32, 9.436789e-32, 9.436806e-32, 
    9.436775e-32, 9.436769e-32, 9.436815e-32, 9.436787e-32, 9.436878e-32, 
    9.436863e-32, 9.436872e-32, 9.436904e-32, 9.436802e-32, 9.436854e-32, 
    9.436758e-32, 9.436786e-32, 9.436703e-32, 9.436744e-32, 9.436664e-32, 
    9.436629e-32, 9.436597e-32, 9.436559e-32, 9.43688e-32, 9.436891e-32, 
    9.436871e-32, 9.436843e-32, 9.436818e-32, 9.436784e-32, 9.43678e-32, 
    9.436774e-32, 9.436758e-32, 9.436744e-32, 9.436772e-32, 9.436741e-32, 
    9.43686e-32, 9.436798e-32, 9.436895e-32, 9.436866e-32, 9.436845e-32, 
    9.436854e-32, 9.436808e-32, 9.436796e-32, 9.436752e-32, 9.436775e-32, 
    9.436638e-32, 9.436698e-32, 9.43653e-32, 9.436577e-32, 9.436895e-32, 
    9.43688e-32, 9.436828e-32, 9.436853e-32, 9.436782e-32, 9.436765e-32, 
    9.436751e-32, 9.436732e-32, 9.436731e-32, 9.436719e-32, 9.436737e-32, 
    9.436721e-32, 9.436784e-32, 9.436756e-32, 9.436834e-32, 9.436815e-32, 
    9.436823e-32, 9.436833e-32, 9.436803e-32, 9.436772e-32, 9.436771e-32, 
    9.436761e-32, 9.436732e-32, 9.436782e-32, 9.43663e-32, 9.436723e-32, 
    9.436863e-32, 9.436835e-32, 9.43683e-32, 9.436842e-32, 9.436766e-32, 
    9.436793e-32, 9.43672e-32, 9.43674e-32, 9.436707e-32, 9.436723e-32, 
    9.436726e-32, 9.436746e-32, 9.436759e-32, 9.436792e-32, 9.436819e-32, 
    9.43684e-32, 9.436835e-32, 9.436812e-32, 9.43677e-32, 9.43673e-32, 
    9.436739e-32, 9.436709e-32, 9.436787e-32, 9.436755e-32, 9.436767e-32, 
    9.436735e-32, 9.436806e-32, 9.436745e-32, 9.436822e-32, 9.436815e-32, 
    9.436794e-32, 9.436752e-32, 9.436743e-32, 9.436733e-32, 9.436739e-32, 
    9.436769e-32, 9.436773e-32, 9.436795e-32, 9.4368e-32, 9.436816e-32, 
    9.43683e-32, 9.436818e-32, 9.436805e-32, 9.436769e-32, 9.436736e-32, 
    9.436701e-32, 9.436692e-32, 9.436651e-32, 9.436685e-32, 9.436629e-32, 
    9.436676e-32, 9.436595e-32, 9.436742e-32, 9.436678e-32, 9.436793e-32, 
    9.43678e-32, 9.436758e-32, 9.436707e-32, 9.436735e-32, 9.436702e-32, 
    9.436774e-32, 9.436811e-32, 9.436821e-32, 9.436839e-32, 9.43682e-32, 
    9.436822e-32, 9.436805e-32, 9.43681e-32, 9.436768e-32, 9.43679e-32, 
    9.436726e-32, 9.436702e-32, 9.436636e-32, 9.436595e-32, 9.436554e-32, 
    9.436535e-32, 9.43653e-32, 9.436528e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1N_TO_SOIL1N =
  4.500506e-14, 4.512833e-14, 4.510439e-14, 4.520373e-14, 4.514865e-14, 
    4.521368e-14, 4.503008e-14, 4.513321e-14, 4.506739e-14, 4.501619e-14, 
    4.53963e-14, 4.520817e-14, 4.559166e-14, 4.547183e-14, 4.577274e-14, 
    4.557299e-14, 4.581298e-14, 4.576702e-14, 4.590542e-14, 4.586579e-14, 
    4.604257e-14, 4.592371e-14, 4.613419e-14, 4.601422e-14, 4.603298e-14, 
    4.591978e-14, 4.524609e-14, 4.537287e-14, 4.523857e-14, 4.525665e-14, 
    4.524855e-14, 4.514977e-14, 4.509994e-14, 4.499567e-14, 4.501461e-14, 
    4.509121e-14, 4.526479e-14, 4.520591e-14, 4.535433e-14, 4.535098e-14, 
    4.551602e-14, 4.544163e-14, 4.571879e-14, 4.564008e-14, 4.586745e-14, 
    4.581029e-14, 4.586475e-14, 4.584825e-14, 4.586497e-14, 4.578114e-14, 
    4.581706e-14, 4.574329e-14, 4.545556e-14, 4.554016e-14, 4.528767e-14, 
    4.513558e-14, 4.50346e-14, 4.496287e-14, 4.497301e-14, 4.499233e-14, 
    4.509166e-14, 4.518503e-14, 4.525613e-14, 4.530367e-14, 4.53505e-14, 
    4.549206e-14, 4.556703e-14, 4.573467e-14, 4.570447e-14, 4.575566e-14, 
    4.580461e-14, 4.588669e-14, 4.587319e-14, 4.590933e-14, 4.575434e-14, 
    4.585735e-14, 4.568726e-14, 4.573379e-14, 4.536308e-14, 4.522181e-14, 
    4.516159e-14, 4.510898e-14, 4.49808e-14, 4.506933e-14, 4.503443e-14, 
    4.511746e-14, 4.517018e-14, 4.514412e-14, 4.530497e-14, 4.524245e-14, 
    4.557147e-14, 4.542983e-14, 4.57989e-14, 4.571068e-14, 4.582004e-14, 
    4.576425e-14, 4.585982e-14, 4.577381e-14, 4.592279e-14, 4.595519e-14, 
    4.593305e-14, 4.601814e-14, 4.576904e-14, 4.586474e-14, 4.514338e-14, 
    4.514763e-14, 4.516745e-14, 4.508031e-14, 4.507499e-14, 4.499514e-14, 
    4.50662e-14, 4.509645e-14, 4.517325e-14, 4.521863e-14, 4.526177e-14, 
    4.535658e-14, 4.546238e-14, 4.561023e-14, 4.571639e-14, 4.57875e-14, 
    4.574391e-14, 4.57824e-14, 4.573937e-14, 4.571921e-14, 4.594304e-14, 
    4.581738e-14, 4.600591e-14, 4.599549e-14, 4.591018e-14, 4.599666e-14, 
    4.515062e-14, 4.512615e-14, 4.504113e-14, 4.510767e-14, 4.498644e-14, 
    4.505429e-14, 4.509328e-14, 4.524372e-14, 4.527679e-14, 4.53074e-14, 
    4.536788e-14, 4.544544e-14, 4.558139e-14, 4.569961e-14, 4.580746e-14, 
    4.579956e-14, 4.580234e-14, 4.582641e-14, 4.576676e-14, 4.58362e-14, 
    4.584784e-14, 4.581739e-14, 4.599409e-14, 4.594363e-14, 4.599527e-14, 
    4.596242e-14, 4.513411e-14, 4.517528e-14, 4.515303e-14, 4.519485e-14, 
    4.516538e-14, 4.529636e-14, 4.533561e-14, 4.551917e-14, 4.54439e-14, 
    4.556372e-14, 4.545609e-14, 4.547516e-14, 4.556757e-14, 4.546192e-14, 
    4.569306e-14, 4.553634e-14, 4.582735e-14, 4.567092e-14, 4.583714e-14, 
    4.580699e-14, 4.585692e-14, 4.59016e-14, 4.595782e-14, 4.606144e-14, 
    4.603746e-14, 4.61241e-14, 4.523664e-14, 4.528999e-14, 4.528532e-14, 
    4.534116e-14, 4.538243e-14, 4.547188e-14, 4.56152e-14, 4.556133e-14, 
    4.566025e-14, 4.568008e-14, 4.552982e-14, 4.562207e-14, 4.532571e-14, 
    4.53736e-14, 4.534511e-14, 4.524084e-14, 4.557371e-14, 4.540295e-14, 
    4.571814e-14, 4.562575e-14, 4.589522e-14, 4.576125e-14, 4.602425e-14, 
    4.613645e-14, 4.62421e-14, 4.63653e-14, 4.531913e-14, 4.528289e-14, 
    4.53478e-14, 4.543752e-14, 4.552079e-14, 4.563139e-14, 4.564271e-14, 
    4.566341e-14, 4.571705e-14, 4.576212e-14, 4.566993e-14, 4.577342e-14, 
    4.538465e-14, 4.558853e-14, 4.526916e-14, 4.536536e-14, 4.543224e-14, 
    4.540293e-14, 4.555518e-14, 4.559103e-14, 4.573661e-14, 4.566139e-14, 
    4.610874e-14, 4.591099e-14, 4.645913e-14, 4.630616e-14, 4.527021e-14, 
    4.531902e-14, 4.548871e-14, 4.5408e-14, 4.563878e-14, 4.569552e-14, 
    4.574166e-14, 4.580056e-14, 4.580694e-14, 4.584183e-14, 4.578465e-14, 
    4.583958e-14, 4.563162e-14, 4.57246e-14, 4.546936e-14, 4.553151e-14, 
    4.550293e-14, 4.547156e-14, 4.556836e-14, 4.567138e-14, 4.567362e-14, 
    4.570663e-14, 4.579952e-14, 4.563972e-14, 4.613416e-14, 4.582893e-14, 
    4.537222e-14, 4.546608e-14, 4.547954e-14, 4.544318e-14, 4.568983e-14, 
    4.56005e-14, 4.584099e-14, 4.577604e-14, 4.588245e-14, 4.582958e-14, 
    4.58218e-14, 4.575387e-14, 4.571155e-14, 4.560459e-14, 4.551752e-14, 
    4.544846e-14, 4.546452e-14, 4.554037e-14, 4.567768e-14, 4.58075e-14, 
    4.577906e-14, 4.587437e-14, 4.562206e-14, 4.572789e-14, 4.568698e-14, 
    4.579363e-14, 4.555989e-14, 4.575882e-14, 4.550898e-14, 4.553091e-14, 
    4.559873e-14, 4.573503e-14, 4.576524e-14, 4.57974e-14, 4.577756e-14, 
    4.568118e-14, 4.56654e-14, 4.559709e-14, 4.55782e-14, 4.552614e-14, 
    4.5483e-14, 4.552241e-14, 4.556377e-14, 4.568124e-14, 4.578699e-14, 
    4.590222e-14, 4.593043e-14, 4.60648e-14, 4.595536e-14, 4.613584e-14, 
    4.598232e-14, 4.624802e-14, 4.57704e-14, 4.59779e-14, 4.560183e-14, 
    4.56424e-14, 4.571571e-14, 4.58838e-14, 4.579313e-14, 4.589919e-14, 
    4.566479e-14, 4.554297e-14, 4.551149e-14, 4.545265e-14, 4.551284e-14, 
    4.550794e-14, 4.556551e-14, 4.554702e-14, 4.568514e-14, 4.561096e-14, 
    4.582159e-14, 4.589836e-14, 4.6115e-14, 4.624761e-14, 4.638253e-14, 
    4.644203e-14, 4.646014e-14, 4.64677e-14 ;

 LITR1N_vr =
  5.557721e-05, 5.557699e-05, 5.557703e-05, 5.557686e-05, 5.557696e-05, 
    5.557685e-05, 5.557716e-05, 5.557698e-05, 5.55771e-05, 5.557719e-05, 
    5.557653e-05, 5.557685e-05, 5.557619e-05, 5.557639e-05, 5.557587e-05, 
    5.557622e-05, 5.55758e-05, 5.557588e-05, 5.557564e-05, 5.557571e-05, 
    5.55754e-05, 5.557561e-05, 5.557524e-05, 5.557545e-05, 5.557542e-05, 
    5.557561e-05, 5.557679e-05, 5.557657e-05, 5.55768e-05, 5.557677e-05, 
    5.557678e-05, 5.557695e-05, 5.557704e-05, 5.557722e-05, 5.557719e-05, 
    5.557706e-05, 5.557675e-05, 5.557686e-05, 5.55766e-05, 5.557661e-05, 
    5.557632e-05, 5.557645e-05, 5.557597e-05, 5.55761e-05, 5.55757e-05, 
    5.557581e-05, 5.557571e-05, 5.557574e-05, 5.557571e-05, 5.557586e-05, 
    5.557579e-05, 5.557592e-05, 5.557642e-05, 5.557627e-05, 5.557671e-05, 
    5.557698e-05, 5.557715e-05, 5.557728e-05, 5.557726e-05, 5.557723e-05, 
    5.557706e-05, 5.557689e-05, 5.557677e-05, 5.557669e-05, 5.557661e-05, 
    5.557636e-05, 5.557623e-05, 5.557594e-05, 5.557599e-05, 5.55759e-05, 
    5.557582e-05, 5.557567e-05, 5.55757e-05, 5.557563e-05, 5.55759e-05, 
    5.557572e-05, 5.557602e-05, 5.557594e-05, 5.557658e-05, 5.557683e-05, 
    5.557693e-05, 5.557703e-05, 5.557725e-05, 5.55771e-05, 5.557715e-05, 
    5.557701e-05, 5.557692e-05, 5.557697e-05, 5.557669e-05, 5.557679e-05, 
    5.557622e-05, 5.557647e-05, 5.557582e-05, 5.557598e-05, 5.557579e-05, 
    5.557589e-05, 5.557572e-05, 5.557587e-05, 5.557561e-05, 5.557555e-05, 
    5.557559e-05, 5.557544e-05, 5.557588e-05, 5.557571e-05, 5.557697e-05, 
    5.557696e-05, 5.557693e-05, 5.557707e-05, 5.557709e-05, 5.557722e-05, 
    5.55771e-05, 5.557705e-05, 5.557691e-05, 5.557683e-05, 5.557676e-05, 
    5.557659e-05, 5.557641e-05, 5.557615e-05, 5.557597e-05, 5.557585e-05, 
    5.557592e-05, 5.557585e-05, 5.557593e-05, 5.557596e-05, 5.557557e-05, 
    5.557579e-05, 5.557546e-05, 5.557548e-05, 5.557563e-05, 5.557548e-05, 
    5.557695e-05, 5.557699e-05, 5.557714e-05, 5.557703e-05, 5.557724e-05, 
    5.557712e-05, 5.557705e-05, 5.557679e-05, 5.557673e-05, 5.557668e-05, 
    5.557658e-05, 5.557644e-05, 5.55762e-05, 5.5576e-05, 5.557581e-05, 
    5.557582e-05, 5.557582e-05, 5.557578e-05, 5.557588e-05, 5.557576e-05, 
    5.557574e-05, 5.557579e-05, 5.557549e-05, 5.557557e-05, 5.557548e-05, 
    5.557554e-05, 5.557698e-05, 5.557691e-05, 5.557695e-05, 5.557688e-05, 
    5.557693e-05, 5.55767e-05, 5.557663e-05, 5.557631e-05, 5.557644e-05, 
    5.557623e-05, 5.557642e-05, 5.557639e-05, 5.557623e-05, 5.557641e-05, 
    5.557601e-05, 5.557628e-05, 5.557578e-05, 5.557605e-05, 5.557576e-05, 
    5.557581e-05, 5.557572e-05, 5.557565e-05, 5.557555e-05, 5.557537e-05, 
    5.557541e-05, 5.557526e-05, 5.557681e-05, 5.557671e-05, 5.557672e-05, 
    5.557662e-05, 5.557655e-05, 5.557639e-05, 5.557614e-05, 5.557624e-05, 
    5.557607e-05, 5.557603e-05, 5.557629e-05, 5.557613e-05, 5.557665e-05, 
    5.557657e-05, 5.557662e-05, 5.55768e-05, 5.557622e-05, 5.557651e-05, 
    5.557597e-05, 5.557613e-05, 5.557566e-05, 5.557589e-05, 5.557543e-05, 
    5.557524e-05, 5.557505e-05, 5.557484e-05, 5.557666e-05, 5.557672e-05, 
    5.557661e-05, 5.557645e-05, 5.557631e-05, 5.557612e-05, 5.55761e-05, 
    5.557606e-05, 5.557597e-05, 5.557589e-05, 5.557605e-05, 5.557587e-05, 
    5.557655e-05, 5.557619e-05, 5.557675e-05, 5.557658e-05, 5.557646e-05, 
    5.557651e-05, 5.557625e-05, 5.557619e-05, 5.557593e-05, 5.557606e-05, 
    5.557528e-05, 5.557563e-05, 5.557467e-05, 5.557494e-05, 5.557674e-05, 
    5.557666e-05, 5.557637e-05, 5.55765e-05, 5.55761e-05, 5.557601e-05, 
    5.557593e-05, 5.557582e-05, 5.557581e-05, 5.557575e-05, 5.557585e-05, 
    5.557575e-05, 5.557611e-05, 5.557595e-05, 5.55764e-05, 5.557629e-05, 
    5.557634e-05, 5.557639e-05, 5.557623e-05, 5.557605e-05, 5.557604e-05, 
    5.557598e-05, 5.557582e-05, 5.55761e-05, 5.557524e-05, 5.557577e-05, 
    5.557657e-05, 5.557641e-05, 5.557638e-05, 5.557645e-05, 5.557602e-05, 
    5.557617e-05, 5.557575e-05, 5.557586e-05, 5.557568e-05, 5.557577e-05, 
    5.557578e-05, 5.55759e-05, 5.557598e-05, 5.557616e-05, 5.557631e-05, 
    5.557643e-05, 5.557641e-05, 5.557627e-05, 5.557603e-05, 5.557581e-05, 
    5.557586e-05, 5.557569e-05, 5.557613e-05, 5.557595e-05, 5.557602e-05, 
    5.557583e-05, 5.557624e-05, 5.557589e-05, 5.557633e-05, 5.557629e-05, 
    5.557617e-05, 5.557594e-05, 5.557588e-05, 5.557583e-05, 5.557586e-05, 
    5.557603e-05, 5.557606e-05, 5.557618e-05, 5.557621e-05, 5.55763e-05, 
    5.557638e-05, 5.557631e-05, 5.557623e-05, 5.557603e-05, 5.557585e-05, 
    5.557565e-05, 5.557559e-05, 5.557536e-05, 5.557555e-05, 5.557524e-05, 
    5.55755e-05, 5.557504e-05, 5.557587e-05, 5.557551e-05, 5.557617e-05, 
    5.55761e-05, 5.557597e-05, 5.557568e-05, 5.557583e-05, 5.557565e-05, 
    5.557606e-05, 5.557627e-05, 5.557633e-05, 5.557643e-05, 5.557632e-05, 
    5.557633e-05, 5.557623e-05, 5.557626e-05, 5.557602e-05, 5.557615e-05, 
    5.557578e-05, 5.557565e-05, 5.557527e-05, 5.557504e-05, 5.557481e-05, 
    5.55747e-05, 5.557467e-05, 5.557466e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR1_HR =
  7.799529e-13, 7.820892e-13, 7.816743e-13, 7.83396e-13, 7.824413e-13, 
    7.835683e-13, 7.803865e-13, 7.821737e-13, 7.810331e-13, 7.801458e-13, 
    7.867332e-13, 7.834728e-13, 7.901189e-13, 7.880421e-13, 7.93257e-13, 
    7.897954e-13, 7.939545e-13, 7.93158e-13, 7.955565e-13, 7.948696e-13, 
    7.979333e-13, 7.958735e-13, 7.995212e-13, 7.97442e-13, 7.977671e-13, 
    7.958054e-13, 7.8413e-13, 7.863272e-13, 7.839996e-13, 7.843131e-13, 
    7.841726e-13, 7.824607e-13, 7.815972e-13, 7.797901e-13, 7.801184e-13, 
    7.814459e-13, 7.84454e-13, 7.834338e-13, 7.860059e-13, 7.859479e-13, 
    7.88808e-13, 7.875188e-13, 7.92322e-13, 7.909579e-13, 7.948983e-13, 
    7.939079e-13, 7.948517e-13, 7.945656e-13, 7.948554e-13, 7.934026e-13, 
    7.940251e-13, 7.927466e-13, 7.877602e-13, 7.892264e-13, 7.848505e-13, 
    7.822149e-13, 7.804648e-13, 7.792217e-13, 7.793974e-13, 7.797323e-13, 
    7.814537e-13, 7.830717e-13, 7.84304e-13, 7.851279e-13, 7.859395e-13, 
    7.883927e-13, 7.896919e-13, 7.925973e-13, 7.920739e-13, 7.929611e-13, 
    7.938093e-13, 7.952318e-13, 7.949979e-13, 7.956242e-13, 7.929382e-13, 
    7.947234e-13, 7.917756e-13, 7.925821e-13, 7.861575e-13, 7.837092e-13, 
    7.826657e-13, 7.817539e-13, 7.795325e-13, 7.810666e-13, 7.804619e-13, 
    7.819009e-13, 7.828145e-13, 7.823628e-13, 7.851504e-13, 7.840669e-13, 
    7.897689e-13, 7.873144e-13, 7.937104e-13, 7.921814e-13, 7.940768e-13, 
    7.931099e-13, 7.947662e-13, 7.932757e-13, 7.958575e-13, 7.96419e-13, 
    7.960352e-13, 7.9751e-13, 7.931929e-13, 7.948514e-13, 7.8235e-13, 
    7.824237e-13, 7.827671e-13, 7.812571e-13, 7.811648e-13, 7.79781e-13, 
    7.810126e-13, 7.815366e-13, 7.828676e-13, 7.836542e-13, 7.844018e-13, 
    7.860449e-13, 7.878783e-13, 7.904407e-13, 7.922805e-13, 7.935129e-13, 
    7.927575e-13, 7.934244e-13, 7.926787e-13, 7.923293e-13, 7.962084e-13, 
    7.940307e-13, 7.972979e-13, 7.971174e-13, 7.95639e-13, 7.971377e-13, 
    7.824754e-13, 7.820515e-13, 7.805781e-13, 7.817312e-13, 7.796303e-13, 
    7.808061e-13, 7.814818e-13, 7.840889e-13, 7.84662e-13, 7.851926e-13, 
    7.862406e-13, 7.875848e-13, 7.899409e-13, 7.919896e-13, 7.938587e-13, 
    7.937219e-13, 7.937701e-13, 7.941871e-13, 7.931535e-13, 7.943568e-13, 
    7.945585e-13, 7.940308e-13, 7.970931e-13, 7.962187e-13, 7.971135e-13, 
    7.965443e-13, 7.821893e-13, 7.829028e-13, 7.825172e-13, 7.832421e-13, 
    7.827312e-13, 7.850012e-13, 7.856814e-13, 7.888627e-13, 7.875582e-13, 
    7.896347e-13, 7.877694e-13, 7.880998e-13, 7.897013e-13, 7.878704e-13, 
    7.918762e-13, 7.891601e-13, 7.942034e-13, 7.914925e-13, 7.943731e-13, 
    7.938507e-13, 7.947159e-13, 7.954901e-13, 7.964645e-13, 7.982603e-13, 
    7.978447e-13, 7.993462e-13, 7.839663e-13, 7.848909e-13, 7.848099e-13, 
    7.857775e-13, 7.864928e-13, 7.88043e-13, 7.905268e-13, 7.895933e-13, 
    7.913075e-13, 7.916513e-13, 7.890472e-13, 7.906459e-13, 7.855098e-13, 
    7.863398e-13, 7.85846e-13, 7.84039e-13, 7.898077e-13, 7.868485e-13, 
    7.923108e-13, 7.907098e-13, 7.953797e-13, 7.930578e-13, 7.976157e-13, 
    7.995603e-13, 8.013912e-13, 8.035263e-13, 7.853958e-13, 7.847678e-13, 
    7.858927e-13, 7.874475e-13, 7.888907e-13, 7.908074e-13, 7.910037e-13, 
    7.913624e-13, 7.92292e-13, 7.930731e-13, 7.914753e-13, 7.932689e-13, 
    7.865313e-13, 7.900647e-13, 7.845298e-13, 7.86197e-13, 7.873561e-13, 
    7.868482e-13, 7.894866e-13, 7.901079e-13, 7.926309e-13, 7.913273e-13, 
    7.9908e-13, 7.95653e-13, 8.051523e-13, 8.025013e-13, 7.845481e-13, 
    7.853939e-13, 7.883347e-13, 7.86936e-13, 7.909355e-13, 7.919188e-13, 
    7.927183e-13, 7.937392e-13, 7.938497e-13, 7.944544e-13, 7.934634e-13, 
    7.944155e-13, 7.908114e-13, 7.924227e-13, 7.879994e-13, 7.890764e-13, 
    7.885811e-13, 7.880374e-13, 7.89715e-13, 7.915003e-13, 7.915393e-13, 
    7.921113e-13, 7.937212e-13, 7.909517e-13, 7.995205e-13, 7.942308e-13, 
    7.863158e-13, 7.879426e-13, 7.881758e-13, 7.875456e-13, 7.918202e-13, 
    7.902721e-13, 7.944398e-13, 7.933143e-13, 7.951584e-13, 7.942421e-13, 
    7.941072e-13, 7.929301e-13, 7.921967e-13, 7.903429e-13, 7.88834e-13, 
    7.876372e-13, 7.879156e-13, 7.892301e-13, 7.916097e-13, 7.938594e-13, 
    7.933666e-13, 7.950182e-13, 7.906457e-13, 7.924797e-13, 7.917707e-13, 
    7.936191e-13, 7.895683e-13, 7.930157e-13, 7.88686e-13, 7.890661e-13, 
    7.902414e-13, 7.926035e-13, 7.93127e-13, 7.936844e-13, 7.933407e-13, 
    7.916702e-13, 7.913968e-13, 7.90213e-13, 7.898857e-13, 7.889834e-13, 
    7.882359e-13, 7.889187e-13, 7.896354e-13, 7.916713e-13, 7.935041e-13, 
    7.95501e-13, 7.959898e-13, 7.983186e-13, 7.96422e-13, 7.995498e-13, 
    7.968891e-13, 8.014938e-13, 7.932166e-13, 7.968125e-13, 7.902951e-13, 
    7.909982e-13, 7.922687e-13, 7.951818e-13, 7.936104e-13, 7.954485e-13, 
    7.913862e-13, 7.89275e-13, 7.887295e-13, 7.877098e-13, 7.887528e-13, 
    7.88668e-13, 7.896657e-13, 7.893452e-13, 7.917389e-13, 7.904534e-13, 
    7.941036e-13, 7.954341e-13, 7.991886e-13, 8.014867e-13, 8.038249e-13, 
    8.048561e-13, 8.051699e-13, 8.05301e-13 ;

 LITR2C =
  1.939613e-05, 1.939611e-05, 1.939611e-05, 1.93961e-05, 1.93961e-05, 
    1.939609e-05, 1.939612e-05, 1.939611e-05, 1.939612e-05, 1.939612e-05, 
    1.939606e-05, 1.939609e-05, 1.939603e-05, 1.939605e-05, 1.9396e-05, 
    1.939603e-05, 1.9396e-05, 1.9396e-05, 1.939598e-05, 1.939599e-05, 
    1.939596e-05, 1.939598e-05, 1.939595e-05, 1.939596e-05, 1.939596e-05, 
    1.939598e-05, 1.939609e-05, 1.939607e-05, 1.939609e-05, 1.939609e-05, 
    1.939609e-05, 1.93961e-05, 1.939611e-05, 1.939613e-05, 1.939612e-05, 
    1.939611e-05, 1.939608e-05, 1.93961e-05, 1.939607e-05, 1.939607e-05, 
    1.939604e-05, 1.939606e-05, 1.939601e-05, 1.939602e-05, 1.939599e-05, 
    1.9396e-05, 1.939599e-05, 1.939599e-05, 1.939599e-05, 1.9396e-05, 
    1.9396e-05, 1.939601e-05, 1.939605e-05, 1.939604e-05, 1.939608e-05, 
    1.939611e-05, 1.939612e-05, 1.939613e-05, 1.939613e-05, 1.939613e-05, 
    1.939611e-05, 1.93961e-05, 1.939609e-05, 1.939608e-05, 1.939607e-05, 
    1.939605e-05, 1.939604e-05, 1.939601e-05, 1.939601e-05, 1.939601e-05, 
    1.9396e-05, 1.939598e-05, 1.939599e-05, 1.939598e-05, 1.939601e-05, 
    1.939599e-05, 1.939602e-05, 1.939601e-05, 1.939607e-05, 1.939609e-05, 
    1.93961e-05, 1.939611e-05, 1.939613e-05, 1.939612e-05, 1.939612e-05, 
    1.939611e-05, 1.93961e-05, 1.93961e-05, 1.939608e-05, 1.939609e-05, 
    1.939603e-05, 1.939606e-05, 1.9396e-05, 1.939601e-05, 1.939599e-05, 
    1.9396e-05, 1.939599e-05, 1.9396e-05, 1.939598e-05, 1.939597e-05, 
    1.939598e-05, 1.939596e-05, 1.9396e-05, 1.939599e-05, 1.93961e-05, 
    1.93961e-05, 1.93961e-05, 1.939612e-05, 1.939612e-05, 1.939613e-05, 
    1.939612e-05, 1.939611e-05, 1.93961e-05, 1.939609e-05, 1.939609e-05, 
    1.939607e-05, 1.939605e-05, 1.939603e-05, 1.939601e-05, 1.9396e-05, 
    1.939601e-05, 1.9396e-05, 1.939601e-05, 1.939601e-05, 1.939597e-05, 
    1.9396e-05, 1.939597e-05, 1.939597e-05, 1.939598e-05, 1.939597e-05, 
    1.93961e-05, 1.939611e-05, 1.939612e-05, 1.939611e-05, 1.939613e-05, 
    1.939612e-05, 1.939611e-05, 1.939609e-05, 1.939608e-05, 1.939608e-05, 
    1.939607e-05, 1.939605e-05, 1.939603e-05, 1.939601e-05, 1.9396e-05, 
    1.9396e-05, 1.9396e-05, 1.939599e-05, 1.9396e-05, 1.939599e-05, 
    1.939599e-05, 1.9396e-05, 1.939597e-05, 1.939597e-05, 1.939597e-05, 
    1.939597e-05, 1.939611e-05, 1.93961e-05, 1.93961e-05, 1.93961e-05, 
    1.93961e-05, 1.939608e-05, 1.939607e-05, 1.939604e-05, 1.939606e-05, 
    1.939604e-05, 1.939605e-05, 1.939605e-05, 1.939604e-05, 1.939605e-05, 
    1.939602e-05, 1.939604e-05, 1.939599e-05, 1.939602e-05, 1.939599e-05, 
    1.9396e-05, 1.939599e-05, 1.939598e-05, 1.939597e-05, 1.939596e-05, 
    1.939596e-05, 1.939595e-05, 1.939609e-05, 1.939608e-05, 1.939608e-05, 
    1.939607e-05, 1.939607e-05, 1.939605e-05, 1.939603e-05, 1.939604e-05, 
    1.939602e-05, 1.939602e-05, 1.939604e-05, 1.939603e-05, 1.939608e-05, 
    1.939607e-05, 1.939607e-05, 1.939609e-05, 1.939603e-05, 1.939606e-05, 
    1.939601e-05, 1.939603e-05, 1.939598e-05, 1.9396e-05, 1.939596e-05, 
    1.939594e-05, 1.939593e-05, 1.939591e-05, 1.939608e-05, 1.939608e-05, 
    1.939607e-05, 1.939606e-05, 1.939604e-05, 1.939603e-05, 1.939602e-05, 
    1.939602e-05, 1.939601e-05, 1.9396e-05, 1.939602e-05, 1.9396e-05, 
    1.939607e-05, 1.939603e-05, 1.939608e-05, 1.939607e-05, 1.939606e-05, 
    1.939606e-05, 1.939604e-05, 1.939603e-05, 1.939601e-05, 1.939602e-05, 
    1.939595e-05, 1.939598e-05, 1.939589e-05, 1.939592e-05, 1.939608e-05, 
    1.939608e-05, 1.939605e-05, 1.939606e-05, 1.939602e-05, 1.939601e-05, 
    1.939601e-05, 1.9396e-05, 1.9396e-05, 1.939599e-05, 1.9396e-05, 
    1.939599e-05, 1.939603e-05, 1.939601e-05, 1.939605e-05, 1.939604e-05, 
    1.939605e-05, 1.939605e-05, 1.939604e-05, 1.939602e-05, 1.939602e-05, 
    1.939601e-05, 1.9396e-05, 1.939602e-05, 1.939595e-05, 1.939599e-05, 
    1.939607e-05, 1.939605e-05, 1.939605e-05, 1.939606e-05, 1.939602e-05, 
    1.939603e-05, 1.939599e-05, 1.9396e-05, 1.939599e-05, 1.939599e-05, 
    1.939599e-05, 1.939601e-05, 1.939601e-05, 1.939603e-05, 1.939604e-05, 
    1.939605e-05, 1.939605e-05, 1.939604e-05, 1.939602e-05, 1.9396e-05, 
    1.9396e-05, 1.939599e-05, 1.939603e-05, 1.939601e-05, 1.939602e-05, 
    1.9396e-05, 1.939604e-05, 1.939601e-05, 1.939605e-05, 1.939604e-05, 
    1.939603e-05, 1.939601e-05, 1.9396e-05, 1.9396e-05, 1.9396e-05, 
    1.939602e-05, 1.939602e-05, 1.939603e-05, 1.939603e-05, 1.939604e-05, 
    1.939605e-05, 1.939604e-05, 1.939604e-05, 1.939602e-05, 1.9396e-05, 
    1.939598e-05, 1.939598e-05, 1.939596e-05, 1.939597e-05, 1.939594e-05, 
    1.939597e-05, 1.939593e-05, 1.9396e-05, 1.939597e-05, 1.939603e-05, 
    1.939602e-05, 1.939601e-05, 1.939599e-05, 1.9396e-05, 1.939598e-05, 
    1.939602e-05, 1.939604e-05, 1.939605e-05, 1.939605e-05, 1.939604e-05, 
    1.939605e-05, 1.939604e-05, 1.939604e-05, 1.939602e-05, 1.939603e-05, 
    1.939599e-05, 1.939598e-05, 1.939595e-05, 1.939593e-05, 1.939591e-05, 
    1.939589e-05, 1.939589e-05, 1.939589e-05 ;

 LITR2C_TO_SOIL1C =
  1.187703e-13, 1.190959e-13, 1.190327e-13, 1.192951e-13, 1.191496e-13, 
    1.193214e-13, 1.188364e-13, 1.191088e-13, 1.189349e-13, 1.187997e-13, 
    1.198038e-13, 1.193068e-13, 1.203199e-13, 1.200033e-13, 1.207983e-13, 
    1.202706e-13, 1.209046e-13, 1.207832e-13, 1.211488e-13, 1.210441e-13, 
    1.215111e-13, 1.211971e-13, 1.217532e-13, 1.214362e-13, 1.214858e-13, 
    1.211867e-13, 1.19407e-13, 1.197419e-13, 1.193871e-13, 1.194349e-13, 
    1.194135e-13, 1.191525e-13, 1.190209e-13, 1.187455e-13, 1.187955e-13, 
    1.189978e-13, 1.194564e-13, 1.193009e-13, 1.196929e-13, 1.196841e-13, 
    1.201201e-13, 1.199236e-13, 1.206558e-13, 1.204478e-13, 1.210485e-13, 
    1.208975e-13, 1.210414e-13, 1.209978e-13, 1.210419e-13, 1.208205e-13, 
    1.209154e-13, 1.207205e-13, 1.199604e-13, 1.201839e-13, 1.195168e-13, 
    1.191151e-13, 1.188483e-13, 1.186588e-13, 1.186856e-13, 1.187366e-13, 
    1.18999e-13, 1.192457e-13, 1.194335e-13, 1.195591e-13, 1.196828e-13, 
    1.200568e-13, 1.202548e-13, 1.206977e-13, 1.206179e-13, 1.207532e-13, 
    1.208825e-13, 1.210993e-13, 1.210636e-13, 1.211591e-13, 1.207497e-13, 
    1.210218e-13, 1.205724e-13, 1.206954e-13, 1.19716e-13, 1.193428e-13, 
    1.191838e-13, 1.190448e-13, 1.187062e-13, 1.1894e-13, 1.188479e-13, 
    1.190672e-13, 1.192065e-13, 1.191376e-13, 1.195625e-13, 1.193974e-13, 
    1.202666e-13, 1.198924e-13, 1.208674e-13, 1.206343e-13, 1.209233e-13, 
    1.207759e-13, 1.210283e-13, 1.208011e-13, 1.211947e-13, 1.212803e-13, 
    1.212218e-13, 1.214466e-13, 1.207885e-13, 1.210413e-13, 1.191357e-13, 
    1.191469e-13, 1.191992e-13, 1.189691e-13, 1.18955e-13, 1.187441e-13, 
    1.189318e-13, 1.190117e-13, 1.192146e-13, 1.193345e-13, 1.194484e-13, 
    1.196989e-13, 1.199784e-13, 1.20369e-13, 1.206494e-13, 1.208373e-13, 
    1.207221e-13, 1.208238e-13, 1.207101e-13, 1.206569e-13, 1.212482e-13, 
    1.209162e-13, 1.214143e-13, 1.213867e-13, 1.211614e-13, 1.213898e-13, 
    1.191548e-13, 1.190901e-13, 1.188656e-13, 1.190413e-13, 1.187211e-13, 
    1.189003e-13, 1.190033e-13, 1.194007e-13, 1.194881e-13, 1.19569e-13, 
    1.197287e-13, 1.199336e-13, 1.202928e-13, 1.206051e-13, 1.2089e-13, 
    1.208691e-13, 1.208765e-13, 1.209401e-13, 1.207825e-13, 1.209659e-13, 
    1.209967e-13, 1.209162e-13, 1.21383e-13, 1.212497e-13, 1.213862e-13, 
    1.212994e-13, 1.191112e-13, 1.192199e-13, 1.191612e-13, 1.192716e-13, 
    1.191938e-13, 1.195398e-13, 1.196435e-13, 1.201284e-13, 1.199296e-13, 
    1.202461e-13, 1.199618e-13, 1.200121e-13, 1.202563e-13, 1.199772e-13, 
    1.205878e-13, 1.201738e-13, 1.209425e-13, 1.205293e-13, 1.209684e-13, 
    1.208888e-13, 1.210207e-13, 1.211387e-13, 1.212872e-13, 1.21561e-13, 
    1.214976e-13, 1.217265e-13, 1.19382e-13, 1.19523e-13, 1.195106e-13, 
    1.196581e-13, 1.197672e-13, 1.200035e-13, 1.203821e-13, 1.202398e-13, 
    1.205011e-13, 1.205535e-13, 1.201565e-13, 1.204002e-13, 1.196173e-13, 
    1.197438e-13, 1.196686e-13, 1.193931e-13, 1.202725e-13, 1.198214e-13, 
    1.20654e-13, 1.2041e-13, 1.211219e-13, 1.207679e-13, 1.214627e-13, 
    1.217591e-13, 1.220382e-13, 1.223637e-13, 1.196e-13, 1.195042e-13, 
    1.196757e-13, 1.199127e-13, 1.201327e-13, 1.204249e-13, 1.204548e-13, 
    1.205095e-13, 1.206512e-13, 1.207702e-13, 1.205267e-13, 1.208001e-13, 
    1.19773e-13, 1.203117e-13, 1.194679e-13, 1.197221e-13, 1.198988e-13, 
    1.198213e-13, 1.202235e-13, 1.203182e-13, 1.207028e-13, 1.205041e-13, 
    1.216859e-13, 1.211635e-13, 1.226116e-13, 1.222075e-13, 1.194707e-13, 
    1.195997e-13, 1.200479e-13, 1.198347e-13, 1.204444e-13, 1.205943e-13, 
    1.207162e-13, 1.208718e-13, 1.208886e-13, 1.209808e-13, 1.208297e-13, 
    1.209749e-13, 1.204255e-13, 1.206711e-13, 1.199968e-13, 1.20161e-13, 
    1.200855e-13, 1.200026e-13, 1.202583e-13, 1.205305e-13, 1.205364e-13, 
    1.206236e-13, 1.20869e-13, 1.204469e-13, 1.217531e-13, 1.209467e-13, 
    1.197402e-13, 1.199882e-13, 1.200237e-13, 1.199277e-13, 1.205793e-13, 
    1.203433e-13, 1.209786e-13, 1.20807e-13, 1.210881e-13, 1.209484e-13, 
    1.209279e-13, 1.207484e-13, 1.206366e-13, 1.203541e-13, 1.20124e-13, 
    1.199416e-13, 1.19984e-13, 1.201844e-13, 1.205472e-13, 1.208901e-13, 
    1.20815e-13, 1.210668e-13, 1.204002e-13, 1.206798e-13, 1.205717e-13, 
    1.208535e-13, 1.20236e-13, 1.207615e-13, 1.201015e-13, 1.201594e-13, 
    1.203386e-13, 1.206987e-13, 1.207785e-13, 1.208634e-13, 1.20811e-13, 
    1.205564e-13, 1.205147e-13, 1.203343e-13, 1.202844e-13, 1.201468e-13, 
    1.200329e-13, 1.20137e-13, 1.202462e-13, 1.205565e-13, 1.208359e-13, 
    1.211403e-13, 1.212149e-13, 1.215699e-13, 1.212807e-13, 1.217575e-13, 
    1.21352e-13, 1.220539e-13, 1.207921e-13, 1.213403e-13, 1.203468e-13, 
    1.20454e-13, 1.206476e-13, 1.210917e-13, 1.208521e-13, 1.211323e-13, 
    1.205131e-13, 1.201913e-13, 1.201081e-13, 1.199527e-13, 1.201117e-13, 
    1.200988e-13, 1.202508e-13, 1.20202e-13, 1.205668e-13, 1.203709e-13, 
    1.209273e-13, 1.211302e-13, 1.217025e-13, 1.220528e-13, 1.224093e-13, 
    1.225664e-13, 1.226143e-13, 1.226343e-13 ;

 LITR2C_vr =
  0.001107539, 0.001107538, 0.001107538, 0.001107537, 0.001107538, 
    0.001107537, 0.001107539, 0.001107538, 0.001107538, 0.001107539, 
    0.001107535, 0.001107537, 0.001107533, 0.001107535, 0.001107532, 
    0.001107534, 0.001107531, 0.001107532, 0.001107531, 0.001107531, 
    0.001107529, 0.00110753, 0.001107528, 0.00110753, 0.001107529, 
    0.00110753, 0.001107537, 0.001107535, 0.001107537, 0.001107537, 
    0.001107537, 0.001107538, 0.001107538, 0.001107539, 0.001107539, 
    0.001107538, 0.001107536, 0.001107537, 0.001107536, 0.001107536, 
    0.001107534, 0.001107535, 0.001107532, 0.001107533, 0.001107531, 
    0.001107531, 0.001107531, 0.001107531, 0.001107531, 0.001107532, 
    0.001107531, 0.001107532, 0.001107535, 0.001107534, 0.001107536, 
    0.001107538, 0.001107539, 0.001107539, 0.001107539, 0.001107539, 
    0.001107538, 0.001107537, 0.001107537, 0.001107536, 0.001107536, 
    0.001107534, 0.001107534, 0.001107532, 0.001107532, 0.001107532, 
    0.001107531, 0.001107531, 0.001107531, 0.001107531, 0.001107532, 
    0.001107531, 0.001107533, 0.001107532, 0.001107536, 0.001107537, 
    0.001107537, 0.001107538, 0.001107539, 0.001107538, 0.001107539, 
    0.001107538, 0.001107537, 0.001107538, 0.001107536, 0.001107537, 
    0.001107534, 0.001107535, 0.001107532, 0.001107532, 0.001107531, 
    0.001107532, 0.001107531, 0.001107532, 0.00110753, 0.00110753, 
    0.00110753, 0.00110753, 0.001107532, 0.001107531, 0.001107538, 
    0.001107538, 0.001107537, 0.001107538, 0.001107538, 0.001107539, 
    0.001107538, 0.001107538, 0.001107537, 0.001107537, 0.001107536, 
    0.001107536, 0.001107535, 0.001107533, 0.001107532, 0.001107532, 
    0.001107532, 0.001107532, 0.001107532, 0.001107532, 0.00110753, 
    0.001107531, 0.00110753, 0.00110753, 0.001107531, 0.00110753, 
    0.001107538, 0.001107538, 0.001107539, 0.001107538, 0.001107539, 
    0.001107538, 0.001107538, 0.001107537, 0.001107536, 0.001107536, 
    0.001107536, 0.001107535, 0.001107534, 0.001107533, 0.001107531, 
    0.001107532, 0.001107532, 0.001107531, 0.001107532, 0.001107531, 
    0.001107531, 0.001107531, 0.00110753, 0.00110753, 0.00110753, 0.00110753, 
    0.001107538, 0.001107537, 0.001107538, 0.001107537, 0.001107537, 
    0.001107536, 0.001107536, 0.001107534, 0.001107535, 0.001107534, 
    0.001107535, 0.001107535, 0.001107534, 0.001107535, 0.001107533, 
    0.001107534, 0.001107531, 0.001107533, 0.001107531, 0.001107531, 
    0.001107531, 0.001107531, 0.00110753, 0.001107529, 0.001107529, 
    0.001107529, 0.001107537, 0.001107536, 0.001107536, 0.001107536, 
    0.001107535, 0.001107535, 0.001107533, 0.001107534, 0.001107533, 
    0.001107533, 0.001107534, 0.001107533, 0.001107536, 0.001107535, 
    0.001107536, 0.001107537, 0.001107534, 0.001107535, 0.001107532, 
    0.001107533, 0.001107531, 0.001107532, 0.00110753, 0.001107528, 
    0.001107528, 0.001107526, 0.001107536, 0.001107536, 0.001107536, 
    0.001107535, 0.001107534, 0.001107533, 0.001107533, 0.001107533, 
    0.001107532, 0.001107532, 0.001107533, 0.001107532, 0.001107535, 
    0.001107533, 0.001107536, 0.001107536, 0.001107535, 0.001107535, 
    0.001107534, 0.001107533, 0.001107532, 0.001107533, 0.001107529, 
    0.001107531, 0.001107526, 0.001107527, 0.001107536, 0.001107536, 
    0.001107534, 0.001107535, 0.001107533, 0.001107533, 0.001107532, 
    0.001107532, 0.001107531, 0.001107531, 0.001107532, 0.001107531, 
    0.001107533, 0.001107532, 0.001107535, 0.001107534, 0.001107534, 
    0.001107535, 0.001107534, 0.001107533, 0.001107533, 0.001107532, 
    0.001107532, 0.001107533, 0.001107528, 0.001107531, 0.001107535, 
    0.001107535, 0.001107535, 0.001107535, 0.001107533, 0.001107533, 
    0.001107531, 0.001107532, 0.001107531, 0.001107531, 0.001107531, 
    0.001107532, 0.001107532, 0.001107533, 0.001107534, 0.001107535, 
    0.001107535, 0.001107534, 0.001107533, 0.001107531, 0.001107532, 
    0.001107531, 0.001107533, 0.001107532, 0.001107533, 0.001107532, 
    0.001107534, 0.001107532, 0.001107534, 0.001107534, 0.001107533, 
    0.001107532, 0.001107532, 0.001107532, 0.001107532, 0.001107533, 
    0.001107533, 0.001107533, 0.001107534, 0.001107534, 0.001107535, 
    0.001107534, 0.001107534, 0.001107533, 0.001107532, 0.001107531, 
    0.00110753, 0.001107529, 0.00110753, 0.001107528, 0.00110753, 
    0.001107527, 0.001107532, 0.00110753, 0.001107533, 0.001107533, 
    0.001107532, 0.001107531, 0.001107532, 0.001107531, 0.001107533, 
    0.001107534, 0.001107534, 0.001107535, 0.001107534, 0.001107534, 
    0.001107534, 0.001107534, 0.001107533, 0.001107533, 0.001107531, 
    0.001107531, 0.001107529, 0.001107527, 0.001107526, 0.001107526, 
    0.001107526, 0.001107525,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N =
  2.684281e-07, 2.684279e-07, 2.684279e-07, 2.684277e-07, 2.684278e-07, 
    2.684277e-07, 2.684281e-07, 2.684278e-07, 2.68428e-07, 2.684281e-07, 
    2.684273e-07, 2.684277e-07, 2.684268e-07, 2.684271e-07, 2.684264e-07, 
    2.684269e-07, 2.684263e-07, 2.684264e-07, 2.684261e-07, 2.684262e-07, 
    2.684258e-07, 2.684261e-07, 2.684256e-07, 2.684259e-07, 2.684259e-07, 
    2.684261e-07, 2.684276e-07, 2.684273e-07, 2.684276e-07, 2.684276e-07, 
    2.684276e-07, 2.684278e-07, 2.684279e-07, 2.684282e-07, 2.684281e-07, 
    2.68428e-07, 2.684276e-07, 2.684277e-07, 2.684274e-07, 2.684274e-07, 
    2.68427e-07, 2.684272e-07, 2.684265e-07, 2.684267e-07, 2.684262e-07, 
    2.684263e-07, 2.684262e-07, 2.684262e-07, 2.684262e-07, 2.684264e-07, 
    2.684263e-07, 2.684265e-07, 2.684271e-07, 2.684269e-07, 2.684275e-07, 
    2.684278e-07, 2.684281e-07, 2.684282e-07, 2.684282e-07, 2.684282e-07, 
    2.68428e-07, 2.684277e-07, 2.684276e-07, 2.684275e-07, 2.684274e-07, 
    2.68427e-07, 2.684269e-07, 2.684265e-07, 2.684266e-07, 2.684264e-07, 
    2.684264e-07, 2.684262e-07, 2.684262e-07, 2.684261e-07, 2.684265e-07, 
    2.684262e-07, 2.684266e-07, 2.684265e-07, 2.684273e-07, 2.684276e-07, 
    2.684278e-07, 2.684279e-07, 2.684282e-07, 2.68428e-07, 2.684281e-07, 
    2.684279e-07, 2.684278e-07, 2.684278e-07, 2.684275e-07, 2.684276e-07, 
    2.684269e-07, 2.684272e-07, 2.684264e-07, 2.684266e-07, 2.684263e-07, 
    2.684264e-07, 2.684262e-07, 2.684264e-07, 2.684261e-07, 2.68426e-07, 
    2.684261e-07, 2.684259e-07, 2.684264e-07, 2.684262e-07, 2.684278e-07, 
    2.684278e-07, 2.684278e-07, 2.68428e-07, 2.68428e-07, 2.684282e-07, 
    2.68428e-07, 2.684279e-07, 2.684278e-07, 2.684277e-07, 2.684276e-07, 
    2.684274e-07, 2.684271e-07, 2.684268e-07, 2.684266e-07, 2.684264e-07, 
    2.684265e-07, 2.684264e-07, 2.684265e-07, 2.684265e-07, 2.68426e-07, 
    2.684263e-07, 2.684259e-07, 2.684259e-07, 2.684261e-07, 2.684259e-07, 
    2.684278e-07, 2.684279e-07, 2.68428e-07, 2.684279e-07, 2.684282e-07, 
    2.68428e-07, 2.684279e-07, 2.684276e-07, 2.684275e-07, 2.684275e-07, 
    2.684273e-07, 2.684272e-07, 2.684268e-07, 2.684266e-07, 2.684263e-07, 
    2.684264e-07, 2.684264e-07, 2.684263e-07, 2.684264e-07, 2.684263e-07, 
    2.684262e-07, 2.684263e-07, 2.684259e-07, 2.68426e-07, 2.684259e-07, 
    2.68426e-07, 2.684278e-07, 2.684278e-07, 2.684278e-07, 2.684277e-07, 
    2.684278e-07, 2.684275e-07, 2.684274e-07, 2.68427e-07, 2.684272e-07, 
    2.684269e-07, 2.684271e-07, 2.684271e-07, 2.684269e-07, 2.684271e-07, 
    2.684266e-07, 2.68427e-07, 2.684263e-07, 2.684266e-07, 2.684263e-07, 
    2.684263e-07, 2.684262e-07, 2.684261e-07, 2.68426e-07, 2.684258e-07, 
    2.684258e-07, 2.684257e-07, 2.684276e-07, 2.684275e-07, 2.684275e-07, 
    2.684274e-07, 2.684273e-07, 2.684271e-07, 2.684268e-07, 2.684269e-07, 
    2.684267e-07, 2.684266e-07, 2.68427e-07, 2.684268e-07, 2.684274e-07, 
    2.684273e-07, 2.684274e-07, 2.684276e-07, 2.684269e-07, 2.684272e-07, 
    2.684265e-07, 2.684268e-07, 2.684261e-07, 2.684264e-07, 2.684259e-07, 
    2.684256e-07, 2.684254e-07, 2.684251e-07, 2.684274e-07, 2.684275e-07, 
    2.684274e-07, 2.684272e-07, 2.68427e-07, 2.684267e-07, 2.684267e-07, 
    2.684267e-07, 2.684265e-07, 2.684264e-07, 2.684266e-07, 2.684264e-07, 
    2.684273e-07, 2.684268e-07, 2.684276e-07, 2.684273e-07, 2.684272e-07, 
    2.684272e-07, 2.684269e-07, 2.684268e-07, 2.684265e-07, 2.684267e-07, 
    2.684257e-07, 2.684261e-07, 2.684249e-07, 2.684252e-07, 2.684276e-07, 
    2.684274e-07, 2.68427e-07, 2.684272e-07, 2.684267e-07, 2.684266e-07, 
    2.684265e-07, 2.684264e-07, 2.684263e-07, 2.684263e-07, 2.684264e-07, 
    2.684263e-07, 2.684267e-07, 2.684265e-07, 2.684271e-07, 2.68427e-07, 
    2.68427e-07, 2.684271e-07, 2.684269e-07, 2.684266e-07, 2.684266e-07, 
    2.684266e-07, 2.684264e-07, 2.684267e-07, 2.684256e-07, 2.684263e-07, 
    2.684273e-07, 2.684271e-07, 2.684271e-07, 2.684272e-07, 2.684266e-07, 
    2.684268e-07, 2.684263e-07, 2.684264e-07, 2.684262e-07, 2.684263e-07, 
    2.684263e-07, 2.684265e-07, 2.684266e-07, 2.684268e-07, 2.68427e-07, 
    2.684272e-07, 2.684271e-07, 2.684269e-07, 2.684266e-07, 2.684263e-07, 
    2.684264e-07, 2.684262e-07, 2.684268e-07, 2.684265e-07, 2.684266e-07, 
    2.684264e-07, 2.684269e-07, 2.684264e-07, 2.68427e-07, 2.68427e-07, 
    2.684268e-07, 2.684265e-07, 2.684264e-07, 2.684264e-07, 2.684264e-07, 
    2.684266e-07, 2.684267e-07, 2.684268e-07, 2.684268e-07, 2.68427e-07, 
    2.684271e-07, 2.68427e-07, 2.684269e-07, 2.684266e-07, 2.684264e-07, 
    2.684261e-07, 2.684261e-07, 2.684258e-07, 2.68426e-07, 2.684256e-07, 
    2.68426e-07, 2.684254e-07, 2.684264e-07, 2.68426e-07, 2.684268e-07, 
    2.684267e-07, 2.684266e-07, 2.684262e-07, 2.684264e-07, 2.684261e-07, 
    2.684267e-07, 2.684269e-07, 2.68427e-07, 2.684271e-07, 2.68427e-07, 
    2.68427e-07, 2.684269e-07, 2.684269e-07, 2.684266e-07, 2.684268e-07, 
    2.684263e-07, 2.684261e-07, 2.684257e-07, 2.684254e-07, 2.684251e-07, 
    2.684249e-07, 2.684249e-07, 2.684249e-07 ;

 LITR2N_TNDNCY_VERT_TRANS =
  -2.450906e-27, 9.313441e-26, 2.205815e-25, 1.151926e-25, 1.715634e-26, 
    2.205815e-26, -2.009742e-25, 1.470543e-26, -4.901811e-26, -1.176435e-25, 
    -1.715634e-25, -5.882173e-26, -1.617598e-25, 9.313441e-26, -3.921449e-26, 
    9.803622e-27, 5.882173e-26, 2.32836e-25, 2.132288e-25, -5.882173e-26, 
    1.225453e-26, 6.862535e-26, 4.41163e-26, -1.004871e-25, 3.676358e-26, 
    8.333079e-26, -1.274471e-25, -1.838179e-25, 8.087988e-26, -2.205815e-26, 
    -9.068351e-26, -1.985233e-25, 1.225453e-26, -1.323489e-25, -1.519561e-25, 
    7.842898e-26, 5.882173e-26, 8.82326e-26, -1.004871e-25, -1.176435e-25, 
    1.593089e-25, 1.789161e-25, 7.107626e-26, 2.475414e-25, 1.347998e-25, 
    -1.715634e-25, 2.009742e-25, -9.803622e-27, -1.02938e-25, -3.333231e-25, 
    5.146902e-26, -1.225453e-25, -1.053889e-25, -2.32836e-25, -7.597807e-26, 
    3.921449e-26, 2.695996e-26, -2.303851e-25, 2.450906e-27, -2.352869e-25, 
    1.397016e-25, -4.41163e-26, -1.960724e-25, 2.695996e-26, 2.524433e-25, 
    1.151926e-25, -9.068351e-26, -1.593089e-25, -1.764652e-25, -2.132288e-25, 
    1.617598e-25, 1.715634e-26, 1.495052e-25, -5.637083e-26, -1.470543e-25, 
    4.166539e-26, 1.102908e-25, 1.862688e-25, -9.313441e-26, 9.803622e-27, 
    -8.578169e-26, 3.921449e-26, 4.901811e-27, -1.715634e-25, -5.146902e-26, 
    6.617445e-26, 3.676358e-26, 2.450905e-26, -1.29898e-25, 4.65672e-26, 
    1.323489e-25, 1.02938e-25, 2.990105e-25, -1.397016e-25, 9.313441e-26, 
    2.009742e-25, 6.617445e-26, -2.941087e-26, -4.901811e-26, 3.186177e-26, 
    2.426396e-25, 3.38225e-25, 7.107626e-26, -1.642107e-25, 9.068351e-26, 
    1.249962e-25, -1.372507e-25, -4.166539e-26, -1.200944e-25, -8.82326e-26, 
    1.593089e-25, 2.181306e-25, 2.59796e-25, -2.769523e-25, 3.676358e-26, 
    -2.941087e-26, -1.274471e-25, -9.313441e-26, 1.176435e-25, 1.446034e-25, 
    2.034252e-25, -2.450906e-27, 5.146902e-26, 3.676358e-26, -5.146902e-26, 
    4.901811e-26, -1.372507e-25, 1.593089e-25, 3.186177e-26, 4.901811e-26, 
    4.901811e-27, -5.882173e-26, -4.901811e-26, 1.617598e-25, 1.764652e-25, 
    3.186177e-26, -6.127264e-26, -4.65672e-26, 2.352869e-25, 8.578169e-26, 
    -1.249962e-25, -5.146902e-26, -1.495052e-25, 9.803622e-27, 1.200944e-25, 
    1.274471e-25, 4.901811e-27, -3.676358e-26, -4.65672e-26, -3.62734e-25, 
    -1.02938e-25, 9.558531e-26, 1.911706e-25, 1.274471e-25, 7.597807e-26, 
    -6.617445e-26, 2.205815e-26, 1.715634e-26, 2.205815e-26, -1.691125e-25, 
    -7.107626e-26, -3.431268e-26, 2.671487e-25, 4.41163e-26, -4.65672e-26, 
    2.377378e-25, 9.558531e-26, 8.333079e-26, 9.803622e-27, -1.985233e-25, 
    -1.29898e-25, -4.65672e-26, 4.901811e-26, 1.593089e-25, 1.470543e-26, 
    -1.323489e-25, -5.882173e-26, 3.676358e-26, 2.009742e-25, -2.450905e-26, 
    -1.519561e-25, 2.941087e-26, -1.053889e-25, -1.29898e-25, 1.470543e-25, 
    -9.803622e-27, -5.391992e-26, 1.397016e-25, 1.004871e-25, -1.078398e-25, 
    1.495052e-25, 1.323489e-25, -2.450905e-26, 2.695996e-26, -7.352717e-27, 
    -1.225453e-26, -1.446034e-25, -7.597807e-26, -7.352717e-27, 
    -6.127264e-26, 7.352717e-26, 2.181306e-25, 1.323489e-25, 1.053889e-25, 
    9.068351e-26, -9.803622e-27, 1.985233e-25, -1.715634e-26, -1.740143e-25, 
    -4.65672e-26, 1.347998e-25, -2.475414e-25, 1.470543e-25, -1.200944e-25, 
    -1.470543e-25, 1.078398e-25, 6.127264e-26, 1.225453e-25, -8.087988e-26, 
    2.303851e-25, 2.450905e-26, -6.862535e-26, -6.862535e-26, 1.053889e-25, 
    2.941087e-26, 1.838179e-25, -3.38225e-25, 2.426396e-25, -7.597807e-26, 
    1.421525e-25, -3.014614e-25, -1.593089e-25, -2.08327e-25, 6.127264e-26, 
    1.495052e-25, -7.597807e-26, -1.642107e-25, 7.842898e-26, -1.372507e-25, 
    -2.695996e-26, -1.764652e-25, -2.695996e-26, -7.107626e-26, 
    -8.578169e-26, -7.597807e-26, -1.102908e-25, 7.352717e-27, -1.078398e-25, 
    5.882173e-26, -1.715634e-26, 2.695996e-26, -4.901811e-27, -1.446034e-25, 
    -1.02938e-25, -2.426396e-25, -7.842898e-26, 9.068351e-26, -9.068351e-26, 
    -1.225453e-26, 1.151926e-25, 5.146902e-26, -2.32836e-25, -4.65672e-26, 
    -1.470543e-26, -5.882173e-26, -5.391992e-26, -7.597807e-26, 1.078398e-25, 
    9.558531e-26, -1.02938e-25, -8.333079e-26, -3.676358e-26, -1.02938e-25, 
    1.740143e-25, 4.65672e-26, 3.431268e-26, 1.225453e-26, -1.495052e-25, 
    1.960724e-25, 1.642107e-25, -9.803622e-26, 1.053889e-25, 4.41163e-26, 
    -2.941087e-26, -2.695996e-25, -1.225453e-25, -4.901811e-27, 3.921449e-26, 
    1.225453e-26, 1.397016e-25, 1.225453e-25, 2.205815e-26, 1.102908e-25, 
    -1.127417e-25, 1.323489e-25, -2.205815e-25, -1.249962e-25, 3.676358e-26, 
    -1.127417e-25, 4.901811e-27, 2.352869e-25, 1.666616e-25, 1.764652e-25, 
    3.431268e-26, 1.225453e-25, -8.333079e-26, -4.901811e-27, 1.764652e-25, 
    -1.004871e-25, 2.450906e-27, -4.901811e-27, -3.431268e-26, -5.637083e-26, 
    -3.014614e-25, -1.764652e-25, -2.230324e-25, -1.764652e-25, 1.715634e-26, 
    9.803622e-27, -2.745014e-25, -1.642107e-25, -1.593089e-25, 2.450906e-27, 
    -5.391992e-26, -1.004871e-25, 2.450906e-27, -5.391992e-26, -3.431268e-26, 
    7.107626e-26, 1.004871e-25, -6.862535e-26, -1.347998e-25, 6.127264e-26, 
    1.470543e-26, -4.65672e-26, -5.391992e-26, 1.372507e-25, -1.838179e-25,
  2.676268e-32, 2.676265e-32, 2.676265e-32, 2.676263e-32, 2.676264e-32, 
    2.676263e-32, 2.676267e-32, 2.676265e-32, 2.676266e-32, 2.676267e-32, 
    2.676259e-32, 2.676263e-32, 2.676254e-32, 2.676257e-32, 2.67625e-32, 
    2.676255e-32, 2.676249e-32, 2.676251e-32, 2.676247e-32, 2.676248e-32, 
    2.676244e-32, 2.676247e-32, 2.676242e-32, 2.676245e-32, 2.676244e-32, 
    2.676247e-32, 2.676262e-32, 2.676259e-32, 2.676262e-32, 2.676262e-32, 
    2.676262e-32, 2.676264e-32, 2.676266e-32, 2.676268e-32, 2.676267e-32, 
    2.676266e-32, 2.676262e-32, 2.676263e-32, 2.67626e-32, 2.67626e-32, 
    2.676256e-32, 2.676258e-32, 2.676252e-32, 2.676253e-32, 2.676248e-32, 
    2.676249e-32, 2.676248e-32, 2.676249e-32, 2.676248e-32, 2.67625e-32, 
    2.676249e-32, 2.676251e-32, 2.676257e-32, 2.676256e-32, 2.676261e-32, 
    2.676265e-32, 2.676267e-32, 2.676269e-32, 2.676268e-32, 2.676268e-32, 
    2.676266e-32, 2.676264e-32, 2.676262e-32, 2.676261e-32, 2.67626e-32, 
    2.676257e-32, 2.676255e-32, 2.676251e-32, 2.676252e-32, 2.676251e-32, 
    2.67625e-32, 2.676248e-32, 2.676248e-32, 2.676247e-32, 2.676251e-32, 
    2.676249e-32, 2.676252e-32, 2.676251e-32, 2.67626e-32, 2.676263e-32, 
    2.676264e-32, 2.676265e-32, 2.676268e-32, 2.676266e-32, 2.676267e-32, 
    2.676265e-32, 2.676264e-32, 2.676264e-32, 2.676261e-32, 2.676262e-32, 
    2.676255e-32, 2.676258e-32, 2.67625e-32, 2.676252e-32, 2.676249e-32, 
    2.676251e-32, 2.676249e-32, 2.67625e-32, 2.676247e-32, 2.676246e-32, 
    2.676247e-32, 2.676245e-32, 2.676251e-32, 2.676248e-32, 2.676264e-32, 
    2.676264e-32, 2.676264e-32, 2.676266e-32, 2.676266e-32, 2.676268e-32, 
    2.676266e-32, 2.676266e-32, 2.676264e-32, 2.676263e-32, 2.676262e-32, 
    2.67626e-32, 2.676257e-32, 2.676254e-32, 2.676252e-32, 2.67625e-32, 
    2.676251e-32, 2.67625e-32, 2.676251e-32, 2.676252e-32, 2.676247e-32, 
    2.676249e-32, 2.676245e-32, 2.676245e-32, 2.676247e-32, 2.676245e-32, 
    2.676264e-32, 2.676265e-32, 2.676267e-32, 2.676265e-32, 2.676268e-32, 
    2.676267e-32, 2.676266e-32, 2.676262e-32, 2.676262e-32, 2.676261e-32, 
    2.676259e-32, 2.676258e-32, 2.676255e-32, 2.676252e-32, 2.67625e-32, 
    2.67625e-32, 2.67625e-32, 2.676249e-32, 2.676251e-32, 2.676249e-32, 
    2.676249e-32, 2.676249e-32, 2.676245e-32, 2.676247e-32, 2.676245e-32, 
    2.676246e-32, 2.676265e-32, 2.676264e-32, 2.676264e-32, 2.676263e-32, 
    2.676264e-32, 2.676261e-32, 2.67626e-32, 2.676256e-32, 2.676258e-32, 
    2.676255e-32, 2.676257e-32, 2.676257e-32, 2.676255e-32, 2.676257e-32, 
    2.676252e-32, 2.676256e-32, 2.676249e-32, 2.676253e-32, 2.676249e-32, 
    2.67625e-32, 2.676249e-32, 2.676247e-32, 2.676246e-32, 2.676244e-32, 
    2.676244e-32, 2.676243e-32, 2.676262e-32, 2.676261e-32, 2.676261e-32, 
    2.67626e-32, 2.676259e-32, 2.676257e-32, 2.676254e-32, 2.676255e-32, 
    2.676253e-32, 2.676252e-32, 2.676256e-32, 2.676254e-32, 2.67626e-32, 
    2.676259e-32, 2.67626e-32, 2.676262e-32, 2.676255e-32, 2.676259e-32, 
    2.676252e-32, 2.676254e-32, 2.676248e-32, 2.676251e-32, 2.676245e-32, 
    2.676242e-32, 2.67624e-32, 2.676237e-32, 2.676261e-32, 2.676262e-32, 
    2.67626e-32, 2.676258e-32, 2.676256e-32, 2.676254e-32, 2.676253e-32, 
    2.676253e-32, 2.676252e-32, 2.676251e-32, 2.676253e-32, 2.67625e-32, 
    2.676259e-32, 2.676254e-32, 2.676262e-32, 2.676259e-32, 2.676258e-32, 
    2.676259e-32, 2.676255e-32, 2.676254e-32, 2.676251e-32, 2.676253e-32, 
    2.676243e-32, 2.676247e-32, 2.676235e-32, 2.676239e-32, 2.676262e-32, 
    2.676261e-32, 2.676257e-32, 2.676259e-32, 2.676254e-32, 2.676252e-32, 
    2.676251e-32, 2.67625e-32, 2.67625e-32, 2.676249e-32, 2.67625e-32, 
    2.676249e-32, 2.676254e-32, 2.676252e-32, 2.676257e-32, 2.676256e-32, 
    2.676257e-32, 2.676257e-32, 2.676255e-32, 2.676253e-32, 2.676253e-32, 
    2.676252e-32, 2.67625e-32, 2.676253e-32, 2.676242e-32, 2.676249e-32, 
    2.676259e-32, 2.676257e-32, 2.676257e-32, 2.676258e-32, 2.676252e-32, 
    2.676254e-32, 2.676249e-32, 2.67625e-32, 2.676248e-32, 2.676249e-32, 
    2.676249e-32, 2.676251e-32, 2.676252e-32, 2.676254e-32, 2.676256e-32, 
    2.676258e-32, 2.676257e-32, 2.676256e-32, 2.676253e-32, 2.67625e-32, 
    2.67625e-32, 2.676248e-32, 2.676254e-32, 2.676252e-32, 2.676252e-32, 
    2.67625e-32, 2.676255e-32, 2.676251e-32, 2.676256e-32, 2.676256e-32, 
    2.676254e-32, 2.676251e-32, 2.676251e-32, 2.67625e-32, 2.67625e-32, 
    2.676252e-32, 2.676253e-32, 2.676254e-32, 2.676255e-32, 2.676256e-32, 
    2.676257e-32, 2.676256e-32, 2.676255e-32, 2.676252e-32, 2.67625e-32, 
    2.676247e-32, 2.676247e-32, 2.676244e-32, 2.676246e-32, 2.676242e-32, 
    2.676246e-32, 2.67624e-32, 2.67625e-32, 2.676246e-32, 2.676254e-32, 
    2.676253e-32, 2.676252e-32, 2.676248e-32, 2.67625e-32, 2.676248e-32, 
    2.676253e-32, 2.676256e-32, 2.676256e-32, 2.676258e-32, 2.676256e-32, 
    2.676256e-32, 2.676255e-32, 2.676256e-32, 2.676252e-32, 2.676254e-32, 
    2.676249e-32, 2.676248e-32, 2.676243e-32, 2.67624e-32, 2.676237e-32, 
    2.676235e-32, 2.676235e-32, 2.676235e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2N_TO_SOIL1N =
  3.287387e-15, 3.2964e-15, 3.294649e-15, 3.301913e-15, 3.297885e-15, 
    3.30264e-15, 3.289216e-15, 3.296756e-15, 3.291944e-15, 3.2882e-15, 
    3.315993e-15, 3.302237e-15, 3.330278e-15, 3.321516e-15, 3.343518e-15, 
    3.328913e-15, 3.346462e-15, 3.343101e-15, 3.353221e-15, 3.350323e-15, 
    3.363249e-15, 3.354558e-15, 3.369949e-15, 3.361176e-15, 3.362548e-15, 
    3.354271e-15, 3.30501e-15, 3.31428e-15, 3.30446e-15, 3.305783e-15, 
    3.30519e-15, 3.297967e-15, 3.294324e-15, 3.2867e-15, 3.288085e-15, 
    3.293685e-15, 3.306377e-15, 3.302073e-15, 3.312925e-15, 3.31268e-15, 
    3.324747e-15, 3.319308e-15, 3.339574e-15, 3.333818e-15, 3.350444e-15, 
    3.346265e-15, 3.350247e-15, 3.34904e-15, 3.350263e-15, 3.344133e-15, 
    3.34676e-15, 3.341365e-15, 3.320326e-15, 3.326512e-15, 3.30805e-15, 
    3.29693e-15, 3.289546e-15, 3.284301e-15, 3.285043e-15, 3.286456e-15, 
    3.293718e-15, 3.300545e-15, 3.305744e-15, 3.30922e-15, 3.312645e-15, 
    3.322995e-15, 3.328477e-15, 3.340735e-15, 3.338527e-15, 3.34227e-15, 
    3.345849e-15, 3.351851e-15, 3.350864e-15, 3.353507e-15, 3.342173e-15, 
    3.349706e-15, 3.337268e-15, 3.340671e-15, 3.313564e-15, 3.303235e-15, 
    3.298832e-15, 3.294985e-15, 3.285613e-15, 3.292085e-15, 3.289534e-15, 
    3.295605e-15, 3.29946e-15, 3.297554e-15, 3.309315e-15, 3.304744e-15, 
    3.328802e-15, 3.318445e-15, 3.345432e-15, 3.338981e-15, 3.346978e-15, 
    3.342898e-15, 3.349886e-15, 3.343597e-15, 3.354491e-15, 3.35686e-15, 
    3.355241e-15, 3.361463e-15, 3.343248e-15, 3.350246e-15, 3.2975e-15, 
    3.297811e-15, 3.29926e-15, 3.292889e-15, 3.292499e-15, 3.286661e-15, 
    3.291857e-15, 3.294068e-15, 3.299684e-15, 3.303002e-15, 3.306157e-15, 
    3.313089e-15, 3.320825e-15, 3.331636e-15, 3.339399e-15, 3.344598e-15, 
    3.341411e-15, 3.344225e-15, 3.341079e-15, 3.339604e-15, 3.355972e-15, 
    3.346783e-15, 3.360568e-15, 3.359807e-15, 3.353569e-15, 3.359892e-15, 
    3.298029e-15, 3.29624e-15, 3.290024e-15, 3.294889e-15, 3.286025e-15, 
    3.290986e-15, 3.293837e-15, 3.304837e-15, 3.307255e-15, 3.309493e-15, 
    3.313915e-15, 3.319586e-15, 3.329527e-15, 3.338171e-15, 3.346058e-15, 
    3.34548e-15, 3.345683e-15, 3.347443e-15, 3.343082e-15, 3.348159e-15, 
    3.34901e-15, 3.346784e-15, 3.359704e-15, 3.356015e-15, 3.35979e-15, 
    3.357389e-15, 3.296822e-15, 3.299832e-15, 3.298206e-15, 3.301264e-15, 
    3.299109e-15, 3.308686e-15, 3.311556e-15, 3.324978e-15, 3.319474e-15, 
    3.328235e-15, 3.320365e-15, 3.32176e-15, 3.328516e-15, 3.320791e-15, 
    3.337693e-15, 3.326233e-15, 3.347512e-15, 3.336074e-15, 3.348228e-15, 
    3.346023e-15, 3.349674e-15, 3.352941e-15, 3.357052e-15, 3.364629e-15, 
    3.362875e-15, 3.369211e-15, 3.30432e-15, 3.30822e-15, 3.307879e-15, 
    3.311961e-15, 3.314979e-15, 3.32152e-15, 3.332e-15, 3.32806e-15, 
    3.335293e-15, 3.336744e-15, 3.325756e-15, 3.332502e-15, 3.310832e-15, 
    3.314333e-15, 3.31225e-15, 3.304626e-15, 3.328965e-15, 3.31648e-15, 
    3.339526e-15, 3.332771e-15, 3.352475e-15, 3.342678e-15, 3.361909e-15, 
    3.370114e-15, 3.377839e-15, 3.386848e-15, 3.310351e-15, 3.307701e-15, 
    3.312447e-15, 3.319007e-15, 3.325096e-15, 3.333183e-15, 3.334011e-15, 
    3.335525e-15, 3.339447e-15, 3.342743e-15, 3.336001e-15, 3.343569e-15, 
    3.315141e-15, 3.330049e-15, 3.306697e-15, 3.313731e-15, 3.318622e-15, 
    3.316479e-15, 3.327611e-15, 3.330232e-15, 3.340877e-15, 3.335377e-15, 
    3.368088e-15, 3.353628e-15, 3.393709e-15, 3.382523e-15, 3.306774e-15, 
    3.310343e-15, 3.322751e-15, 3.316849e-15, 3.333724e-15, 3.337873e-15, 
    3.341246e-15, 3.345553e-15, 3.34602e-15, 3.348571e-15, 3.34439e-15, 
    3.348407e-15, 3.3332e-15, 3.339999e-15, 3.321336e-15, 3.32588e-15, 
    3.32379e-15, 3.321496e-15, 3.328574e-15, 3.336107e-15, 3.336271e-15, 
    3.338685e-15, 3.345477e-15, 3.333792e-15, 3.369946e-15, 3.347628e-15, 
    3.314232e-15, 3.321096e-15, 3.32208e-15, 3.319421e-15, 3.337457e-15, 
    3.330925e-15, 3.348509e-15, 3.34376e-15, 3.351541e-15, 3.347675e-15, 
    3.347106e-15, 3.342139e-15, 3.339045e-15, 3.331224e-15, 3.324857e-15, 
    3.319807e-15, 3.320982e-15, 3.326528e-15, 3.336568e-15, 3.34606e-15, 
    3.343981e-15, 3.35095e-15, 3.332501e-15, 3.340239e-15, 3.337248e-15, 
    3.345046e-15, 3.327955e-15, 3.342501e-15, 3.324233e-15, 3.325836e-15, 
    3.330795e-15, 3.340761e-15, 3.34297e-15, 3.345322e-15, 3.343872e-15, 
    3.336824e-15, 3.33567e-15, 3.330675e-15, 3.329294e-15, 3.325488e-15, 
    3.322333e-15, 3.325214e-15, 3.328239e-15, 3.336828e-15, 3.344561e-15, 
    3.352987e-15, 3.355049e-15, 3.364875e-15, 3.356872e-15, 3.37007e-15, 
    3.358844e-15, 3.378272e-15, 3.343348e-15, 3.35852e-15, 3.331022e-15, 
    3.333988e-15, 3.339349e-15, 3.35164e-15, 3.34501e-15, 3.352765e-15, 
    3.335625e-15, 3.326718e-15, 3.324416e-15, 3.320114e-15, 3.324515e-15, 
    3.324157e-15, 3.328366e-15, 3.327014e-15, 3.337113e-15, 3.33169e-15, 
    3.347091e-15, 3.352705e-15, 3.368546e-15, 3.378242e-15, 3.388108e-15, 
    3.392459e-15, 3.393783e-15, 3.394336e-15 ;

 LITR2N_vr =
  1.532752e-05, 1.532751e-05, 1.532751e-05, 1.53275e-05, 1.532751e-05, 
    1.53275e-05, 1.532752e-05, 1.532751e-05, 1.532752e-05, 1.532752e-05, 
    1.532747e-05, 1.53275e-05, 1.532745e-05, 1.532747e-05, 1.532743e-05, 
    1.532745e-05, 1.532742e-05, 1.532743e-05, 1.532741e-05, 1.532741e-05, 
    1.532739e-05, 1.532741e-05, 1.532738e-05, 1.53274e-05, 1.532739e-05, 
    1.532741e-05, 1.532749e-05, 1.532748e-05, 1.532749e-05, 1.532749e-05, 
    1.532749e-05, 1.532751e-05, 1.532751e-05, 1.532753e-05, 1.532752e-05, 
    1.532751e-05, 1.532749e-05, 1.53275e-05, 1.532748e-05, 1.532748e-05, 
    1.532746e-05, 1.532747e-05, 1.532743e-05, 1.532744e-05, 1.532741e-05, 
    1.532742e-05, 1.532741e-05, 1.532742e-05, 1.532741e-05, 1.532742e-05, 
    1.532742e-05, 1.532743e-05, 1.532747e-05, 1.532746e-05, 1.532749e-05, 
    1.532751e-05, 1.532752e-05, 1.532753e-05, 1.532753e-05, 1.532753e-05, 
    1.532751e-05, 1.53275e-05, 1.532749e-05, 1.532749e-05, 1.532748e-05, 
    1.532746e-05, 1.532745e-05, 1.532743e-05, 1.532743e-05, 1.532743e-05, 
    1.532742e-05, 1.532741e-05, 1.532741e-05, 1.532741e-05, 1.532743e-05, 
    1.532742e-05, 1.532744e-05, 1.532743e-05, 1.532748e-05, 1.53275e-05, 
    1.53275e-05, 1.532751e-05, 1.532753e-05, 1.532752e-05, 1.532752e-05, 
    1.532751e-05, 1.53275e-05, 1.532751e-05, 1.532749e-05, 1.532749e-05, 
    1.532745e-05, 1.532747e-05, 1.532742e-05, 1.532743e-05, 1.532742e-05, 
    1.532743e-05, 1.532741e-05, 1.532743e-05, 1.532741e-05, 1.53274e-05, 
    1.53274e-05, 1.532739e-05, 1.532743e-05, 1.532741e-05, 1.532751e-05, 
    1.532751e-05, 1.53275e-05, 1.532751e-05, 1.532751e-05, 1.532753e-05, 
    1.532752e-05, 1.532751e-05, 1.53275e-05, 1.53275e-05, 1.532749e-05, 
    1.532748e-05, 1.532747e-05, 1.532745e-05, 1.532743e-05, 1.532742e-05, 
    1.532743e-05, 1.532742e-05, 1.532743e-05, 1.532743e-05, 1.53274e-05, 
    1.532742e-05, 1.53274e-05, 1.53274e-05, 1.532741e-05, 1.53274e-05, 
    1.532751e-05, 1.532751e-05, 1.532752e-05, 1.532751e-05, 1.532753e-05, 
    1.532752e-05, 1.532751e-05, 1.532749e-05, 1.532749e-05, 1.532749e-05, 
    1.532748e-05, 1.532747e-05, 1.532745e-05, 1.532744e-05, 1.532742e-05, 
    1.532742e-05, 1.532742e-05, 1.532742e-05, 1.532743e-05, 1.532742e-05, 
    1.532742e-05, 1.532742e-05, 1.53274e-05, 1.53274e-05, 1.53274e-05, 
    1.53274e-05, 1.532751e-05, 1.53275e-05, 1.532751e-05, 1.53275e-05, 
    1.53275e-05, 1.532749e-05, 1.532748e-05, 1.532746e-05, 1.532747e-05, 
    1.532745e-05, 1.532747e-05, 1.532746e-05, 1.532745e-05, 1.532747e-05, 
    1.532744e-05, 1.532746e-05, 1.532742e-05, 1.532744e-05, 1.532742e-05, 
    1.532742e-05, 1.532742e-05, 1.532741e-05, 1.53274e-05, 1.532739e-05, 
    1.532739e-05, 1.532738e-05, 1.532749e-05, 1.532749e-05, 1.532749e-05, 
    1.532748e-05, 1.532748e-05, 1.532747e-05, 1.532745e-05, 1.532745e-05, 
    1.532744e-05, 1.532744e-05, 1.532746e-05, 1.532744e-05, 1.532748e-05, 
    1.532748e-05, 1.532748e-05, 1.532749e-05, 1.532745e-05, 1.532747e-05, 
    1.532743e-05, 1.532744e-05, 1.532741e-05, 1.532743e-05, 1.532739e-05, 
    1.532738e-05, 1.532737e-05, 1.532735e-05, 1.532748e-05, 1.532749e-05, 
    1.532748e-05, 1.532747e-05, 1.532746e-05, 1.532744e-05, 1.532744e-05, 
    1.532744e-05, 1.532743e-05, 1.532743e-05, 1.532744e-05, 1.532743e-05, 
    1.532748e-05, 1.532745e-05, 1.532749e-05, 1.532748e-05, 1.532747e-05, 
    1.532747e-05, 1.532745e-05, 1.532745e-05, 1.532743e-05, 1.532744e-05, 
    1.532738e-05, 1.532741e-05, 1.532734e-05, 1.532736e-05, 1.532749e-05, 
    1.532748e-05, 1.532746e-05, 1.532747e-05, 1.532744e-05, 1.532744e-05, 
    1.532743e-05, 1.532742e-05, 1.532742e-05, 1.532742e-05, 1.532742e-05, 
    1.532742e-05, 1.532744e-05, 1.532743e-05, 1.532747e-05, 1.532746e-05, 
    1.532746e-05, 1.532747e-05, 1.532745e-05, 1.532744e-05, 1.532744e-05, 
    1.532743e-05, 1.532742e-05, 1.532744e-05, 1.532738e-05, 1.532742e-05, 
    1.532748e-05, 1.532747e-05, 1.532746e-05, 1.532747e-05, 1.532744e-05, 
    1.532745e-05, 1.532742e-05, 1.532742e-05, 1.532741e-05, 1.532742e-05, 
    1.532742e-05, 1.532743e-05, 1.532743e-05, 1.532745e-05, 1.532746e-05, 
    1.532747e-05, 1.532747e-05, 1.532746e-05, 1.532744e-05, 1.532742e-05, 
    1.532742e-05, 1.532741e-05, 1.532744e-05, 1.532743e-05, 1.532744e-05, 
    1.532742e-05, 1.532745e-05, 1.532743e-05, 1.532746e-05, 1.532746e-05, 
    1.532745e-05, 1.532743e-05, 1.532743e-05, 1.532742e-05, 1.532742e-05, 
    1.532744e-05, 1.532744e-05, 1.532745e-05, 1.532745e-05, 1.532746e-05, 
    1.532746e-05, 1.532746e-05, 1.532745e-05, 1.532744e-05, 1.532742e-05, 
    1.532741e-05, 1.532741e-05, 1.532739e-05, 1.53274e-05, 1.532738e-05, 
    1.53274e-05, 1.532736e-05, 1.532743e-05, 1.53274e-05, 1.532745e-05, 
    1.532744e-05, 1.532743e-05, 1.532741e-05, 1.532742e-05, 1.532741e-05, 
    1.532744e-05, 1.532746e-05, 1.532746e-05, 1.532747e-05, 1.532746e-05, 
    1.532746e-05, 1.532745e-05, 1.532745e-05, 1.532744e-05, 1.532745e-05, 
    1.532742e-05, 1.532741e-05, 1.532738e-05, 1.532736e-05, 1.532735e-05, 
    1.532734e-05, 1.532734e-05, 1.532734e-05,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR2_HR =
  1.187703e-13, 1.190959e-13, 1.190327e-13, 1.192951e-13, 1.191496e-13, 
    1.193214e-13, 1.188364e-13, 1.191088e-13, 1.189349e-13, 1.187997e-13, 
    1.198038e-13, 1.193068e-13, 1.203199e-13, 1.200033e-13, 1.207983e-13, 
    1.202706e-13, 1.209046e-13, 1.207832e-13, 1.211488e-13, 1.210441e-13, 
    1.215111e-13, 1.211971e-13, 1.217532e-13, 1.214362e-13, 1.214858e-13, 
    1.211867e-13, 1.19407e-13, 1.197419e-13, 1.193871e-13, 1.194349e-13, 
    1.194135e-13, 1.191525e-13, 1.190209e-13, 1.187455e-13, 1.187955e-13, 
    1.189978e-13, 1.194564e-13, 1.193009e-13, 1.196929e-13, 1.196841e-13, 
    1.201201e-13, 1.199236e-13, 1.206558e-13, 1.204478e-13, 1.210485e-13, 
    1.208975e-13, 1.210414e-13, 1.209978e-13, 1.210419e-13, 1.208205e-13, 
    1.209154e-13, 1.207205e-13, 1.199604e-13, 1.201839e-13, 1.195168e-13, 
    1.191151e-13, 1.188483e-13, 1.186588e-13, 1.186856e-13, 1.187366e-13, 
    1.18999e-13, 1.192457e-13, 1.194335e-13, 1.195591e-13, 1.196828e-13, 
    1.200568e-13, 1.202548e-13, 1.206977e-13, 1.206179e-13, 1.207532e-13, 
    1.208825e-13, 1.210993e-13, 1.210636e-13, 1.211591e-13, 1.207497e-13, 
    1.210218e-13, 1.205724e-13, 1.206954e-13, 1.19716e-13, 1.193428e-13, 
    1.191838e-13, 1.190448e-13, 1.187062e-13, 1.1894e-13, 1.188479e-13, 
    1.190672e-13, 1.192065e-13, 1.191376e-13, 1.195625e-13, 1.193974e-13, 
    1.202666e-13, 1.198924e-13, 1.208674e-13, 1.206343e-13, 1.209233e-13, 
    1.207759e-13, 1.210283e-13, 1.208011e-13, 1.211947e-13, 1.212803e-13, 
    1.212218e-13, 1.214466e-13, 1.207885e-13, 1.210413e-13, 1.191357e-13, 
    1.191469e-13, 1.191992e-13, 1.189691e-13, 1.18955e-13, 1.187441e-13, 
    1.189318e-13, 1.190117e-13, 1.192146e-13, 1.193345e-13, 1.194484e-13, 
    1.196989e-13, 1.199784e-13, 1.20369e-13, 1.206494e-13, 1.208373e-13, 
    1.207221e-13, 1.208238e-13, 1.207101e-13, 1.206569e-13, 1.212482e-13, 
    1.209162e-13, 1.214143e-13, 1.213867e-13, 1.211614e-13, 1.213898e-13, 
    1.191548e-13, 1.190901e-13, 1.188656e-13, 1.190413e-13, 1.187211e-13, 
    1.189003e-13, 1.190033e-13, 1.194007e-13, 1.194881e-13, 1.19569e-13, 
    1.197287e-13, 1.199336e-13, 1.202928e-13, 1.206051e-13, 1.2089e-13, 
    1.208691e-13, 1.208765e-13, 1.209401e-13, 1.207825e-13, 1.209659e-13, 
    1.209967e-13, 1.209162e-13, 1.21383e-13, 1.212497e-13, 1.213862e-13, 
    1.212994e-13, 1.191112e-13, 1.192199e-13, 1.191612e-13, 1.192716e-13, 
    1.191938e-13, 1.195398e-13, 1.196435e-13, 1.201284e-13, 1.199296e-13, 
    1.202461e-13, 1.199618e-13, 1.200121e-13, 1.202563e-13, 1.199772e-13, 
    1.205878e-13, 1.201738e-13, 1.209425e-13, 1.205293e-13, 1.209684e-13, 
    1.208888e-13, 1.210207e-13, 1.211387e-13, 1.212872e-13, 1.21561e-13, 
    1.214976e-13, 1.217265e-13, 1.19382e-13, 1.19523e-13, 1.195106e-13, 
    1.196581e-13, 1.197672e-13, 1.200035e-13, 1.203821e-13, 1.202398e-13, 
    1.205011e-13, 1.205535e-13, 1.201565e-13, 1.204002e-13, 1.196173e-13, 
    1.197438e-13, 1.196686e-13, 1.193931e-13, 1.202725e-13, 1.198214e-13, 
    1.20654e-13, 1.2041e-13, 1.211219e-13, 1.207679e-13, 1.214627e-13, 
    1.217591e-13, 1.220382e-13, 1.223637e-13, 1.196e-13, 1.195042e-13, 
    1.196757e-13, 1.199127e-13, 1.201327e-13, 1.204249e-13, 1.204548e-13, 
    1.205095e-13, 1.206512e-13, 1.207702e-13, 1.205267e-13, 1.208001e-13, 
    1.19773e-13, 1.203117e-13, 1.194679e-13, 1.197221e-13, 1.198988e-13, 
    1.198213e-13, 1.202235e-13, 1.203182e-13, 1.207028e-13, 1.205041e-13, 
    1.216859e-13, 1.211635e-13, 1.226116e-13, 1.222075e-13, 1.194707e-13, 
    1.195997e-13, 1.200479e-13, 1.198347e-13, 1.204444e-13, 1.205943e-13, 
    1.207162e-13, 1.208718e-13, 1.208886e-13, 1.209808e-13, 1.208297e-13, 
    1.209749e-13, 1.204255e-13, 1.206711e-13, 1.199968e-13, 1.20161e-13, 
    1.200855e-13, 1.200026e-13, 1.202583e-13, 1.205305e-13, 1.205364e-13, 
    1.206236e-13, 1.20869e-13, 1.204469e-13, 1.217531e-13, 1.209467e-13, 
    1.197402e-13, 1.199882e-13, 1.200237e-13, 1.199277e-13, 1.205793e-13, 
    1.203433e-13, 1.209786e-13, 1.20807e-13, 1.210881e-13, 1.209484e-13, 
    1.209279e-13, 1.207484e-13, 1.206366e-13, 1.203541e-13, 1.20124e-13, 
    1.199416e-13, 1.19984e-13, 1.201844e-13, 1.205472e-13, 1.208901e-13, 
    1.20815e-13, 1.210668e-13, 1.204002e-13, 1.206798e-13, 1.205717e-13, 
    1.208535e-13, 1.20236e-13, 1.207615e-13, 1.201015e-13, 1.201594e-13, 
    1.203386e-13, 1.206987e-13, 1.207785e-13, 1.208634e-13, 1.20811e-13, 
    1.205564e-13, 1.205147e-13, 1.203343e-13, 1.202844e-13, 1.201468e-13, 
    1.200329e-13, 1.20137e-13, 1.202462e-13, 1.205565e-13, 1.208359e-13, 
    1.211403e-13, 1.212149e-13, 1.215699e-13, 1.212807e-13, 1.217575e-13, 
    1.21352e-13, 1.220539e-13, 1.207921e-13, 1.213403e-13, 1.203468e-13, 
    1.20454e-13, 1.206476e-13, 1.210917e-13, 1.208521e-13, 1.211323e-13, 
    1.205131e-13, 1.201913e-13, 1.201081e-13, 1.199527e-13, 1.201117e-13, 
    1.200988e-13, 1.202508e-13, 1.20202e-13, 1.205668e-13, 1.203709e-13, 
    1.209273e-13, 1.211302e-13, 1.217025e-13, 1.220528e-13, 1.224093e-13, 
    1.225664e-13, 1.226143e-13, 1.226343e-13 ;

 LITR3C =
  9.69806e-06, 9.69805e-06, 9.698052e-06, 9.698045e-06, 9.698048e-06, 
    9.698044e-06, 9.698058e-06, 9.69805e-06, 9.698056e-06, 9.698059e-06, 
    9.698029e-06, 9.698044e-06, 9.698013e-06, 9.698023e-06, 9.697998e-06, 
    9.698015e-06, 9.697996e-06, 9.697999e-06, 9.697988e-06, 9.697991e-06, 
    9.697977e-06, 9.697987e-06, 9.697969e-06, 9.697979e-06, 9.697977e-06, 
    9.697987e-06, 9.698041e-06, 9.698031e-06, 9.698042e-06, 9.69804e-06, 
    9.698041e-06, 9.698048e-06, 9.698053e-06, 9.698061e-06, 9.698059e-06, 
    9.698054e-06, 9.698039e-06, 9.698044e-06, 9.698032e-06, 9.698033e-06, 
    9.698019e-06, 9.698026e-06, 9.698003e-06, 9.698009e-06, 9.697991e-06, 
    9.697996e-06, 9.697991e-06, 9.697993e-06, 9.697991e-06, 9.697998e-06, 
    9.697995e-06, 9.698001e-06, 9.698024e-06, 9.698017e-06, 9.698038e-06, 
    9.69805e-06, 9.698058e-06, 9.698064e-06, 9.698063e-06, 9.698061e-06, 
    9.698054e-06, 9.698046e-06, 9.69804e-06, 9.698037e-06, 9.698033e-06, 
    9.698021e-06, 9.698015e-06, 9.698002e-06, 9.698004e-06, 9.698e-06, 
    9.697996e-06, 9.697989e-06, 9.69799e-06, 9.697987e-06, 9.698e-06, 
    9.697992e-06, 9.698006e-06, 9.698002e-06, 9.698032e-06, 9.698043e-06, 
    9.698048e-06, 9.698052e-06, 9.698062e-06, 9.698055e-06, 9.698058e-06, 
    9.698051e-06, 9.698048e-06, 9.698049e-06, 9.698037e-06, 9.698041e-06, 
    9.698015e-06, 9.698027e-06, 9.697997e-06, 9.698004e-06, 9.697995e-06, 
    9.697999e-06, 9.697992e-06, 9.697998e-06, 9.697987e-06, 9.697984e-06, 
    9.697986e-06, 9.697979e-06, 9.697999e-06, 9.697991e-06, 9.698049e-06, 
    9.698049e-06, 9.698048e-06, 9.698055e-06, 9.698055e-06, 9.698061e-06, 
    9.698056e-06, 9.698053e-06, 9.698047e-06, 9.698043e-06, 9.698039e-06, 
    9.698032e-06, 9.698024e-06, 9.698012e-06, 9.698003e-06, 9.697997e-06, 
    9.698001e-06, 9.697997e-06, 9.698001e-06, 9.698003e-06, 9.697985e-06, 
    9.697995e-06, 9.69798e-06, 9.697981e-06, 9.697987e-06, 9.69798e-06, 
    9.698048e-06, 9.69805e-06, 9.698058e-06, 9.698052e-06, 9.698062e-06, 
    9.698057e-06, 9.698053e-06, 9.698041e-06, 9.698038e-06, 9.698036e-06, 
    9.698031e-06, 9.698025e-06, 9.698014e-06, 9.698005e-06, 9.697996e-06, 
    9.697997e-06, 9.697997e-06, 9.697995e-06, 9.697999e-06, 9.697994e-06, 
    9.697993e-06, 9.697995e-06, 9.697981e-06, 9.697985e-06, 9.697981e-06, 
    9.697983e-06, 9.69805e-06, 9.698047e-06, 9.698048e-06, 9.698045e-06, 
    9.698048e-06, 9.698037e-06, 9.698034e-06, 9.698019e-06, 9.698025e-06, 
    9.698016e-06, 9.698024e-06, 9.698023e-06, 9.698015e-06, 9.698024e-06, 
    9.698005e-06, 9.698017e-06, 9.697994e-06, 9.698007e-06, 9.697994e-06, 
    9.697996e-06, 9.697992e-06, 9.697988e-06, 9.697984e-06, 9.697976e-06, 
    9.697977e-06, 9.69797e-06, 9.698042e-06, 9.698038e-06, 9.698038e-06, 
    9.698033e-06, 9.69803e-06, 9.698023e-06, 9.698011e-06, 9.698016e-06, 
    9.698007e-06, 9.698006e-06, 9.698018e-06, 9.698011e-06, 9.698035e-06, 
    9.698031e-06, 9.698033e-06, 9.698041e-06, 9.698015e-06, 9.698028e-06, 
    9.698003e-06, 9.69801e-06, 9.697988e-06, 9.697999e-06, 9.697978e-06, 
    9.697969e-06, 9.697961e-06, 9.697951e-06, 9.698035e-06, 9.698038e-06, 
    9.698033e-06, 9.698026e-06, 9.698019e-06, 9.69801e-06, 9.698009e-06, 
    9.698007e-06, 9.698003e-06, 9.697999e-06, 9.698007e-06, 9.697998e-06, 
    9.69803e-06, 9.698014e-06, 9.698039e-06, 9.698031e-06, 9.698026e-06, 
    9.698028e-06, 9.698017e-06, 9.698013e-06, 9.698001e-06, 9.698007e-06, 
    9.697972e-06, 9.697987e-06, 9.697944e-06, 9.697956e-06, 9.698039e-06, 
    9.698035e-06, 9.698021e-06, 9.698028e-06, 9.698009e-06, 9.698005e-06, 
    9.698001e-06, 9.697997e-06, 9.697996e-06, 9.697993e-06, 9.697997e-06, 
    9.697993e-06, 9.69801e-06, 9.698003e-06, 9.698023e-06, 9.698018e-06, 
    9.69802e-06, 9.698023e-06, 9.698015e-06, 9.698007e-06, 9.698007e-06, 
    9.698004e-06, 9.697997e-06, 9.698009e-06, 9.697969e-06, 9.697994e-06, 
    9.698031e-06, 9.698023e-06, 9.698022e-06, 9.698025e-06, 9.698006e-06, 
    9.698013e-06, 9.697993e-06, 9.697998e-06, 9.69799e-06, 9.697994e-06, 
    9.697995e-06, 9.698e-06, 9.698004e-06, 9.698012e-06, 9.698019e-06, 
    9.698025e-06, 9.698024e-06, 9.698017e-06, 9.698007e-06, 9.697996e-06, 
    9.697998e-06, 9.69799e-06, 9.698011e-06, 9.698002e-06, 9.698006e-06, 
    9.697997e-06, 9.698016e-06, 9.698e-06, 9.69802e-06, 9.698018e-06, 
    9.698013e-06, 9.698002e-06, 9.697999e-06, 9.697997e-06, 9.697998e-06, 
    9.698006e-06, 9.698007e-06, 9.698013e-06, 9.698014e-06, 9.698018e-06, 
    9.698022e-06, 9.698018e-06, 9.698016e-06, 9.698006e-06, 9.697997e-06, 
    9.697988e-06, 9.697986e-06, 9.697975e-06, 9.697984e-06, 9.697969e-06, 
    9.697982e-06, 9.69796e-06, 9.697998e-06, 9.697982e-06, 9.698012e-06, 
    9.698009e-06, 9.698003e-06, 9.697989e-06, 9.697997e-06, 9.697988e-06, 
    9.698007e-06, 9.698017e-06, 9.698019e-06, 9.698025e-06, 9.698019e-06, 
    9.69802e-06, 9.698016e-06, 9.698017e-06, 9.698006e-06, 9.698012e-06, 
    9.697995e-06, 9.697988e-06, 9.697971e-06, 9.69796e-06, 9.697949e-06, 
    9.697945e-06, 9.697943e-06, 9.697943e-06 ;

 LITR3C_TO_SOIL2C =
  5.938512e-14, 5.954794e-14, 5.951631e-14, 5.964753e-14, 5.957477e-14, 
    5.966066e-14, 5.941816e-14, 5.955438e-14, 5.946745e-14, 5.939982e-14, 
    5.990189e-14, 5.965339e-14, 6.015994e-14, 6.000165e-14, 6.039911e-14, 
    6.013528e-14, 6.045228e-14, 6.039157e-14, 6.057439e-14, 6.052204e-14, 
    6.075555e-14, 6.059855e-14, 6.087658e-14, 6.07181e-14, 6.074287e-14, 
    6.059336e-14, 5.970348e-14, 5.987095e-14, 5.969354e-14, 5.971744e-14, 
    5.970673e-14, 5.957625e-14, 5.951043e-14, 5.937271e-14, 5.939773e-14, 
    5.949891e-14, 5.972818e-14, 5.965042e-14, 5.984646e-14, 5.984203e-14, 
    6.006002e-14, 5.996177e-14, 6.032785e-14, 6.022389e-14, 6.052422e-14, 
    6.044872e-14, 6.052067e-14, 6.049886e-14, 6.052095e-14, 6.041022e-14, 
    6.045767e-14, 6.036022e-14, 5.998016e-14, 6.009191e-14, 5.97584e-14, 
    5.955752e-14, 5.942413e-14, 5.932939e-14, 5.934278e-14, 5.936831e-14, 
    5.94995e-14, 5.962283e-14, 5.971674e-14, 5.977953e-14, 5.984139e-14, 
    6.002837e-14, 6.012739e-14, 6.034884e-14, 6.030895e-14, 6.037657e-14, 
    6.044122e-14, 6.054964e-14, 6.053181e-14, 6.057955e-14, 6.037482e-14, 
    6.051089e-14, 6.028621e-14, 6.034768e-14, 5.985801e-14, 5.967141e-14, 
    5.959187e-14, 5.952238e-14, 5.935308e-14, 5.947e-14, 5.942391e-14, 
    5.953358e-14, 5.960321e-14, 5.956879e-14, 5.978125e-14, 5.969867e-14, 
    6.013326e-14, 5.994618e-14, 6.043368e-14, 6.031714e-14, 6.04616e-14, 
    6.038791e-14, 6.051415e-14, 6.040054e-14, 6.059733e-14, 6.064013e-14, 
    6.061087e-14, 6.072328e-14, 6.039424e-14, 6.052065e-14, 5.956782e-14, 
    5.957343e-14, 5.95996e-14, 5.948452e-14, 5.947748e-14, 5.937202e-14, 
    5.946588e-14, 5.950582e-14, 5.960727e-14, 5.966721e-14, 5.972419e-14, 
    5.984943e-14, 5.998917e-14, 6.018447e-14, 6.03247e-14, 6.041862e-14, 
    6.036105e-14, 6.041188e-14, 6.035505e-14, 6.032841e-14, 6.062408e-14, 
    6.045809e-14, 6.070712e-14, 6.069335e-14, 6.058067e-14, 6.06949e-14, 
    5.957737e-14, 5.954506e-14, 5.943276e-14, 5.952065e-14, 5.936053e-14, 
    5.945015e-14, 5.950165e-14, 5.970035e-14, 5.974403e-14, 5.978447e-14, 
    5.986434e-14, 5.99668e-14, 6.014637e-14, 6.030252e-14, 6.044498e-14, 
    6.043455e-14, 6.043823e-14, 6.047001e-14, 6.039123e-14, 6.048295e-14, 
    6.049832e-14, 6.04581e-14, 6.069151e-14, 6.062486e-14, 6.069306e-14, 
    6.064967e-14, 5.955557e-14, 5.960994e-14, 5.958056e-14, 5.96358e-14, 
    5.959687e-14, 5.976988e-14, 5.982172e-14, 6.006419e-14, 5.996477e-14, 
    6.012304e-14, 5.998086e-14, 6.000605e-14, 6.012811e-14, 5.998856e-14, 
    6.029387e-14, 6.008686e-14, 6.047125e-14, 6.026463e-14, 6.048419e-14, 
    6.044437e-14, 6.051031e-14, 6.056933e-14, 6.064359e-14, 6.078047e-14, 
    6.074879e-14, 6.086323e-14, 5.969101e-14, 5.976147e-14, 5.97553e-14, 
    5.982905e-14, 5.988356e-14, 6.000172e-14, 6.019104e-14, 6.011988e-14, 
    6.025053e-14, 6.027673e-14, 6.007825e-14, 6.020011e-14, 5.980864e-14, 
    5.98719e-14, 5.983427e-14, 5.969654e-14, 6.013622e-14, 5.991067e-14, 
    6.0327e-14, 6.020497e-14, 6.056091e-14, 6.038394e-14, 6.073134e-14, 
    6.087955e-14, 6.101911e-14, 6.118185e-14, 5.979996e-14, 5.975209e-14, 
    5.983783e-14, 5.995633e-14, 6.006633e-14, 6.021241e-14, 6.022737e-14, 
    6.025471e-14, 6.032556e-14, 6.03851e-14, 6.026332e-14, 6.040002e-14, 
    5.98865e-14, 6.015581e-14, 5.973395e-14, 5.986102e-14, 5.994937e-14, 
    5.991065e-14, 6.011175e-14, 6.015911e-14, 6.03514e-14, 6.025204e-14, 
    6.084295e-14, 6.058174e-14, 6.130578e-14, 6.110372e-14, 5.973535e-14, 
    5.979981e-14, 6.002395e-14, 5.991734e-14, 6.022218e-14, 6.029712e-14, 
    6.035806e-14, 6.043587e-14, 6.04443e-14, 6.049038e-14, 6.041485e-14, 
    6.048742e-14, 6.021272e-14, 6.033553e-14, 5.999839e-14, 6.008048e-14, 
    6.004273e-14, 6.000129e-14, 6.012916e-14, 6.026523e-14, 6.02682e-14, 
    6.03118e-14, 6.04345e-14, 6.022341e-14, 6.087652e-14, 6.047334e-14, 
    5.987008e-14, 5.999406e-14, 6.001184e-14, 5.996381e-14, 6.028961e-14, 
    6.017161e-14, 6.048927e-14, 6.040348e-14, 6.054404e-14, 6.04742e-14, 
    6.046392e-14, 6.03742e-14, 6.03183e-14, 6.017702e-14, 6.0062e-14, 
    5.997079e-14, 5.9992e-14, 6.00922e-14, 6.027356e-14, 6.044503e-14, 
    6.040748e-14, 6.053336e-14, 6.020009e-14, 6.033988e-14, 6.028584e-14, 
    6.042671e-14, 6.011797e-14, 6.038073e-14, 6.005073e-14, 6.007969e-14, 
    6.016928e-14, 6.034932e-14, 6.038921e-14, 6.043169e-14, 6.04055e-14, 
    6.027818e-14, 6.025734e-14, 6.016712e-14, 6.014216e-14, 6.007339e-14, 
    6.001642e-14, 6.006846e-14, 6.012309e-14, 6.027826e-14, 6.041795e-14, 
    6.057016e-14, 6.060742e-14, 6.078491e-14, 6.064035e-14, 6.087875e-14, 
    6.067596e-14, 6.102693e-14, 6.039604e-14, 6.067012e-14, 6.017337e-14, 
    6.022696e-14, 6.032379e-14, 6.054583e-14, 6.042606e-14, 6.056615e-14, 
    6.025653e-14, 6.009562e-14, 6.005404e-14, 5.997632e-14, 6.005582e-14, 
    6.004936e-14, 6.012539e-14, 6.010097e-14, 6.028341e-14, 6.018543e-14, 
    6.046365e-14, 6.056506e-14, 6.085122e-14, 6.102639e-14, 6.120461e-14, 
    6.12832e-14, 6.130712e-14, 6.131711e-14 ;

 LITR3C_vr =
  0.0005537693, 0.0005537687, 0.0005537688, 0.0005537684, 0.0005537686, 
    0.0005537683, 0.0005537692, 0.0005537687, 0.000553769, 0.0005537692, 
    0.0005537675, 0.0005537684, 0.0005537666, 0.0005537671, 0.0005537657, 
    0.0005537667, 0.0005537656, 0.0005537657, 0.0005537652, 0.0005537653, 
    0.0005537645, 0.000553765, 0.0005537641, 0.0005537646, 0.0005537646, 
    0.000553765, 0.0005537682, 0.0005537676, 0.0005537682, 0.0005537681, 
    0.0005537681, 0.0005537686, 0.0005537688, 0.0005537693, 0.0005537692, 
    0.0005537689, 0.0005537681, 0.0005537684, 0.0005537677, 0.0005537677, 
    0.0005537669, 0.0005537673, 0.000553766, 0.0005537664, 0.0005537653, 
    0.0005537656, 0.0005537653, 0.0005537654, 0.0005537653, 0.0005537657, 
    0.0005537656, 0.0005537659, 0.0005537672, 0.0005537668, 0.000553768, 
    0.0005537687, 0.0005537691, 0.0005537695, 0.0005537694, 0.0005537694, 
    0.0005537689, 0.0005537684, 0.0005537681, 0.0005537679, 0.0005537677, 
    0.000553767, 0.0005537667, 0.0005537659, 0.000553766, 0.0005537658, 
    0.0005537656, 0.0005537652, 0.0005537653, 0.0005537651, 0.0005537658, 
    0.0005537653, 0.0005537661, 0.0005537659, 0.0005537676, 0.0005537683, 
    0.0005537685, 0.0005537688, 0.0005537694, 0.000553769, 0.0005537691, 
    0.0005537688, 0.0005537685, 0.0005537687, 0.0005537679, 0.0005537682, 
    0.0005537667, 0.0005537673, 0.0005537656, 0.000553766, 0.0005537655, 
    0.0005537658, 0.0005537653, 0.0005537657, 0.000553765, 0.0005537649, 
    0.000553765, 0.0005537646, 0.0005537657, 0.0005537653, 0.0005537687, 
    0.0005537686, 0.0005537685, 0.0005537689, 0.0005537689, 0.0005537693, 
    0.000553769, 0.0005537688, 0.0005537685, 0.0005537683, 0.0005537681, 
    0.0005537677, 0.0005537672, 0.0005537665, 0.000553766, 0.0005537657, 
    0.0005537659, 0.0005537657, 0.0005537659, 0.000553766, 0.000553765, 
    0.0005537656, 0.0005537647, 0.0005537647, 0.0005537651, 0.0005537647, 
    0.0005537686, 0.0005537687, 0.0005537691, 0.0005537688, 0.0005537694, 
    0.0005537691, 0.0005537689, 0.0005537682, 0.000553768, 0.0005537679, 
    0.0005537676, 0.0005537673, 0.0005537666, 0.0005537661, 0.0005537656, 
    0.0005537656, 0.0005537656, 0.0005537655, 0.0005537658, 0.0005537655, 
    0.0005537654, 0.0005537656, 0.0005537648, 0.000553765, 0.0005537647, 
    0.0005537649, 0.0005537687, 0.0005537685, 0.0005537686, 0.0005537684, 
    0.0005537685, 0.000553768, 0.0005537678, 0.0005537669, 0.0005537673, 
    0.0005537667, 0.0005537672, 0.0005537671, 0.0005537667, 0.0005537672, 
    0.0005537661, 0.0005537668, 0.0005537655, 0.0005537662, 0.0005537655, 
    0.0005537656, 0.0005537653, 0.0005537652, 0.0005537649, 0.0005537644, 
    0.0005537645, 0.0005537641, 0.0005537682, 0.000553768, 0.000553768, 
    0.0005537677, 0.0005537675, 0.0005537671, 0.0005537664, 0.0005537667, 
    0.0005537663, 0.0005537661, 0.0005537668, 0.0005537664, 0.0005537678, 
    0.0005537676, 0.0005537677, 0.0005537682, 0.0005537667, 0.0005537674, 
    0.000553766, 0.0005537664, 0.0005537652, 0.0005537658, 0.0005537646, 
    0.0005537641, 0.0005537636, 0.000553763, 0.0005537678, 0.000553768, 
    0.0005537677, 0.0005537673, 0.0005537669, 0.0005537664, 0.0005537663, 
    0.0005537663, 0.000553766, 0.0005537658, 0.0005537662, 0.0005537657, 
    0.0005537675, 0.0005537666, 0.0005537681, 0.0005537676, 0.0005537673, 
    0.0005537674, 0.0005537667, 0.0005537666, 0.0005537659, 0.0005537663, 
    0.0005537642, 0.0005537651, 0.0005537626, 0.0005537633, 0.0005537681, 
    0.0005537678, 0.000553767, 0.0005537674, 0.0005537664, 0.0005537661, 
    0.0005537659, 0.0005537656, 0.0005537656, 0.0005537655, 0.0005537657, 
    0.0005537655, 0.0005537664, 0.000553766, 0.0005537671, 0.0005537668, 
    0.000553767, 0.0005537671, 0.0005537667, 0.0005537662, 0.0005537662, 
    0.000553766, 0.0005537656, 0.0005537664, 0.0005537641, 0.0005537655, 
    0.0005537676, 0.0005537671, 0.0005537671, 0.0005537673, 0.0005537661, 
    0.0005537666, 0.0005537655, 0.0005537657, 0.0005537652, 0.0005537655, 
    0.0005537655, 0.0005537659, 0.000553766, 0.0005537665, 0.0005537669, 
    0.0005537673, 0.0005537671, 0.0005537668, 0.0005537662, 0.0005537656, 
    0.0005537657, 0.0005537653, 0.0005537664, 0.000553766, 0.0005537661, 
    0.0005537656, 0.0005537667, 0.0005537658, 0.000553767, 0.0005537668, 
    0.0005537666, 0.0005537659, 0.0005537658, 0.0005537656, 0.0005537657, 
    0.0005537661, 0.0005537663, 0.0005537666, 0.0005537666, 0.0005537669, 
    0.0005537671, 0.0005537669, 0.0005537667, 0.0005537661, 0.0005537657, 
    0.0005537652, 0.000553765, 0.0005537644, 0.0005537649, 0.0005537641, 
    0.0005537648, 0.0005537636, 0.0005537657, 0.0005537648, 0.0005537666, 
    0.0005537663, 0.000553766, 0.0005537652, 0.0005537656, 0.0005537652, 
    0.0005537663, 0.0005537668, 0.000553767, 0.0005537672, 0.000553767, 
    0.000553767, 0.0005537667, 0.0005537668, 0.0005537661, 0.0005537665, 
    0.0005537655, 0.0005537652, 0.0005537642, 0.0005537636, 0.0005537629, 
    0.0005537627, 0.0005537626, 0.0005537625,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N =
  1.342141e-07, 1.342139e-07, 1.342139e-07, 1.342138e-07, 1.342139e-07, 
    1.342138e-07, 1.34214e-07, 1.342139e-07, 1.34214e-07, 1.34214e-07, 
    1.342136e-07, 1.342138e-07, 1.342134e-07, 1.342135e-07, 1.342132e-07, 
    1.342134e-07, 1.342132e-07, 1.342132e-07, 1.342131e-07, 1.342131e-07, 
    1.342129e-07, 1.34213e-07, 1.342128e-07, 1.342129e-07, 1.342129e-07, 
    1.34213e-07, 1.342138e-07, 1.342136e-07, 1.342138e-07, 1.342138e-07, 
    1.342138e-07, 1.342139e-07, 1.342139e-07, 1.342141e-07, 1.34214e-07, 
    1.34214e-07, 1.342138e-07, 1.342138e-07, 1.342137e-07, 1.342137e-07, 
    1.342135e-07, 1.342136e-07, 1.342133e-07, 1.342134e-07, 1.342131e-07, 
    1.342132e-07, 1.342131e-07, 1.342131e-07, 1.342131e-07, 1.342132e-07, 
    1.342132e-07, 1.342132e-07, 1.342136e-07, 1.342135e-07, 1.342137e-07, 
    1.342139e-07, 1.34214e-07, 1.342141e-07, 1.342141e-07, 1.342141e-07, 
    1.34214e-07, 1.342139e-07, 1.342138e-07, 1.342137e-07, 1.342137e-07, 
    1.342135e-07, 1.342134e-07, 1.342133e-07, 1.342133e-07, 1.342132e-07, 
    1.342132e-07, 1.342131e-07, 1.342131e-07, 1.342131e-07, 1.342132e-07, 
    1.342131e-07, 1.342133e-07, 1.342133e-07, 1.342137e-07, 1.342138e-07, 
    1.342139e-07, 1.342139e-07, 1.342141e-07, 1.34214e-07, 1.34214e-07, 
    1.342139e-07, 1.342139e-07, 1.342139e-07, 1.342137e-07, 1.342138e-07, 
    1.342134e-07, 1.342136e-07, 1.342132e-07, 1.342133e-07, 1.342132e-07, 
    1.342132e-07, 1.342131e-07, 1.342132e-07, 1.34213e-07, 1.34213e-07, 
    1.34213e-07, 1.342129e-07, 1.342132e-07, 1.342131e-07, 1.342139e-07, 
    1.342139e-07, 1.342139e-07, 1.34214e-07, 1.34214e-07, 1.342141e-07, 
    1.34214e-07, 1.34214e-07, 1.342139e-07, 1.342138e-07, 1.342138e-07, 
    1.342137e-07, 1.342136e-07, 1.342134e-07, 1.342133e-07, 1.342132e-07, 
    1.342132e-07, 1.342132e-07, 1.342132e-07, 1.342133e-07, 1.34213e-07, 
    1.342132e-07, 1.342129e-07, 1.34213e-07, 1.342131e-07, 1.34213e-07, 
    1.342139e-07, 1.342139e-07, 1.34214e-07, 1.342139e-07, 1.342141e-07, 
    1.34214e-07, 1.34214e-07, 1.342138e-07, 1.342138e-07, 1.342137e-07, 
    1.342136e-07, 1.342136e-07, 1.342134e-07, 1.342133e-07, 1.342132e-07, 
    1.342132e-07, 1.342132e-07, 1.342131e-07, 1.342132e-07, 1.342131e-07, 
    1.342131e-07, 1.342132e-07, 1.34213e-07, 1.34213e-07, 1.34213e-07, 
    1.34213e-07, 1.342139e-07, 1.342139e-07, 1.342139e-07, 1.342138e-07, 
    1.342139e-07, 1.342137e-07, 1.342137e-07, 1.342135e-07, 1.342136e-07, 
    1.342134e-07, 1.342136e-07, 1.342135e-07, 1.342134e-07, 1.342136e-07, 
    1.342133e-07, 1.342135e-07, 1.342131e-07, 1.342133e-07, 1.342131e-07, 
    1.342132e-07, 1.342131e-07, 1.342131e-07, 1.34213e-07, 1.342129e-07, 
    1.342129e-07, 1.342128e-07, 1.342138e-07, 1.342137e-07, 1.342137e-07, 
    1.342137e-07, 1.342136e-07, 1.342135e-07, 1.342134e-07, 1.342134e-07, 
    1.342133e-07, 1.342133e-07, 1.342135e-07, 1.342134e-07, 1.342137e-07, 
    1.342136e-07, 1.342137e-07, 1.342138e-07, 1.342134e-07, 1.342136e-07, 
    1.342133e-07, 1.342134e-07, 1.342131e-07, 1.342132e-07, 1.342129e-07, 
    1.342128e-07, 1.342127e-07, 1.342125e-07, 1.342137e-07, 1.342137e-07, 
    1.342137e-07, 1.342136e-07, 1.342135e-07, 1.342134e-07, 1.342134e-07, 
    1.342133e-07, 1.342133e-07, 1.342132e-07, 1.342133e-07, 1.342132e-07, 
    1.342136e-07, 1.342134e-07, 1.342138e-07, 1.342137e-07, 1.342136e-07, 
    1.342136e-07, 1.342135e-07, 1.342134e-07, 1.342133e-07, 1.342133e-07, 
    1.342128e-07, 1.342131e-07, 1.342124e-07, 1.342126e-07, 1.342138e-07, 
    1.342137e-07, 1.342135e-07, 1.342136e-07, 1.342134e-07, 1.342133e-07, 
    1.342132e-07, 1.342132e-07, 1.342132e-07, 1.342131e-07, 1.342132e-07, 
    1.342131e-07, 1.342134e-07, 1.342133e-07, 1.342135e-07, 1.342135e-07, 
    1.342135e-07, 1.342135e-07, 1.342134e-07, 1.342133e-07, 1.342133e-07, 
    1.342133e-07, 1.342132e-07, 1.342134e-07, 1.342128e-07, 1.342131e-07, 
    1.342136e-07, 1.342136e-07, 1.342135e-07, 1.342136e-07, 1.342133e-07, 
    1.342134e-07, 1.342131e-07, 1.342132e-07, 1.342131e-07, 1.342131e-07, 
    1.342132e-07, 1.342132e-07, 1.342133e-07, 1.342134e-07, 1.342135e-07, 
    1.342136e-07, 1.342136e-07, 1.342135e-07, 1.342133e-07, 1.342132e-07, 
    1.342132e-07, 1.342131e-07, 1.342134e-07, 1.342133e-07, 1.342133e-07, 
    1.342132e-07, 1.342134e-07, 1.342132e-07, 1.342135e-07, 1.342135e-07, 
    1.342134e-07, 1.342133e-07, 1.342132e-07, 1.342132e-07, 1.342132e-07, 
    1.342133e-07, 1.342133e-07, 1.342134e-07, 1.342134e-07, 1.342135e-07, 
    1.342135e-07, 1.342135e-07, 1.342134e-07, 1.342133e-07, 1.342132e-07, 
    1.342131e-07, 1.34213e-07, 1.342129e-07, 1.34213e-07, 1.342128e-07, 
    1.34213e-07, 1.342127e-07, 1.342132e-07, 1.34213e-07, 1.342134e-07, 
    1.342134e-07, 1.342133e-07, 1.342131e-07, 1.342132e-07, 1.342131e-07, 
    1.342133e-07, 1.342135e-07, 1.342135e-07, 1.342136e-07, 1.342135e-07, 
    1.342135e-07, 1.342134e-07, 1.342135e-07, 1.342133e-07, 1.342134e-07, 
    1.342132e-07, 1.342131e-07, 1.342128e-07, 1.342127e-07, 1.342125e-07, 
    1.342125e-07, 1.342124e-07, 1.342124e-07 ;

 LITR3N_TNDNCY_VERT_TRANS =
  1.715634e-26, -3.798904e-26, 1.225453e-26, -5.882173e-26, 8.700715e-26, 
    5.269447e-26, 7.352717e-27, -1.372507e-25, -1.225453e-26, -3.063632e-26, 
    -1.02938e-25, 4.779266e-26, -5.269447e-26, -4.779266e-26, -6.004719e-26, 
    3.553813e-26, -2.941087e-26, -3.186177e-26, 1.249962e-25, -4.166539e-26, 
    1.960724e-26, -1.556325e-25, -2.941087e-26, 1.397016e-25, 3.308722e-26, 
    2.941087e-26, -3.676358e-26, -1.041635e-25, 1.225453e-27, -7.965443e-26, 
    3.676358e-26, 4.41163e-26, -7.720352e-26, 1.274471e-25, 5.024356e-26, 
    -1.347998e-26, 5.882173e-26, -4.289085e-26, -8.333079e-26, -6.862535e-26, 
    3.553813e-26, 2.08327e-26, -2.450905e-26, -4.901811e-26, -6.617445e-26, 
    -3.063632e-26, 8.82326e-26, 7.720352e-26, 7.842898e-26, -4.534175e-26, 
    2.941087e-26, -1.838179e-26, -1.004871e-25, 1.838179e-26, -1.102908e-26, 
    -1.225453e-26, 5.146902e-26, -3.431268e-26, 4.901811e-26, -9.803622e-27, 
    4.779266e-26, 3.308722e-26, -4.779266e-26, -4.043994e-26, 3.063632e-26, 
    -4.289085e-26, -1.102908e-26, -6.004719e-26, 2.941087e-26, -2.205815e-26, 
    -4.41163e-26, -8.087988e-26, 5.882173e-26, 1.715634e-26, 4.289085e-26, 
    1.838179e-26, -7.652491e-42, 1.715634e-26, -1.593089e-26, -1.225453e-27, 
    4.534175e-26, -6.127264e-27, -6.127264e-27, -1.593089e-26, 1.311234e-25, 
    1.225453e-27, 1.838179e-26, -1.960724e-26, 6.372354e-26, -2.695996e-26, 
    -3.676358e-26, 1.593089e-26, -3.921449e-26, -2.818541e-26, -6.4949e-26, 
    5.269447e-26, 2.32836e-26, 6.127264e-26, 5.269447e-26, -6.617445e-26, 
    -5.269447e-26, 4.901811e-27, 9.803622e-27, -3.431268e-26, 6.127264e-26, 
    -3.676358e-27, -4.289085e-26, -1.053889e-25, -7.107626e-26, 4.779266e-26, 
    -1.470543e-26, 5.637083e-26, -2.941087e-26, 3.676358e-27, -6.4949e-26, 
    -4.289085e-26, -1.127417e-25, 9.926167e-26, 1.151926e-25, -1.347998e-26, 
    -4.289085e-26, -6.862535e-26, -4.534175e-26, 4.043994e-26, 6.617445e-26, 
    1.139671e-25, -4.901811e-26, -8.578169e-26, -2.818541e-26, 3.676358e-27, 
    1.960724e-26, -4.901811e-27, 2.941087e-26, -5.637083e-26, -3.063632e-26, 
    -6.617445e-26, -7.352717e-26, -2.695996e-26, 2.450905e-26, -3.921449e-26, 
    1.470543e-26, 1.213198e-25, 6.127264e-27, 5.514538e-26, -3.063632e-26, 
    7.842898e-26, 5.146902e-26, 3.798904e-26, 2.205815e-26, 8.578169e-27, 
    6.98508e-26, -2.818541e-26, 5.269447e-26, 5.269447e-26, 6.372354e-26, 
    -7.597807e-26, -8.945805e-26, -4.65672e-26, 1.838179e-26, 6.004719e-26, 
    1.838179e-26, 9.068351e-26, 6.73999e-26, -5.882173e-26, 1.470543e-26, 
    -7.352717e-27, 3.676358e-27, -6.249809e-26, 7.230172e-26, -7.352717e-27, 
    8.578169e-27, 2.32836e-26, -4.65672e-26, -6.127264e-26, 3.676358e-27, 
    1.102908e-26, 8.333079e-26, 2.573451e-26, 3.308722e-26, 2.573451e-26, 
    -1.115162e-25, 5.146902e-26, -3.431268e-26, -9.190896e-26, -1.102908e-26, 
    -1.593089e-26, 2.32836e-26, 9.926167e-26, -1.078398e-25, -1.347998e-26, 
    7.230172e-26, -2.08327e-26, 2.32836e-26, 6.617445e-26, -5.759628e-26, 
    -2.941087e-26, 1.225453e-27, 9.803622e-26, 1.347998e-26, 2.450905e-26, 
    -6.372354e-26, -8.210533e-26, 4.289085e-26, 1.776906e-25, -1.102908e-26, 
    4.901811e-26, -1.593089e-26, 4.166539e-26, 7.107626e-26, 2.450906e-27, 
    2.450905e-26, -5.024356e-26, -2.695996e-26, 1.225453e-26, -1.16418e-25, 
    -6.004719e-26, 4.289085e-26, 2.08327e-26, 2.941087e-26, -5.391992e-26, 
    -5.637083e-26, -6.617445e-26, 3.308722e-26, -8.333079e-26, -3.921449e-26, 
    -6.862535e-26, 7.352717e-27, 9.803622e-27, -6.127264e-26, -5.882173e-26, 
    -5.146902e-26, -5.024356e-26, 1.347998e-26, -9.803622e-26, -5.024356e-26, 
    8.578169e-27, 4.901811e-26, -8.210533e-26, -1.102908e-26, -5.146902e-26, 
    0, 7.475262e-26, 3.186177e-26, -7.230172e-26, 1.740143e-25, 4.901811e-26, 
    -2.009742e-25, -2.450905e-26, -2.573451e-26, -6.127264e-27, 
    -8.455624e-26, 2.08327e-26, 8.578169e-27, -7.107626e-26, 7.352717e-27, 
    -6.73999e-26, 4.41163e-26, -1.838179e-26, 5.514538e-26, 5.146902e-26, 
    4.779266e-26, -5.146902e-26, 3.826946e-42, -1.470543e-25, 7.352717e-27, 
    1.004871e-25, 2.205815e-26, -4.41163e-26, 1.43378e-25, -5.882173e-26, 
    9.803622e-27, -1.078398e-25, -1.43378e-25, 1.519561e-25, -8.578169e-27, 
    -4.901811e-27, 9.681077e-26, -4.534175e-26, -8.210533e-26, 2.941087e-26, 
    2.941087e-26, -1.470543e-25, -1.470543e-26, 5.514538e-26, 3.676358e-27, 
    -5.269447e-26, 4.779266e-26, -3.921449e-26, 9.558531e-26, 2.08327e-26, 
    -1.139671e-25, -5.391992e-26, -3.553813e-26, 1.666616e-25, 1.225453e-27, 
    2.695996e-26, 3.431268e-26, -4.166539e-26, -9.068351e-26, -2.450905e-26, 
    -1.960724e-26, 1.347998e-26, 3.431268e-26, 1.960724e-26, -1.151926e-25, 
    -3.308722e-26, 6.127264e-26, 8.578169e-27, -1.102908e-26, -1.29898e-25, 
    -2.941087e-26, -9.068351e-26, -4.166539e-26, 8.578169e-27, -1.421525e-25, 
    -8.210533e-26, -5.759628e-26, 4.166539e-26, -4.779266e-26, -4.166539e-26, 
    -1.102908e-26, -2.695996e-26, -7.842898e-26, 8.210533e-26, 1.225453e-27, 
    4.41163e-26, 3.921449e-26, -4.41163e-26, 4.534175e-26, -1.115162e-25, 
    2.450906e-27, -1.347998e-25, -9.435986e-26, 1.151926e-25, 5.146902e-26, 
    4.901811e-26, -4.41163e-26, 2.695996e-26,
  1.338134e-32, 1.338132e-32, 1.338133e-32, 1.338131e-32, 1.338132e-32, 
    1.338131e-32, 1.338134e-32, 1.338132e-32, 1.338133e-32, 1.338134e-32, 
    1.338129e-32, 1.338131e-32, 1.338127e-32, 1.338129e-32, 1.338125e-32, 
    1.338127e-32, 1.338125e-32, 1.338125e-32, 1.338124e-32, 1.338124e-32, 
    1.338122e-32, 1.338123e-32, 1.338121e-32, 1.338123e-32, 1.338122e-32, 
    1.338124e-32, 1.338131e-32, 1.33813e-32, 1.338131e-32, 1.338131e-32, 
    1.338131e-32, 1.338132e-32, 1.338133e-32, 1.338134e-32, 1.338134e-32, 
    1.338133e-32, 1.338131e-32, 1.338131e-32, 1.33813e-32, 1.33813e-32, 
    1.338128e-32, 1.338129e-32, 1.338126e-32, 1.338127e-32, 1.338124e-32, 
    1.338125e-32, 1.338124e-32, 1.338124e-32, 1.338124e-32, 1.338125e-32, 
    1.338125e-32, 1.338125e-32, 1.338129e-32, 1.338128e-32, 1.338131e-32, 
    1.338132e-32, 1.338133e-32, 1.338134e-32, 1.338134e-32, 1.338134e-32, 
    1.338133e-32, 1.338132e-32, 1.338131e-32, 1.33813e-32, 1.33813e-32, 
    1.338128e-32, 1.338128e-32, 1.338126e-32, 1.338126e-32, 1.338125e-32, 
    1.338125e-32, 1.338124e-32, 1.338124e-32, 1.338124e-32, 1.338125e-32, 
    1.338124e-32, 1.338126e-32, 1.338126e-32, 1.33813e-32, 1.338131e-32, 
    1.338132e-32, 1.338133e-32, 1.338134e-32, 1.338133e-32, 1.338133e-32, 
    1.338133e-32, 1.338132e-32, 1.338132e-32, 1.33813e-32, 1.338131e-32, 
    1.338127e-32, 1.338129e-32, 1.338125e-32, 1.338126e-32, 1.338125e-32, 
    1.338125e-32, 1.338124e-32, 1.338125e-32, 1.338123e-32, 1.338123e-32, 
    1.338123e-32, 1.338122e-32, 1.338125e-32, 1.338124e-32, 1.338132e-32, 
    1.338132e-32, 1.338132e-32, 1.338133e-32, 1.338133e-32, 1.338134e-32, 
    1.338133e-32, 1.338133e-32, 1.338132e-32, 1.338131e-32, 1.338131e-32, 
    1.33813e-32, 1.338129e-32, 1.338127e-32, 1.338126e-32, 1.338125e-32, 
    1.338125e-32, 1.338125e-32, 1.338125e-32, 1.338126e-32, 1.338123e-32, 
    1.338125e-32, 1.338123e-32, 1.338123e-32, 1.338124e-32, 1.338123e-32, 
    1.338132e-32, 1.338132e-32, 1.338133e-32, 1.338133e-32, 1.338134e-32, 
    1.338133e-32, 1.338133e-32, 1.338131e-32, 1.338131e-32, 1.33813e-32, 
    1.33813e-32, 1.338129e-32, 1.338127e-32, 1.338126e-32, 1.338125e-32, 
    1.338125e-32, 1.338125e-32, 1.338125e-32, 1.338125e-32, 1.338124e-32, 
    1.338124e-32, 1.338125e-32, 1.338123e-32, 1.338123e-32, 1.338123e-32, 
    1.338123e-32, 1.338132e-32, 1.338132e-32, 1.338132e-32, 1.338132e-32, 
    1.338132e-32, 1.33813e-32, 1.33813e-32, 1.338128e-32, 1.338129e-32, 
    1.338128e-32, 1.338129e-32, 1.338129e-32, 1.338128e-32, 1.338129e-32, 
    1.338126e-32, 1.338128e-32, 1.338125e-32, 1.338126e-32, 1.338124e-32, 
    1.338125e-32, 1.338124e-32, 1.338124e-32, 1.338123e-32, 1.338122e-32, 
    1.338122e-32, 1.338121e-32, 1.338131e-32, 1.338131e-32, 1.338131e-32, 
    1.33813e-32, 1.33813e-32, 1.338129e-32, 1.338127e-32, 1.338128e-32, 
    1.338126e-32, 1.338126e-32, 1.338128e-32, 1.338127e-32, 1.33813e-32, 
    1.33813e-32, 1.33813e-32, 1.338131e-32, 1.338127e-32, 1.338129e-32, 
    1.338126e-32, 1.338127e-32, 1.338124e-32, 1.338125e-32, 1.338122e-32, 
    1.338121e-32, 1.33812e-32, 1.338119e-32, 1.33813e-32, 1.338131e-32, 
    1.33813e-32, 1.338129e-32, 1.338128e-32, 1.338127e-32, 1.338127e-32, 
    1.338126e-32, 1.338126e-32, 1.338125e-32, 1.338126e-32, 1.338125e-32, 
    1.338129e-32, 1.338127e-32, 1.338131e-32, 1.33813e-32, 1.338129e-32, 
    1.338129e-32, 1.338128e-32, 1.338127e-32, 1.338126e-32, 1.338126e-32, 
    1.338121e-32, 1.338124e-32, 1.338118e-32, 1.338119e-32, 1.338131e-32, 
    1.33813e-32, 1.338128e-32, 1.338129e-32, 1.338127e-32, 1.338126e-32, 
    1.338125e-32, 1.338125e-32, 1.338125e-32, 1.338124e-32, 1.338125e-32, 
    1.338124e-32, 1.338127e-32, 1.338126e-32, 1.338129e-32, 1.338128e-32, 
    1.338128e-32, 1.338129e-32, 1.338127e-32, 1.338126e-32, 1.338126e-32, 
    1.338126e-32, 1.338125e-32, 1.338127e-32, 1.338121e-32, 1.338125e-32, 
    1.33813e-32, 1.338129e-32, 1.338128e-32, 1.338129e-32, 1.338126e-32, 
    1.338127e-32, 1.338124e-32, 1.338125e-32, 1.338124e-32, 1.338125e-32, 
    1.338125e-32, 1.338125e-32, 1.338126e-32, 1.338127e-32, 1.338128e-32, 
    1.338129e-32, 1.338129e-32, 1.338128e-32, 1.338126e-32, 1.338125e-32, 
    1.338125e-32, 1.338124e-32, 1.338127e-32, 1.338126e-32, 1.338126e-32, 
    1.338125e-32, 1.338128e-32, 1.338125e-32, 1.338128e-32, 1.338128e-32, 
    1.338127e-32, 1.338126e-32, 1.338125e-32, 1.338125e-32, 1.338125e-32, 
    1.338126e-32, 1.338126e-32, 1.338127e-32, 1.338127e-32, 1.338128e-32, 
    1.338128e-32, 1.338128e-32, 1.338128e-32, 1.338126e-32, 1.338125e-32, 
    1.338124e-32, 1.338123e-32, 1.338122e-32, 1.338123e-32, 1.338121e-32, 
    1.338123e-32, 1.33812e-32, 1.338125e-32, 1.338123e-32, 1.338127e-32, 
    1.338127e-32, 1.338126e-32, 1.338124e-32, 1.338125e-32, 1.338124e-32, 
    1.338126e-32, 1.338128e-32, 1.338128e-32, 1.338129e-32, 1.338128e-32, 
    1.338128e-32, 1.338128e-32, 1.338128e-32, 1.338126e-32, 1.338127e-32, 
    1.338125e-32, 1.338124e-32, 1.338121e-32, 1.33812e-32, 1.338118e-32, 
    1.338118e-32, 1.338118e-32, 1.338117e-32,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3N_TO_SOIL2N =
  1.643693e-15, 1.6482e-15, 1.647324e-15, 1.650956e-15, 1.648943e-15, 
    1.65132e-15, 1.644608e-15, 1.648378e-15, 1.645972e-15, 1.6441e-15, 
    1.657997e-15, 1.651119e-15, 1.665139e-15, 1.660758e-15, 1.671759e-15, 
    1.664457e-15, 1.673231e-15, 1.67155e-15, 1.67661e-15, 1.675161e-15, 
    1.681625e-15, 1.677279e-15, 1.684974e-15, 1.680588e-15, 1.681274e-15, 
    1.677135e-15, 1.652505e-15, 1.65714e-15, 1.65223e-15, 1.652891e-15, 
    1.652595e-15, 1.648984e-15, 1.647162e-15, 1.64335e-15, 1.644042e-15, 
    1.646843e-15, 1.653189e-15, 1.651036e-15, 1.656462e-15, 1.65634e-15, 
    1.662374e-15, 1.659654e-15, 1.669787e-15, 1.666909e-15, 1.675222e-15, 
    1.673132e-15, 1.675123e-15, 1.67452e-15, 1.675131e-15, 1.672066e-15, 
    1.67338e-15, 1.670682e-15, 1.660163e-15, 1.663256e-15, 1.654025e-15, 
    1.648465e-15, 1.644773e-15, 1.642151e-15, 1.642521e-15, 1.643228e-15, 
    1.646859e-15, 1.650272e-15, 1.652872e-15, 1.65461e-15, 1.656322e-15, 
    1.661497e-15, 1.664238e-15, 1.670368e-15, 1.669263e-15, 1.671135e-15, 
    1.672924e-15, 1.675925e-15, 1.675432e-15, 1.676753e-15, 1.671087e-15, 
    1.674853e-15, 1.668634e-15, 1.670335e-15, 1.656782e-15, 1.651617e-15, 
    1.649416e-15, 1.647492e-15, 1.642806e-15, 1.646043e-15, 1.644767e-15, 
    1.647803e-15, 1.64973e-15, 1.648777e-15, 1.654658e-15, 1.652372e-15, 
    1.664401e-15, 1.659223e-15, 1.672716e-15, 1.66949e-15, 1.673489e-15, 
    1.671449e-15, 1.674943e-15, 1.671799e-15, 1.677245e-15, 1.67843e-15, 
    1.67762e-15, 1.680731e-15, 1.671624e-15, 1.675123e-15, 1.64875e-15, 
    1.648905e-15, 1.64963e-15, 1.646444e-15, 1.64625e-15, 1.64333e-15, 
    1.645928e-15, 1.647034e-15, 1.649842e-15, 1.651501e-15, 1.653078e-15, 
    1.656545e-15, 1.660412e-15, 1.665818e-15, 1.669699e-15, 1.672299e-15, 
    1.670705e-15, 1.672112e-15, 1.670539e-15, 1.669802e-15, 1.677986e-15, 
    1.673392e-15, 1.680284e-15, 1.679903e-15, 1.676784e-15, 1.679946e-15, 
    1.649015e-15, 1.64812e-15, 1.645012e-15, 1.647444e-15, 1.643013e-15, 
    1.645493e-15, 1.646918e-15, 1.652418e-15, 1.653627e-15, 1.654747e-15, 
    1.656958e-15, 1.659793e-15, 1.664764e-15, 1.669086e-15, 1.673029e-15, 
    1.67274e-15, 1.672842e-15, 1.673722e-15, 1.671541e-15, 1.67408e-15, 
    1.674505e-15, 1.673392e-15, 1.679852e-15, 1.678007e-15, 1.679895e-15, 
    1.678694e-15, 1.648411e-15, 1.649916e-15, 1.649103e-15, 1.650632e-15, 
    1.649554e-15, 1.654343e-15, 1.655778e-15, 1.662489e-15, 1.659737e-15, 
    1.664118e-15, 1.660183e-15, 1.66088e-15, 1.664258e-15, 1.660396e-15, 
    1.668846e-15, 1.663116e-15, 1.673756e-15, 1.668037e-15, 1.674114e-15, 
    1.673012e-15, 1.674837e-15, 1.67647e-15, 1.678526e-15, 1.682314e-15, 
    1.681438e-15, 1.684605e-15, 1.65216e-15, 1.65411e-15, 1.653939e-15, 
    1.655981e-15, 1.657489e-15, 1.66076e-15, 1.666e-15, 1.66403e-15, 
    1.667647e-15, 1.668372e-15, 1.662878e-15, 1.666251e-15, 1.655416e-15, 
    1.657167e-15, 1.656125e-15, 1.652313e-15, 1.664483e-15, 1.65824e-15, 
    1.669763e-15, 1.666386e-15, 1.676237e-15, 1.671339e-15, 1.680955e-15, 
    1.685057e-15, 1.68892e-15, 1.693424e-15, 1.655175e-15, 1.65385e-15, 
    1.656224e-15, 1.659504e-15, 1.662548e-15, 1.666591e-15, 1.667006e-15, 
    1.667762e-15, 1.669723e-15, 1.671371e-15, 1.668001e-15, 1.671784e-15, 
    1.657571e-15, 1.665025e-15, 1.653348e-15, 1.656865e-15, 1.659311e-15, 
    1.658239e-15, 1.663805e-15, 1.665116e-15, 1.670439e-15, 1.667688e-15, 
    1.684044e-15, 1.676814e-15, 1.696854e-15, 1.691261e-15, 1.653387e-15, 
    1.655171e-15, 1.661375e-15, 1.658424e-15, 1.666862e-15, 1.668936e-15, 
    1.670623e-15, 1.672776e-15, 1.67301e-15, 1.674285e-15, 1.672195e-15, 
    1.674203e-15, 1.6666e-15, 1.669999e-15, 1.660668e-15, 1.66294e-15, 
    1.661895e-15, 1.660748e-15, 1.664287e-15, 1.668053e-15, 1.668136e-15, 
    1.669342e-15, 1.672739e-15, 1.666896e-15, 1.684973e-15, 1.673814e-15, 
    1.657116e-15, 1.660548e-15, 1.66104e-15, 1.659711e-15, 1.668728e-15, 
    1.665462e-15, 1.674255e-15, 1.67188e-15, 1.67577e-15, 1.673837e-15, 
    1.673553e-15, 1.671069e-15, 1.669522e-15, 1.665612e-15, 1.662428e-15, 
    1.659904e-15, 1.660491e-15, 1.663264e-15, 1.668284e-15, 1.67303e-15, 
    1.671991e-15, 1.675475e-15, 1.66625e-15, 1.67012e-15, 1.668624e-15, 
    1.672523e-15, 1.663977e-15, 1.67125e-15, 1.662116e-15, 1.662918e-15, 
    1.665397e-15, 1.670381e-15, 1.671485e-15, 1.672661e-15, 1.671936e-15, 
    1.668412e-15, 1.667835e-15, 1.665338e-15, 1.664647e-15, 1.662744e-15, 
    1.661167e-15, 1.662607e-15, 1.664119e-15, 1.668414e-15, 1.672281e-15, 
    1.676493e-15, 1.677525e-15, 1.682437e-15, 1.678436e-15, 1.685035e-15, 
    1.679422e-15, 1.689136e-15, 1.671674e-15, 1.67926e-15, 1.665511e-15, 
    1.666994e-15, 1.669674e-15, 1.67582e-15, 1.672505e-15, 1.676382e-15, 
    1.667813e-15, 1.663359e-15, 1.662208e-15, 1.660057e-15, 1.662257e-15, 
    1.662078e-15, 1.664183e-15, 1.663507e-15, 1.668557e-15, 1.665845e-15, 
    1.673545e-15, 1.676352e-15, 1.684273e-15, 1.689121e-15, 1.694054e-15, 
    1.696229e-15, 1.696891e-15, 1.697168e-15 ;

 LITR3N_vr =
  7.663762e-06, 7.663753e-06, 7.663755e-06, 7.663749e-06, 7.663753e-06, 
    7.663748e-06, 7.66376e-06, 7.663753e-06, 7.663758e-06, 7.663761e-06, 
    7.663737e-06, 7.663749e-06, 7.663724e-06, 7.663732e-06, 7.663712e-06, 
    7.663725e-06, 7.66371e-06, 7.663713e-06, 7.663704e-06, 7.663707e-06, 
    7.663695e-06, 7.663703e-06, 7.66369e-06, 7.663697e-06, 7.663696e-06, 
    7.663703e-06, 7.663746e-06, 7.663738e-06, 7.663747e-06, 7.663745e-06, 
    7.663746e-06, 7.663753e-06, 7.663755e-06, 7.663763e-06, 7.663761e-06, 
    7.663756e-06, 7.663745e-06, 7.663749e-06, 7.663739e-06, 7.66374e-06, 
    7.663729e-06, 7.663733e-06, 7.663716e-06, 7.663722e-06, 7.663707e-06, 
    7.663711e-06, 7.663707e-06, 7.663708e-06, 7.663707e-06, 7.663712e-06, 
    7.66371e-06, 7.663714e-06, 7.663733e-06, 7.663727e-06, 7.663743e-06, 
    7.663753e-06, 7.66376e-06, 7.663764e-06, 7.663763e-06, 7.663763e-06, 
    7.663756e-06, 7.66375e-06, 7.663745e-06, 7.663743e-06, 7.66374e-06, 
    7.663731e-06, 7.663726e-06, 7.663715e-06, 7.663717e-06, 7.663713e-06, 
    7.663711e-06, 7.663705e-06, 7.663706e-06, 7.663704e-06, 7.663714e-06, 
    7.663707e-06, 7.663718e-06, 7.663715e-06, 7.663739e-06, 7.663748e-06, 
    7.663752e-06, 7.663755e-06, 7.663763e-06, 7.663757e-06, 7.66376e-06, 
    7.663754e-06, 7.663751e-06, 7.663753e-06, 7.663743e-06, 7.663746e-06, 
    7.663725e-06, 7.663734e-06, 7.663711e-06, 7.663717e-06, 7.66371e-06, 
    7.663713e-06, 7.663707e-06, 7.663712e-06, 7.663703e-06, 7.663701e-06, 
    7.663702e-06, 7.663697e-06, 7.663712e-06, 7.663707e-06, 7.663753e-06, 
    7.663753e-06, 7.663752e-06, 7.663757e-06, 7.663757e-06, 7.663763e-06, 
    7.663758e-06, 7.663756e-06, 7.663751e-06, 7.663748e-06, 7.663745e-06, 
    7.663739e-06, 7.663733e-06, 7.663723e-06, 7.663716e-06, 7.663712e-06, 
    7.663714e-06, 7.663712e-06, 7.663715e-06, 7.663716e-06, 7.663702e-06, 
    7.66371e-06, 7.663698e-06, 7.663699e-06, 7.663704e-06, 7.663699e-06, 
    7.663753e-06, 7.663753e-06, 7.663759e-06, 7.663755e-06, 7.663763e-06, 
    7.663758e-06, 7.663756e-06, 7.663746e-06, 7.663744e-06, 7.663743e-06, 
    7.663739e-06, 7.663733e-06, 7.663725e-06, 7.663717e-06, 7.663711e-06, 
    7.663711e-06, 7.663711e-06, 7.663709e-06, 7.663713e-06, 7.663709e-06, 
    7.663708e-06, 7.66371e-06, 7.663699e-06, 7.663702e-06, 7.663699e-06, 
    7.663701e-06, 7.663753e-06, 7.663751e-06, 7.663753e-06, 7.66375e-06, 
    7.663752e-06, 7.663743e-06, 7.663741e-06, 7.663729e-06, 7.663733e-06, 
    7.663726e-06, 7.663733e-06, 7.663732e-06, 7.663726e-06, 7.663733e-06, 
    7.663718e-06, 7.663728e-06, 7.663709e-06, 7.663719e-06, 7.663709e-06, 
    7.663711e-06, 7.663707e-06, 7.663704e-06, 7.663701e-06, 7.663694e-06, 
    7.663696e-06, 7.663691e-06, 7.663747e-06, 7.663743e-06, 7.663743e-06, 
    7.66374e-06, 7.663738e-06, 7.663732e-06, 7.663722e-06, 7.663726e-06, 
    7.66372e-06, 7.663719e-06, 7.663728e-06, 7.663722e-06, 7.663742e-06, 
    7.663738e-06, 7.66374e-06, 7.663746e-06, 7.663725e-06, 7.663736e-06, 
    7.663716e-06, 7.663722e-06, 7.663705e-06, 7.663713e-06, 7.663697e-06, 
    7.66369e-06, 7.663682e-06, 7.663675e-06, 7.663742e-06, 7.663743e-06, 
    7.66374e-06, 7.663734e-06, 7.663729e-06, 7.663722e-06, 7.663721e-06, 
    7.66372e-06, 7.663716e-06, 7.663713e-06, 7.663719e-06, 7.663712e-06, 
    7.663737e-06, 7.663724e-06, 7.663744e-06, 7.663739e-06, 7.663734e-06, 
    7.663736e-06, 7.663726e-06, 7.663724e-06, 7.663715e-06, 7.66372e-06, 
    7.663692e-06, 7.663704e-06, 7.663669e-06, 7.663679e-06, 7.663744e-06, 
    7.663742e-06, 7.663731e-06, 7.663736e-06, 7.663722e-06, 7.663718e-06, 
    7.663714e-06, 7.663711e-06, 7.663711e-06, 7.663708e-06, 7.663712e-06, 
    7.663709e-06, 7.663722e-06, 7.663716e-06, 7.663732e-06, 7.663728e-06, 
    7.66373e-06, 7.663732e-06, 7.663726e-06, 7.663719e-06, 7.663719e-06, 
    7.663717e-06, 7.663711e-06, 7.663722e-06, 7.66369e-06, 7.663709e-06, 
    7.663738e-06, 7.663733e-06, 7.663732e-06, 7.663733e-06, 7.663718e-06, 
    7.663723e-06, 7.663708e-06, 7.663712e-06, 7.663706e-06, 7.663709e-06, 
    7.66371e-06, 7.663714e-06, 7.663716e-06, 7.663723e-06, 7.663729e-06, 
    7.663733e-06, 7.663733e-06, 7.663727e-06, 7.663719e-06, 7.663711e-06, 
    7.663712e-06, 7.663706e-06, 7.663722e-06, 7.663715e-06, 7.663718e-06, 
    7.663712e-06, 7.663726e-06, 7.663713e-06, 7.66373e-06, 7.663728e-06, 
    7.663723e-06, 7.663715e-06, 7.663713e-06, 7.663711e-06, 7.663712e-06, 
    7.663719e-06, 7.66372e-06, 7.663724e-06, 7.663725e-06, 7.663728e-06, 
    7.663731e-06, 7.663729e-06, 7.663726e-06, 7.663719e-06, 7.663712e-06, 
    7.663704e-06, 7.663702e-06, 7.663694e-06, 7.663701e-06, 7.66369e-06, 
    7.6637e-06, 7.663682e-06, 7.663712e-06, 7.6637e-06, 7.663723e-06, 
    7.663721e-06, 7.663716e-06, 7.663705e-06, 7.663712e-06, 7.663704e-06, 
    7.66372e-06, 7.663727e-06, 7.66373e-06, 7.663733e-06, 7.663729e-06, 
    7.66373e-06, 7.663726e-06, 7.663727e-06, 7.663718e-06, 7.663723e-06, 
    7.66371e-06, 7.663704e-06, 7.663691e-06, 7.663682e-06, 7.663674e-06, 
    7.66367e-06, 7.663669e-06, 7.663669e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LITR3_HR =
  5.938512e-14, 5.954794e-14, 5.951631e-14, 5.964753e-14, 5.957477e-14, 
    5.966066e-14, 5.941816e-14, 5.955438e-14, 5.946745e-14, 5.939982e-14, 
    5.990189e-14, 5.965339e-14, 6.015994e-14, 6.000165e-14, 6.039911e-14, 
    6.013528e-14, 6.045228e-14, 6.039157e-14, 6.057439e-14, 6.052204e-14, 
    6.075555e-14, 6.059855e-14, 6.087658e-14, 6.07181e-14, 6.074287e-14, 
    6.059336e-14, 5.970348e-14, 5.987095e-14, 5.969354e-14, 5.971744e-14, 
    5.970673e-14, 5.957625e-14, 5.951043e-14, 5.937271e-14, 5.939773e-14, 
    5.949891e-14, 5.972818e-14, 5.965042e-14, 5.984646e-14, 5.984203e-14, 
    6.006002e-14, 5.996177e-14, 6.032785e-14, 6.022389e-14, 6.052422e-14, 
    6.044872e-14, 6.052067e-14, 6.049886e-14, 6.052095e-14, 6.041022e-14, 
    6.045767e-14, 6.036022e-14, 5.998016e-14, 6.009191e-14, 5.97584e-14, 
    5.955752e-14, 5.942413e-14, 5.932939e-14, 5.934278e-14, 5.936831e-14, 
    5.94995e-14, 5.962283e-14, 5.971674e-14, 5.977953e-14, 5.984139e-14, 
    6.002837e-14, 6.012739e-14, 6.034884e-14, 6.030895e-14, 6.037657e-14, 
    6.044122e-14, 6.054964e-14, 6.053181e-14, 6.057955e-14, 6.037482e-14, 
    6.051089e-14, 6.028621e-14, 6.034768e-14, 5.985801e-14, 5.967141e-14, 
    5.959187e-14, 5.952238e-14, 5.935308e-14, 5.947e-14, 5.942391e-14, 
    5.953358e-14, 5.960321e-14, 5.956879e-14, 5.978125e-14, 5.969867e-14, 
    6.013326e-14, 5.994618e-14, 6.043368e-14, 6.031714e-14, 6.04616e-14, 
    6.038791e-14, 6.051415e-14, 6.040054e-14, 6.059733e-14, 6.064013e-14, 
    6.061087e-14, 6.072328e-14, 6.039424e-14, 6.052065e-14, 5.956782e-14, 
    5.957343e-14, 5.95996e-14, 5.948452e-14, 5.947748e-14, 5.937202e-14, 
    5.946588e-14, 5.950582e-14, 5.960727e-14, 5.966721e-14, 5.972419e-14, 
    5.984943e-14, 5.998917e-14, 6.018447e-14, 6.03247e-14, 6.041862e-14, 
    6.036105e-14, 6.041188e-14, 6.035505e-14, 6.032841e-14, 6.062408e-14, 
    6.045809e-14, 6.070712e-14, 6.069335e-14, 6.058067e-14, 6.06949e-14, 
    5.957737e-14, 5.954506e-14, 5.943276e-14, 5.952065e-14, 5.936053e-14, 
    5.945015e-14, 5.950165e-14, 5.970035e-14, 5.974403e-14, 5.978447e-14, 
    5.986434e-14, 5.99668e-14, 6.014637e-14, 6.030252e-14, 6.044498e-14, 
    6.043455e-14, 6.043823e-14, 6.047001e-14, 6.039123e-14, 6.048295e-14, 
    6.049832e-14, 6.04581e-14, 6.069151e-14, 6.062486e-14, 6.069306e-14, 
    6.064967e-14, 5.955557e-14, 5.960994e-14, 5.958056e-14, 5.96358e-14, 
    5.959687e-14, 5.976988e-14, 5.982172e-14, 6.006419e-14, 5.996477e-14, 
    6.012304e-14, 5.998086e-14, 6.000605e-14, 6.012811e-14, 5.998856e-14, 
    6.029387e-14, 6.008686e-14, 6.047125e-14, 6.026463e-14, 6.048419e-14, 
    6.044437e-14, 6.051031e-14, 6.056933e-14, 6.064359e-14, 6.078047e-14, 
    6.074879e-14, 6.086323e-14, 5.969101e-14, 5.976147e-14, 5.97553e-14, 
    5.982905e-14, 5.988356e-14, 6.000172e-14, 6.019104e-14, 6.011988e-14, 
    6.025053e-14, 6.027673e-14, 6.007825e-14, 6.020011e-14, 5.980864e-14, 
    5.98719e-14, 5.983427e-14, 5.969654e-14, 6.013622e-14, 5.991067e-14, 
    6.0327e-14, 6.020497e-14, 6.056091e-14, 6.038394e-14, 6.073134e-14, 
    6.087955e-14, 6.101911e-14, 6.118185e-14, 5.979996e-14, 5.975209e-14, 
    5.983783e-14, 5.995633e-14, 6.006633e-14, 6.021241e-14, 6.022737e-14, 
    6.025471e-14, 6.032556e-14, 6.03851e-14, 6.026332e-14, 6.040002e-14, 
    5.98865e-14, 6.015581e-14, 5.973395e-14, 5.986102e-14, 5.994937e-14, 
    5.991065e-14, 6.011175e-14, 6.015911e-14, 6.03514e-14, 6.025204e-14, 
    6.084295e-14, 6.058174e-14, 6.130578e-14, 6.110372e-14, 5.973535e-14, 
    5.979981e-14, 6.002395e-14, 5.991734e-14, 6.022218e-14, 6.029712e-14, 
    6.035806e-14, 6.043587e-14, 6.04443e-14, 6.049038e-14, 6.041485e-14, 
    6.048742e-14, 6.021272e-14, 6.033553e-14, 5.999839e-14, 6.008048e-14, 
    6.004273e-14, 6.000129e-14, 6.012916e-14, 6.026523e-14, 6.02682e-14, 
    6.03118e-14, 6.04345e-14, 6.022341e-14, 6.087652e-14, 6.047334e-14, 
    5.987008e-14, 5.999406e-14, 6.001184e-14, 5.996381e-14, 6.028961e-14, 
    6.017161e-14, 6.048927e-14, 6.040348e-14, 6.054404e-14, 6.04742e-14, 
    6.046392e-14, 6.03742e-14, 6.03183e-14, 6.017702e-14, 6.0062e-14, 
    5.997079e-14, 5.9992e-14, 6.00922e-14, 6.027356e-14, 6.044503e-14, 
    6.040748e-14, 6.053336e-14, 6.020009e-14, 6.033988e-14, 6.028584e-14, 
    6.042671e-14, 6.011797e-14, 6.038073e-14, 6.005073e-14, 6.007969e-14, 
    6.016928e-14, 6.034932e-14, 6.038921e-14, 6.043169e-14, 6.04055e-14, 
    6.027818e-14, 6.025734e-14, 6.016712e-14, 6.014216e-14, 6.007339e-14, 
    6.001642e-14, 6.006846e-14, 6.012309e-14, 6.027826e-14, 6.041795e-14, 
    6.057016e-14, 6.060742e-14, 6.078491e-14, 6.064035e-14, 6.087875e-14, 
    6.067596e-14, 6.102693e-14, 6.039604e-14, 6.067012e-14, 6.017337e-14, 
    6.022696e-14, 6.032379e-14, 6.054583e-14, 6.042606e-14, 6.056615e-14, 
    6.025653e-14, 6.009562e-14, 6.005404e-14, 5.997632e-14, 6.005582e-14, 
    6.004936e-14, 6.012539e-14, 6.010097e-14, 6.028341e-14, 6.018543e-14, 
    6.046365e-14, 6.056506e-14, 6.085122e-14, 6.102639e-14, 6.120461e-14, 
    6.12832e-14, 6.130712e-14, 6.131711e-14 ;

 LITTERC =
  5.976298e-05, 5.976283e-05, 5.976286e-05, 5.976274e-05, 5.976281e-05, 
    5.976273e-05, 5.976295e-05, 5.976282e-05, 5.97629e-05, 5.976297e-05, 
    5.976251e-05, 5.976273e-05, 5.976227e-05, 5.976242e-05, 5.976206e-05, 
    5.97623e-05, 5.976201e-05, 5.976206e-05, 5.97619e-05, 5.976194e-05, 
    5.976173e-05, 5.976187e-05, 5.976162e-05, 5.976177e-05, 5.976174e-05, 
    5.976188e-05, 5.976269e-05, 5.976254e-05, 5.97627e-05, 5.976267e-05, 
    5.976269e-05, 5.976281e-05, 5.976286e-05, 5.976299e-05, 5.976297e-05, 
    5.976288e-05, 5.976267e-05, 5.976274e-05, 5.976256e-05, 5.976256e-05, 
    5.976236e-05, 5.976245e-05, 5.976212e-05, 5.976221e-05, 5.976194e-05, 
    5.976201e-05, 5.976194e-05, 5.976197e-05, 5.976194e-05, 5.976205e-05, 
    5.9762e-05, 5.976209e-05, 5.976243e-05, 5.976234e-05, 5.976264e-05, 
    5.976282e-05, 5.976294e-05, 5.976303e-05, 5.976302e-05, 5.9763e-05, 
    5.976288e-05, 5.976276e-05, 5.976267e-05, 5.976262e-05, 5.976256e-05, 
    5.976239e-05, 5.97623e-05, 5.97621e-05, 5.976214e-05, 5.976207e-05, 
    5.976202e-05, 5.976192e-05, 5.976193e-05, 5.976189e-05, 5.976208e-05, 
    5.976195e-05, 5.976216e-05, 5.97621e-05, 5.976255e-05, 5.976272e-05, 
    5.976279e-05, 5.976285e-05, 5.976301e-05, 5.97629e-05, 5.976294e-05, 
    5.976284e-05, 5.976278e-05, 5.976281e-05, 5.976262e-05, 5.976269e-05, 
    5.97623e-05, 5.976247e-05, 5.976202e-05, 5.976213e-05, 5.9762e-05, 
    5.976206e-05, 5.976195e-05, 5.976205e-05, 5.976187e-05, 5.976183e-05, 
    5.976186e-05, 5.976176e-05, 5.976206e-05, 5.976194e-05, 5.976281e-05, 
    5.976281e-05, 5.976278e-05, 5.976289e-05, 5.976289e-05, 5.976299e-05, 
    5.97629e-05, 5.976287e-05, 5.976278e-05, 5.976272e-05, 5.976267e-05, 
    5.976255e-05, 5.976243e-05, 5.976225e-05, 5.976212e-05, 5.976204e-05, 
    5.976209e-05, 5.976204e-05, 5.97621e-05, 5.976212e-05, 5.976185e-05, 
    5.9762e-05, 5.976178e-05, 5.976179e-05, 5.976189e-05, 5.976179e-05, 
    5.97628e-05, 5.976283e-05, 5.976293e-05, 5.976285e-05, 5.9763e-05, 
    5.976292e-05, 5.976287e-05, 5.976269e-05, 5.976265e-05, 5.976261e-05, 
    5.976254e-05, 5.976245e-05, 5.976229e-05, 5.976214e-05, 5.976201e-05, 
    5.976202e-05, 5.976202e-05, 5.976199e-05, 5.976206e-05, 5.976198e-05, 
    5.976197e-05, 5.9762e-05, 5.976179e-05, 5.976185e-05, 5.976179e-05, 
    5.976183e-05, 5.976282e-05, 5.976277e-05, 5.97628e-05, 5.976275e-05, 
    5.976278e-05, 5.976263e-05, 5.976258e-05, 5.976236e-05, 5.976245e-05, 
    5.976231e-05, 5.976243e-05, 5.976241e-05, 5.97623e-05, 5.976243e-05, 
    5.976215e-05, 5.976234e-05, 5.976199e-05, 5.976218e-05, 5.976198e-05, 
    5.976201e-05, 5.976195e-05, 5.97619e-05, 5.976183e-05, 5.976171e-05, 
    5.976174e-05, 5.976163e-05, 5.97627e-05, 5.976263e-05, 5.976264e-05, 
    5.976257e-05, 5.976253e-05, 5.976242e-05, 5.976225e-05, 5.976231e-05, 
    5.976219e-05, 5.976217e-05, 5.976235e-05, 5.976223e-05, 5.976259e-05, 
    5.976254e-05, 5.976257e-05, 5.976269e-05, 5.976229e-05, 5.97625e-05, 
    5.976212e-05, 5.976223e-05, 5.976191e-05, 5.976207e-05, 5.976175e-05, 
    5.976162e-05, 5.976149e-05, 5.976134e-05, 5.97626e-05, 5.976265e-05, 
    5.976257e-05, 5.976246e-05, 5.976236e-05, 5.976222e-05, 5.976221e-05, 
    5.976219e-05, 5.976212e-05, 5.976207e-05, 5.976218e-05, 5.976205e-05, 
    5.976252e-05, 5.976228e-05, 5.976266e-05, 5.976254e-05, 5.976246e-05, 
    5.97625e-05, 5.976232e-05, 5.976227e-05, 5.97621e-05, 5.976219e-05, 
    5.976165e-05, 5.976189e-05, 5.976123e-05, 5.976141e-05, 5.976266e-05, 
    5.97626e-05, 5.97624e-05, 5.976249e-05, 5.976222e-05, 5.976215e-05, 
    5.976209e-05, 5.976202e-05, 5.976201e-05, 5.976197e-05, 5.976204e-05, 
    5.976198e-05, 5.976222e-05, 5.976211e-05, 5.976242e-05, 5.976234e-05, 
    5.976238e-05, 5.976242e-05, 5.97623e-05, 5.976218e-05, 5.976217e-05, 
    5.976213e-05, 5.976202e-05, 5.976222e-05, 5.976162e-05, 5.976199e-05, 
    5.976254e-05, 5.976242e-05, 5.976241e-05, 5.976245e-05, 5.976215e-05, 
    5.976226e-05, 5.976197e-05, 5.976205e-05, 5.976192e-05, 5.976199e-05, 
    5.976199e-05, 5.976208e-05, 5.976213e-05, 5.976226e-05, 5.976236e-05, 
    5.976245e-05, 5.976243e-05, 5.976233e-05, 5.976217e-05, 5.976201e-05, 
    5.976205e-05, 5.976193e-05, 5.976223e-05, 5.976211e-05, 5.976216e-05, 
    5.976203e-05, 5.976231e-05, 5.976207e-05, 5.976237e-05, 5.976235e-05, 
    5.976226e-05, 5.97621e-05, 5.976206e-05, 5.976202e-05, 5.976205e-05, 
    5.976217e-05, 5.976218e-05, 5.976227e-05, 5.976229e-05, 5.976235e-05, 
    5.97624e-05, 5.976235e-05, 5.976231e-05, 5.976217e-05, 5.976204e-05, 
    5.97619e-05, 5.976186e-05, 5.97617e-05, 5.976183e-05, 5.976162e-05, 
    5.97618e-05, 5.976148e-05, 5.976206e-05, 5.976181e-05, 5.976226e-05, 
    5.976221e-05, 5.976212e-05, 5.976192e-05, 5.976203e-05, 5.97619e-05, 
    5.976218e-05, 5.976233e-05, 5.976237e-05, 5.976244e-05, 5.976237e-05, 
    5.976237e-05, 5.97623e-05, 5.976233e-05, 5.976216e-05, 5.976225e-05, 
    5.976199e-05, 5.97619e-05, 5.976164e-05, 5.976149e-05, 5.976132e-05, 
    5.976125e-05, 5.976123e-05, 5.976122e-05 ;

 LITTERC_HR =
  9.581084e-13, 9.607331e-13, 9.602232e-13, 9.623386e-13, 9.611656e-13, 
    9.625504e-13, 9.58641e-13, 9.608369e-13, 9.594355e-13, 9.583453e-13, 
    9.664388e-13, 9.62433e-13, 9.705987e-13, 9.680471e-13, 9.744543e-13, 
    9.702012e-13, 9.753114e-13, 9.743327e-13, 9.772797e-13, 9.764358e-13, 
    9.802e-13, 9.776691e-13, 9.82151e-13, 9.795963e-13, 9.799957e-13, 
    9.775854e-13, 9.632404e-13, 9.659401e-13, 9.630803e-13, 9.634654e-13, 
    9.632928e-13, 9.611896e-13, 9.601286e-13, 9.579082e-13, 9.583117e-13, 
    9.599426e-13, 9.636387e-13, 9.623851e-13, 9.655452e-13, 9.65474e-13, 
    9.689881e-13, 9.674041e-13, 9.733056e-13, 9.716297e-13, 9.764711e-13, 
    9.752541e-13, 9.764137e-13, 9.760622e-13, 9.764183e-13, 9.746334e-13, 
    9.753981e-13, 9.738274e-13, 9.677006e-13, 9.695021e-13, 9.641258e-13, 
    9.608874e-13, 9.587372e-13, 9.572099e-13, 9.574259e-13, 9.578373e-13, 
    9.599522e-13, 9.619403e-13, 9.634543e-13, 9.644665e-13, 9.654637e-13, 
    9.684779e-13, 9.700742e-13, 9.736439e-13, 9.730008e-13, 9.740908e-13, 
    9.75133e-13, 9.768808e-13, 9.765933e-13, 9.773628e-13, 9.740626e-13, 
    9.762561e-13, 9.726342e-13, 9.736252e-13, 9.657315e-13, 9.627235e-13, 
    9.614413e-13, 9.603211e-13, 9.575918e-13, 9.594766e-13, 9.587336e-13, 
    9.605016e-13, 9.616241e-13, 9.610692e-13, 9.644942e-13, 9.631629e-13, 
    9.701687e-13, 9.671529e-13, 9.750114e-13, 9.731329e-13, 9.754617e-13, 
    9.742737e-13, 9.763087e-13, 9.744773e-13, 9.776495e-13, 9.783394e-13, 
    9.778679e-13, 9.796799e-13, 9.743756e-13, 9.764134e-13, 9.610535e-13, 
    9.611439e-13, 9.61566e-13, 9.597106e-13, 9.595973e-13, 9.578971e-13, 
    9.594102e-13, 9.600541e-13, 9.616895e-13, 9.626558e-13, 9.635744e-13, 
    9.655932e-13, 9.678459e-13, 9.709942e-13, 9.732547e-13, 9.747688e-13, 
    9.738407e-13, 9.7466e-13, 9.737439e-13, 9.733145e-13, 9.780807e-13, 
    9.754051e-13, 9.794193e-13, 9.791974e-13, 9.77381e-13, 9.792225e-13, 
    9.612076e-13, 9.606866e-13, 9.588764e-13, 9.602932e-13, 9.577119e-13, 
    9.591566e-13, 9.599868e-13, 9.6319e-13, 9.638942e-13, 9.64546e-13, 
    9.658337e-13, 9.674852e-13, 9.7038e-13, 9.728972e-13, 9.751938e-13, 
    9.750256e-13, 9.750848e-13, 9.755972e-13, 9.743272e-13, 9.758057e-13, 
    9.760535e-13, 9.754052e-13, 9.791677e-13, 9.780933e-13, 9.791927e-13, 
    9.784933e-13, 9.608561e-13, 9.617326e-13, 9.61259e-13, 9.621495e-13, 
    9.615219e-13, 9.643109e-13, 9.651466e-13, 9.690552e-13, 9.674525e-13, 
    9.700038e-13, 9.67712e-13, 9.681181e-13, 9.700857e-13, 9.678362e-13, 
    9.727578e-13, 9.694207e-13, 9.756172e-13, 9.722864e-13, 9.758256e-13, 
    9.751838e-13, 9.762469e-13, 9.771981e-13, 9.783952e-13, 9.806018e-13, 
    9.800911e-13, 9.819359e-13, 9.630393e-13, 9.641754e-13, 9.640759e-13, 
    9.652648e-13, 9.661435e-13, 9.680481e-13, 9.710999e-13, 9.69953e-13, 
    9.720591e-13, 9.724815e-13, 9.692819e-13, 9.712463e-13, 9.649358e-13, 
    9.659555e-13, 9.653489e-13, 9.631287e-13, 9.702164e-13, 9.665804e-13, 
    9.732919e-13, 9.713247e-13, 9.770625e-13, 9.742096e-13, 9.798098e-13, 
    9.821989e-13, 9.844485e-13, 9.870719e-13, 9.647957e-13, 9.64024e-13, 
    9.654062e-13, 9.673165e-13, 9.690897e-13, 9.714446e-13, 9.716858e-13, 
    9.721266e-13, 9.732687e-13, 9.742284e-13, 9.722653e-13, 9.74469e-13, 
    9.661908e-13, 9.705321e-13, 9.637317e-13, 9.657801e-13, 9.672042e-13, 
    9.665802e-13, 9.698219e-13, 9.705853e-13, 9.736852e-13, 9.720834e-13, 
    9.816089e-13, 9.773983e-13, 9.890697e-13, 9.858125e-13, 9.637543e-13, 
    9.647933e-13, 9.684067e-13, 9.666881e-13, 9.716021e-13, 9.728103e-13, 
    9.737926e-13, 9.750469e-13, 9.751826e-13, 9.759256e-13, 9.747079e-13, 
    9.758778e-13, 9.714496e-13, 9.734293e-13, 9.679946e-13, 9.693178e-13, 
    9.687094e-13, 9.680413e-13, 9.701026e-13, 9.72296e-13, 9.72344e-13, 
    9.730467e-13, 9.750247e-13, 9.71622e-13, 9.821501e-13, 9.756509e-13, 
    9.659261e-13, 9.679249e-13, 9.682114e-13, 9.674372e-13, 9.726891e-13, 
    9.70787e-13, 9.759076e-13, 9.745247e-13, 9.767905e-13, 9.756648e-13, 
    9.75499e-13, 9.740527e-13, 9.731516e-13, 9.708741e-13, 9.6902e-13, 
    9.675496e-13, 9.678916e-13, 9.695067e-13, 9.724305e-13, 9.751945e-13, 
    9.745891e-13, 9.766184e-13, 9.71246e-13, 9.734994e-13, 9.726283e-13, 
    9.748992e-13, 9.699222e-13, 9.741579e-13, 9.688383e-13, 9.693053e-13, 
    9.707492e-13, 9.736515e-13, 9.742946e-13, 9.749795e-13, 9.745571e-13, 
    9.725048e-13, 9.721689e-13, 9.707144e-13, 9.703122e-13, 9.692037e-13, 
    9.682851e-13, 9.691241e-13, 9.700048e-13, 9.72506e-13, 9.747579e-13, 
    9.772116e-13, 9.778121e-13, 9.806733e-13, 9.783431e-13, 9.821861e-13, 
    9.78917e-13, 9.845746e-13, 9.744047e-13, 9.788228e-13, 9.708152e-13, 
    9.716791e-13, 9.732402e-13, 9.768193e-13, 9.748886e-13, 9.77147e-13, 
    9.721557e-13, 9.695619e-13, 9.688916e-13, 9.676388e-13, 9.689203e-13, 
    9.688162e-13, 9.700419e-13, 9.696481e-13, 9.725891e-13, 9.710097e-13, 
    9.754946e-13, 9.771293e-13, 9.817422e-13, 9.845659e-13, 9.874389e-13, 
    9.887056e-13, 9.890913e-13, 9.892524e-13 ;

 LITTERC_LOSS =
  1.774407e-12, 1.779268e-12, 1.778324e-12, 1.782242e-12, 1.780069e-12, 
    1.782634e-12, 1.775394e-12, 1.77946e-12, 1.776865e-12, 1.774846e-12, 
    1.789835e-12, 1.782416e-12, 1.79754e-12, 1.792814e-12, 1.80468e-12, 
    1.796803e-12, 1.806267e-12, 1.804455e-12, 1.809913e-12, 1.80835e-12, 
    1.815321e-12, 1.810634e-12, 1.818934e-12, 1.814203e-12, 1.814943e-12, 
    1.810479e-12, 1.783912e-12, 1.788912e-12, 1.783615e-12, 1.784328e-12, 
    1.784009e-12, 1.780113e-12, 1.778148e-12, 1.774037e-12, 1.774784e-12, 
    1.777804e-12, 1.784649e-12, 1.782328e-12, 1.78818e-12, 1.788048e-12, 
    1.794557e-12, 1.791623e-12, 1.802553e-12, 1.799449e-12, 1.808415e-12, 
    1.806161e-12, 1.808309e-12, 1.807658e-12, 1.808317e-12, 1.805012e-12, 
    1.806428e-12, 1.803519e-12, 1.792172e-12, 1.795509e-12, 1.785551e-12, 
    1.779554e-12, 1.775572e-12, 1.772743e-12, 1.773143e-12, 1.773905e-12, 
    1.777822e-12, 1.781504e-12, 1.784308e-12, 1.786183e-12, 1.788029e-12, 
    1.793612e-12, 1.796568e-12, 1.803179e-12, 1.801988e-12, 1.804007e-12, 
    1.805937e-12, 1.809174e-12, 1.808641e-12, 1.810067e-12, 1.803955e-12, 
    1.808017e-12, 1.801309e-12, 1.803144e-12, 1.788525e-12, 1.782954e-12, 
    1.78058e-12, 1.778505e-12, 1.77345e-12, 1.776941e-12, 1.775565e-12, 
    1.77884e-12, 1.780918e-12, 1.779891e-12, 1.786234e-12, 1.783768e-12, 
    1.796743e-12, 1.791158e-12, 1.805712e-12, 1.802233e-12, 1.806546e-12, 
    1.804346e-12, 1.808114e-12, 1.804723e-12, 1.810598e-12, 1.811875e-12, 
    1.811002e-12, 1.814358e-12, 1.804534e-12, 1.808308e-12, 1.779862e-12, 
    1.780029e-12, 1.780811e-12, 1.777374e-12, 1.777165e-12, 1.774016e-12, 
    1.776818e-12, 1.778011e-12, 1.781039e-12, 1.782829e-12, 1.78453e-12, 
    1.788269e-12, 1.792441e-12, 1.798272e-12, 1.802458e-12, 1.805263e-12, 
    1.803544e-12, 1.805061e-12, 1.803364e-12, 1.802569e-12, 1.811396e-12, 
    1.806441e-12, 1.813875e-12, 1.813464e-12, 1.8101e-12, 1.813511e-12, 
    1.780147e-12, 1.779182e-12, 1.775829e-12, 1.778453e-12, 1.773673e-12, 
    1.776348e-12, 1.777886e-12, 1.783818e-12, 1.785123e-12, 1.78633e-12, 
    1.788715e-12, 1.791773e-12, 1.797134e-12, 1.801796e-12, 1.80605e-12, 
    1.805738e-12, 1.805848e-12, 1.806797e-12, 1.804445e-12, 1.807183e-12, 
    1.807642e-12, 1.806441e-12, 1.813409e-12, 1.81142e-12, 1.813456e-12, 
    1.81216e-12, 1.779496e-12, 1.781119e-12, 1.780242e-12, 1.781891e-12, 
    1.780729e-12, 1.785894e-12, 1.787442e-12, 1.794681e-12, 1.791713e-12, 
    1.796438e-12, 1.792193e-12, 1.792945e-12, 1.796589e-12, 1.792423e-12, 
    1.801538e-12, 1.795358e-12, 1.806834e-12, 1.800665e-12, 1.80722e-12, 
    1.806031e-12, 1.808e-12, 1.809762e-12, 1.811979e-12, 1.816065e-12, 
    1.815119e-12, 1.818536e-12, 1.783539e-12, 1.785643e-12, 1.785459e-12, 
    1.787661e-12, 1.789288e-12, 1.792816e-12, 1.798468e-12, 1.796343e-12, 
    1.800244e-12, 1.801026e-12, 1.795101e-12, 1.798739e-12, 1.787052e-12, 
    1.78894e-12, 1.787817e-12, 1.783705e-12, 1.796831e-12, 1.790098e-12, 
    1.802527e-12, 1.798884e-12, 1.80951e-12, 1.804227e-12, 1.814598e-12, 
    1.819023e-12, 1.82319e-12, 1.828048e-12, 1.786792e-12, 1.785363e-12, 
    1.787923e-12, 1.791461e-12, 1.794745e-12, 1.799106e-12, 1.799553e-12, 
    1.800369e-12, 1.802484e-12, 1.804262e-12, 1.800626e-12, 1.804707e-12, 
    1.789376e-12, 1.797416e-12, 1.784822e-12, 1.788615e-12, 1.791253e-12, 
    1.790097e-12, 1.796101e-12, 1.797515e-12, 1.803256e-12, 1.800289e-12, 
    1.817931e-12, 1.810132e-12, 1.831748e-12, 1.825716e-12, 1.784863e-12, 
    1.786788e-12, 1.79348e-12, 1.790297e-12, 1.799398e-12, 1.801635e-12, 
    1.803455e-12, 1.805777e-12, 1.806029e-12, 1.807405e-12, 1.80515e-12, 
    1.807316e-12, 1.799115e-12, 1.802782e-12, 1.792717e-12, 1.795167e-12, 
    1.79404e-12, 1.792803e-12, 1.796621e-12, 1.800683e-12, 1.800772e-12, 
    1.802073e-12, 1.805737e-12, 1.799435e-12, 1.818933e-12, 1.806896e-12, 
    1.788886e-12, 1.792587e-12, 1.793118e-12, 1.791684e-12, 1.801411e-12, 
    1.797888e-12, 1.807372e-12, 1.804811e-12, 1.809007e-12, 1.806922e-12, 
    1.806615e-12, 1.803936e-12, 1.802267e-12, 1.798049e-12, 1.794616e-12, 
    1.791892e-12, 1.792526e-12, 1.795517e-12, 1.800932e-12, 1.806051e-12, 
    1.80493e-12, 1.808688e-12, 1.798738e-12, 1.802912e-12, 1.801298e-12, 
    1.805504e-12, 1.796287e-12, 1.804131e-12, 1.794279e-12, 1.795144e-12, 
    1.797818e-12, 1.803193e-12, 1.804384e-12, 1.805653e-12, 1.804871e-12, 
    1.80107e-12, 1.800447e-12, 1.797754e-12, 1.797009e-12, 1.794956e-12, 
    1.793255e-12, 1.794808e-12, 1.796439e-12, 1.801072e-12, 1.805242e-12, 
    1.809787e-12, 1.810899e-12, 1.816198e-12, 1.811882e-12, 1.818999e-12, 
    1.812945e-12, 1.823423e-12, 1.804588e-12, 1.812771e-12, 1.79794e-12, 
    1.79954e-12, 1.802431e-12, 1.80906e-12, 1.805484e-12, 1.809667e-12, 
    1.800423e-12, 1.795619e-12, 1.794378e-12, 1.792058e-12, 1.794431e-12, 
    1.794238e-12, 1.796508e-12, 1.795779e-12, 1.801226e-12, 1.798301e-12, 
    1.806607e-12, 1.809634e-12, 1.818178e-12, 1.823407e-12, 1.828728e-12, 
    1.831074e-12, 1.831788e-12, 1.832086e-12 ;

 LIVECROOTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVECROOTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 LIVESTEMN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 MEG_acetaldehyde =
  1.676205e-18, 1.676468e-18, 1.676418e-18, 1.676627e-18, 1.676513e-18, 
    1.676648e-18, 1.676261e-18, 1.676476e-18, 1.67634e-18, 1.676232e-18, 
    1.677027e-18, 1.676637e-18, 1.677455e-18, 1.677202e-18, 1.677845e-18, 
    1.677412e-18, 1.677933e-18, 1.677838e-18, 1.678138e-18, 1.678052e-18, 
    1.678426e-18, 1.678178e-18, 1.678629e-18, 1.67837e-18, 1.678408e-18, 
    1.678169e-18, 1.67672e-18, 1.676977e-18, 1.676704e-18, 1.676741e-18, 
    1.676726e-18, 1.676514e-18, 1.676403e-18, 1.676189e-18, 1.676229e-18, 
    1.676388e-18, 1.676758e-18, 1.676635e-18, 1.676953e-18, 1.676946e-18, 
    1.677297e-18, 1.677139e-18, 1.677733e-18, 1.677565e-18, 1.678056e-18, 
    1.677932e-18, 1.678049e-18, 1.678014e-18, 1.67805e-18, 1.677868e-18, 
    1.677945e-18, 1.677787e-18, 1.677167e-18, 1.677348e-18, 1.676808e-18, 
    1.676476e-18, 1.676269e-18, 1.676119e-18, 1.67614e-18, 1.676179e-18, 
    1.676389e-18, 1.676591e-18, 1.676743e-18, 1.676845e-18, 1.676945e-18, 
    1.677236e-18, 1.677402e-18, 1.677765e-18, 1.677704e-18, 1.677811e-18, 
    1.677919e-18, 1.678096e-18, 1.678068e-18, 1.678145e-18, 1.677811e-18, 
    1.678031e-18, 1.677668e-18, 1.677767e-18, 1.676955e-18, 1.676669e-18, 
    1.676533e-18, 1.676427e-18, 1.676156e-18, 1.676342e-18, 1.676268e-18, 
    1.676448e-18, 1.676559e-18, 1.676505e-18, 1.676847e-18, 1.676713e-18, 
    1.677412e-18, 1.677111e-18, 1.677907e-18, 1.677717e-18, 1.677953e-18, 
    1.677833e-18, 1.678037e-18, 1.677854e-18, 1.678175e-18, 1.678242e-18, 
    1.678196e-18, 1.678382e-18, 1.677843e-18, 1.678048e-18, 1.676502e-18, 
    1.676511e-18, 1.676554e-18, 1.676365e-18, 1.676355e-18, 1.676187e-18, 
    1.676338e-18, 1.6764e-18, 1.676567e-18, 1.676662e-18, 1.676754e-18, 
    1.676956e-18, 1.67718e-18, 1.677497e-18, 1.677729e-18, 1.677883e-18, 
    1.67779e-18, 1.677872e-18, 1.677779e-18, 1.677737e-18, 1.678216e-18, 
    1.677945e-18, 1.678355e-18, 1.678333e-18, 1.678146e-18, 1.678335e-18, 
    1.676517e-18, 1.676466e-18, 1.676284e-18, 1.676427e-18, 1.676169e-18, 
    1.676311e-18, 1.676391e-18, 1.676712e-18, 1.676787e-18, 1.676851e-18, 
    1.676981e-18, 1.677147e-18, 1.677436e-18, 1.677691e-18, 1.677926e-18, 
    1.67791e-18, 1.677915e-18, 1.677966e-18, 1.677838e-18, 1.677987e-18, 
    1.678011e-18, 1.677947e-18, 1.67833e-18, 1.67822e-18, 1.678332e-18, 
    1.678261e-18, 1.676484e-18, 1.67657e-18, 1.676523e-18, 1.676611e-18, 
    1.676548e-18, 1.676824e-18, 1.676906e-18, 1.677299e-18, 1.677142e-18, 
    1.677397e-18, 1.67717e-18, 1.677209e-18, 1.677398e-18, 1.677183e-18, 
    1.677673e-18, 1.677334e-18, 1.677968e-18, 1.677622e-18, 1.67799e-18, 
    1.677925e-18, 1.678033e-18, 1.678128e-18, 1.678251e-18, 1.678472e-18, 
    1.678422e-18, 1.67861e-18, 1.676701e-18, 1.676812e-18, 1.676806e-18, 
    1.676924e-18, 1.677011e-18, 1.677204e-18, 1.67751e-18, 1.677396e-18, 
    1.677609e-18, 1.677651e-18, 1.677329e-18, 1.677523e-18, 1.676889e-18, 
    1.676988e-18, 1.676931e-18, 1.676708e-18, 1.677418e-18, 1.677051e-18, 
    1.677732e-18, 1.677533e-18, 1.678114e-18, 1.677822e-18, 1.678393e-18, 
    1.678629e-18, 1.678868e-18, 1.679129e-18, 1.676876e-18, 1.676801e-18, 
    1.676939e-18, 1.677125e-18, 1.677308e-18, 1.677545e-18, 1.677571e-18, 
    1.677615e-18, 1.677732e-18, 1.677828e-18, 1.677625e-18, 1.677853e-18, 
    1.677004e-18, 1.677451e-18, 1.676769e-18, 1.67697e-18, 1.677116e-18, 
    1.677055e-18, 1.677384e-18, 1.67746e-18, 1.67777e-18, 1.677612e-18, 
    1.678568e-18, 1.678144e-18, 1.679339e-18, 1.679002e-18, 1.676773e-18, 
    1.676878e-18, 1.677237e-18, 1.677066e-18, 1.677563e-18, 1.677683e-18, 
    1.677785e-18, 1.677909e-18, 1.677925e-18, 1.677999e-18, 1.677877e-18, 
    1.677995e-18, 1.677545e-18, 1.677747e-18, 1.6772e-18, 1.677331e-18, 
    1.677271e-18, 1.677204e-18, 1.677412e-18, 1.677628e-18, 1.677638e-18, 
    1.677706e-18, 1.677889e-18, 1.677565e-18, 1.678613e-18, 1.677956e-18, 
    1.676991e-18, 1.677185e-18, 1.67722e-18, 1.677143e-18, 1.677671e-18, 
    1.677479e-18, 1.677998e-18, 1.677859e-18, 1.678088e-18, 1.677974e-18, 
    1.677956e-18, 1.677811e-18, 1.677718e-18, 1.677487e-18, 1.6773e-18, 
    1.677155e-18, 1.677189e-18, 1.677349e-18, 1.677642e-18, 1.677924e-18, 
    1.677861e-18, 1.678071e-18, 1.677526e-18, 1.677752e-18, 1.677663e-18, 
    1.677896e-18, 1.677392e-18, 1.677805e-18, 1.677285e-18, 1.677331e-18, 
    1.677475e-18, 1.677763e-18, 1.677835e-18, 1.677902e-18, 1.677862e-18, 
    1.67765e-18, 1.677618e-18, 1.677473e-18, 1.67743e-18, 1.677321e-18, 
    1.677229e-18, 1.677312e-18, 1.677399e-18, 1.677653e-18, 1.677879e-18, 
    1.678129e-18, 1.678192e-18, 1.678471e-18, 1.678236e-18, 1.678616e-18, 
    1.678282e-18, 1.678866e-18, 1.677836e-18, 1.678283e-18, 1.677484e-18, 
    1.677571e-18, 1.677723e-18, 1.678084e-18, 1.677895e-18, 1.678119e-18, 
    1.677617e-18, 1.677352e-18, 1.67729e-18, 1.677163e-18, 1.677292e-18, 
    1.677282e-18, 1.677406e-18, 1.677366e-18, 1.677661e-18, 1.677503e-18, 
    1.677955e-18, 1.678118e-18, 1.678588e-18, 1.678874e-18, 1.679174e-18, 
    1.679304e-18, 1.679344e-18, 1.67936e-18 ;

 MEG_acetic_acid =
  2.514308e-19, 2.514702e-19, 2.514627e-19, 2.514941e-19, 2.514769e-19, 
    2.514973e-19, 2.514391e-19, 2.514714e-19, 2.51451e-19, 2.514348e-19, 
    2.515541e-19, 2.514955e-19, 2.516182e-19, 2.515803e-19, 2.516767e-19, 
    2.516119e-19, 2.5169e-19, 2.516756e-19, 2.517207e-19, 2.517078e-19, 
    2.517639e-19, 2.517266e-19, 2.517944e-19, 2.517555e-19, 2.517613e-19, 
    2.517253e-19, 2.51508e-19, 2.515465e-19, 2.515056e-19, 2.515111e-19, 
    2.515088e-19, 2.51477e-19, 2.514605e-19, 2.514283e-19, 2.514343e-19, 
    2.514582e-19, 2.515136e-19, 2.514953e-19, 2.51543e-19, 2.515419e-19, 
    2.515945e-19, 2.515708e-19, 2.5166e-19, 2.516348e-19, 2.517084e-19, 
    2.516897e-19, 2.517074e-19, 2.517021e-19, 2.517074e-19, 2.516801e-19, 
    2.516918e-19, 2.51668e-19, 2.515751e-19, 2.516021e-19, 2.515212e-19, 
    2.514714e-19, 2.514404e-19, 2.514178e-19, 2.51421e-19, 2.514269e-19, 
    2.514584e-19, 2.514886e-19, 2.515115e-19, 2.515267e-19, 2.515417e-19, 
    2.515854e-19, 2.516103e-19, 2.516647e-19, 2.516555e-19, 2.516716e-19, 
    2.516879e-19, 2.517144e-19, 2.517101e-19, 2.517217e-19, 2.516717e-19, 
    2.517046e-19, 2.516502e-19, 2.51665e-19, 2.515432e-19, 2.515004e-19, 
    2.514799e-19, 2.51464e-19, 2.514234e-19, 2.514513e-19, 2.514402e-19, 
    2.514671e-19, 2.514838e-19, 2.514757e-19, 2.515271e-19, 2.51507e-19, 
    2.516117e-19, 2.515666e-19, 2.51686e-19, 2.516575e-19, 2.516929e-19, 
    2.51675e-19, 2.517056e-19, 2.51678e-19, 2.517262e-19, 2.517364e-19, 
    2.517293e-19, 2.517572e-19, 2.516764e-19, 2.517071e-19, 2.514753e-19, 
    2.514767e-19, 2.514831e-19, 2.514547e-19, 2.514532e-19, 2.51428e-19, 
    2.514506e-19, 2.514601e-19, 2.51485e-19, 2.514993e-19, 2.515131e-19, 
    2.515434e-19, 2.515769e-19, 2.516246e-19, 2.516593e-19, 2.516825e-19, 
    2.516684e-19, 2.516808e-19, 2.516669e-19, 2.516605e-19, 2.517324e-19, 
    2.516917e-19, 2.517532e-19, 2.517499e-19, 2.517218e-19, 2.517503e-19, 
    2.514776e-19, 2.5147e-19, 2.514426e-19, 2.51464e-19, 2.514253e-19, 
    2.514466e-19, 2.514587e-19, 2.515069e-19, 2.515181e-19, 2.515276e-19, 
    2.515472e-19, 2.51572e-19, 2.516154e-19, 2.516536e-19, 2.51689e-19, 
    2.516864e-19, 2.516873e-19, 2.516949e-19, 2.516757e-19, 2.516981e-19, 
    2.517016e-19, 2.51692e-19, 2.517494e-19, 2.517331e-19, 2.517498e-19, 
    2.517392e-19, 2.514725e-19, 2.514855e-19, 2.514784e-19, 2.514916e-19, 
    2.514821e-19, 2.515235e-19, 2.51536e-19, 2.515949e-19, 2.515713e-19, 
    2.516096e-19, 2.515754e-19, 2.515813e-19, 2.516097e-19, 2.515774e-19, 
    2.51651e-19, 2.516001e-19, 2.516952e-19, 2.516433e-19, 2.516984e-19, 
    2.516888e-19, 2.51705e-19, 2.517192e-19, 2.517376e-19, 2.517708e-19, 
    2.517633e-19, 2.517915e-19, 2.515052e-19, 2.515218e-19, 2.515208e-19, 
    2.515386e-19, 2.515517e-19, 2.515806e-19, 2.516265e-19, 2.516094e-19, 
    2.516413e-19, 2.516476e-19, 2.515993e-19, 2.516285e-19, 2.515333e-19, 
    2.515482e-19, 2.515397e-19, 2.515062e-19, 2.516127e-19, 2.515576e-19, 
    2.516598e-19, 2.5163e-19, 2.517171e-19, 2.516732e-19, 2.51759e-19, 
    2.517944e-19, 2.518301e-19, 2.518693e-19, 2.515315e-19, 2.515201e-19, 
    2.515409e-19, 2.515688e-19, 2.515961e-19, 2.516317e-19, 2.516357e-19, 
    2.516422e-19, 2.516597e-19, 2.516743e-19, 2.516438e-19, 2.516779e-19, 
    2.515506e-19, 2.516176e-19, 2.515153e-19, 2.515454e-19, 2.515674e-19, 
    2.515582e-19, 2.516076e-19, 2.51619e-19, 2.516655e-19, 2.516417e-19, 
    2.517852e-19, 2.517215e-19, 2.519008e-19, 2.518502e-19, 2.51516e-19, 
    2.515316e-19, 2.515855e-19, 2.515599e-19, 2.516344e-19, 2.516525e-19, 
    2.516677e-19, 2.516863e-19, 2.516887e-19, 2.516998e-19, 2.516816e-19, 
    2.516993e-19, 2.516318e-19, 2.51662e-19, 2.515799e-19, 2.515996e-19, 
    2.515907e-19, 2.515806e-19, 2.516117e-19, 2.516441e-19, 2.516456e-19, 
    2.516559e-19, 2.516834e-19, 2.516347e-19, 2.51792e-19, 2.516933e-19, 
    2.515487e-19, 2.515778e-19, 2.515829e-19, 2.515715e-19, 2.516507e-19, 
    2.516218e-19, 2.516997e-19, 2.516788e-19, 2.517132e-19, 2.51696e-19, 
    2.516935e-19, 2.516716e-19, 2.516578e-19, 2.51623e-19, 2.51595e-19, 
    2.515732e-19, 2.515783e-19, 2.516023e-19, 2.516463e-19, 2.516886e-19, 
    2.516792e-19, 2.517106e-19, 2.516289e-19, 2.516627e-19, 2.516494e-19, 
    2.516843e-19, 2.516087e-19, 2.516707e-19, 2.515927e-19, 2.515997e-19, 
    2.516213e-19, 2.516645e-19, 2.516753e-19, 2.516853e-19, 2.516793e-19, 
    2.516476e-19, 2.516427e-19, 2.516209e-19, 2.516145e-19, 2.515982e-19, 
    2.515843e-19, 2.515968e-19, 2.516098e-19, 2.516479e-19, 2.516819e-19, 
    2.517193e-19, 2.517288e-19, 2.517706e-19, 2.517355e-19, 2.517924e-19, 
    2.517423e-19, 2.518299e-19, 2.516754e-19, 2.517425e-19, 2.516225e-19, 
    2.516356e-19, 2.516584e-19, 2.517126e-19, 2.516842e-19, 2.517178e-19, 
    2.516426e-19, 2.516027e-19, 2.515934e-19, 2.515744e-19, 2.515939e-19, 
    2.515923e-19, 2.516109e-19, 2.516049e-19, 2.516492e-19, 2.516254e-19, 
    2.516932e-19, 2.517177e-19, 2.517882e-19, 2.518311e-19, 2.518761e-19, 
    2.518955e-19, 2.519015e-19, 2.51904e-19 ;

 MEG_acetone =
  8.435203e-17, 8.436062e-17, 8.435899e-17, 8.436584e-17, 8.43621e-17, 
    8.436654e-17, 8.435385e-17, 8.436089e-17, 8.435644e-17, 8.435291e-17, 
    8.437893e-17, 8.436616e-17, 8.439293e-17, 8.438465e-17, 8.44057e-17, 
    8.439154e-17, 8.44086e-17, 8.440547e-17, 8.441531e-17, 8.44125e-17, 
    8.442475e-17, 8.441661e-17, 8.44314e-17, 8.44229e-17, 8.442416e-17, 
    8.441632e-17, 8.436889e-17, 8.437728e-17, 8.436835e-17, 8.436956e-17, 
    8.436905e-17, 8.436212e-17, 8.435851e-17, 8.435149e-17, 8.43528e-17, 
    8.435802e-17, 8.437011e-17, 8.436611e-17, 8.437651e-17, 8.437628e-17, 
    8.438777e-17, 8.438259e-17, 8.440206e-17, 8.439656e-17, 8.441262e-17, 
    8.440855e-17, 8.44124e-17, 8.441125e-17, 8.441241e-17, 8.440646e-17, 
    8.4409e-17, 8.440381e-17, 8.438352e-17, 8.438942e-17, 8.437175e-17, 
    8.43609e-17, 8.435413e-17, 8.43492e-17, 8.434989e-17, 8.435119e-17, 
    8.435805e-17, 8.436465e-17, 8.436964e-17, 8.437296e-17, 8.437625e-17, 
    8.438578e-17, 8.43912e-17, 8.440309e-17, 8.440108e-17, 8.440459e-17, 
    8.440815e-17, 8.441393e-17, 8.441301e-17, 8.441552e-17, 8.44046e-17, 
    8.44118e-17, 8.439991e-17, 8.440314e-17, 8.437657e-17, 8.436721e-17, 
    8.436275e-17, 8.435928e-17, 8.435041e-17, 8.435651e-17, 8.435409e-17, 
    8.435996e-17, 8.436361e-17, 8.436183e-17, 8.437304e-17, 8.436866e-17, 
    8.439152e-17, 8.438167e-17, 8.440773e-17, 8.440151e-17, 8.440925e-17, 
    8.440532e-17, 8.441201e-17, 8.4406e-17, 8.44165e-17, 8.441873e-17, 
    8.44172e-17, 8.442328e-17, 8.440565e-17, 8.441235e-17, 8.436176e-17, 
    8.436204e-17, 8.436344e-17, 8.435726e-17, 8.435691e-17, 8.435143e-17, 
    8.435636e-17, 8.435842e-17, 8.436387e-17, 8.436699e-17, 8.436999e-17, 
    8.437662e-17, 8.438392e-17, 8.439433e-17, 8.44019e-17, 8.440697e-17, 
    8.44039e-17, 8.44066e-17, 8.440356e-17, 8.440216e-17, 8.441786e-17, 
    8.440898e-17, 8.442241e-17, 8.442168e-17, 8.441556e-17, 8.442177e-17, 
    8.436225e-17, 8.436058e-17, 8.43546e-17, 8.435928e-17, 8.435084e-17, 
    8.435549e-17, 8.435812e-17, 8.436862e-17, 8.437108e-17, 8.437317e-17, 
    8.437744e-17, 8.438284e-17, 8.439231e-17, 8.440067e-17, 8.440838e-17, 
    8.440783e-17, 8.440802e-17, 8.440969e-17, 8.440548e-17, 8.441038e-17, 
    8.441115e-17, 8.440906e-17, 8.442158e-17, 8.441801e-17, 8.442167e-17, 
    8.441935e-17, 8.436114e-17, 8.436397e-17, 8.436243e-17, 8.43653e-17, 
    8.436324e-17, 8.437227e-17, 8.437498e-17, 8.438785e-17, 8.438271e-17, 
    8.439105e-17, 8.43836e-17, 8.438488e-17, 8.439108e-17, 8.438404e-17, 
    8.440009e-17, 8.438899e-17, 8.440975e-17, 8.43984e-17, 8.441045e-17, 
    8.440835e-17, 8.441188e-17, 8.441499e-17, 8.4419e-17, 8.442626e-17, 
    8.44246e-17, 8.443076e-17, 8.436826e-17, 8.437189e-17, 8.437168e-17, 
    8.437557e-17, 8.437841e-17, 8.438472e-17, 8.439474e-17, 8.439101e-17, 
    8.439799e-17, 8.439935e-17, 8.438881e-17, 8.439518e-17, 8.437441e-17, 
    8.437765e-17, 8.43758e-17, 8.436849e-17, 8.439172e-17, 8.437971e-17, 
    8.440201e-17, 8.439551e-17, 8.441453e-17, 8.440495e-17, 8.442366e-17, 
    8.44314e-17, 8.443921e-17, 8.444776e-17, 8.4374e-17, 8.437152e-17, 
    8.437606e-17, 8.438215e-17, 8.438811e-17, 8.439589e-17, 8.439674e-17, 
    8.439817e-17, 8.4402e-17, 8.440517e-17, 8.439852e-17, 8.440597e-17, 
    8.437818e-17, 8.439281e-17, 8.437048e-17, 8.437705e-17, 8.438184e-17, 
    8.437985e-17, 8.439061e-17, 8.439311e-17, 8.440325e-17, 8.439807e-17, 
    8.442939e-17, 8.441549e-17, 8.445464e-17, 8.444359e-17, 8.437062e-17, 
    8.437404e-17, 8.43858e-17, 8.438022e-17, 8.439646e-17, 8.440043e-17, 
    8.440374e-17, 8.440781e-17, 8.440833e-17, 8.441075e-17, 8.440677e-17, 
    8.441064e-17, 8.43959e-17, 8.44025e-17, 8.438458e-17, 8.438887e-17, 
    8.438693e-17, 8.438473e-17, 8.439152e-17, 8.439859e-17, 8.439892e-17, 
    8.440116e-17, 8.440716e-17, 8.439654e-17, 8.443087e-17, 8.440933e-17, 
    8.437776e-17, 8.438412e-17, 8.438523e-17, 8.438273e-17, 8.440002e-17, 
    8.439373e-17, 8.441072e-17, 8.440616e-17, 8.441368e-17, 8.440992e-17, 
    8.440936e-17, 8.440458e-17, 8.440157e-17, 8.439398e-17, 8.438787e-17, 
    8.438312e-17, 8.438423e-17, 8.438946e-17, 8.439906e-17, 8.44083e-17, 
    8.440624e-17, 8.441311e-17, 8.439528e-17, 8.440266e-17, 8.439975e-17, 
    8.440737e-17, 8.439087e-17, 8.440438e-17, 8.438736e-17, 8.438889e-17, 
    8.43936e-17, 8.440303e-17, 8.440539e-17, 8.440758e-17, 8.440626e-17, 
    8.439934e-17, 8.439829e-17, 8.439353e-17, 8.439214e-17, 8.438857e-17, 
    8.438554e-17, 8.438826e-17, 8.439109e-17, 8.439942e-17, 8.440684e-17, 
    8.441501e-17, 8.441708e-17, 8.44262e-17, 8.441853e-17, 8.443095e-17, 
    8.442003e-17, 8.443915e-17, 8.440543e-17, 8.442006e-17, 8.439388e-17, 
    8.439673e-17, 8.440171e-17, 8.441354e-17, 8.440734e-17, 8.441467e-17, 
    8.439826e-17, 8.438956e-17, 8.438752e-17, 8.438337e-17, 8.438762e-17, 
    8.438728e-17, 8.439134e-17, 8.439004e-17, 8.43997e-17, 8.439451e-17, 
    8.44093e-17, 8.441466e-17, 8.443005e-17, 8.443941e-17, 8.444924e-17, 
    8.445349e-17, 8.44548e-17, 8.445534e-17 ;

 MEG_carene_3 =
  3.259629e-17, 3.259968e-17, 3.259904e-17, 3.260175e-17, 3.260027e-17, 
    3.260202e-17, 3.259701e-17, 3.259979e-17, 3.259803e-17, 3.259663e-17, 
    3.260692e-17, 3.260187e-17, 3.261246e-17, 3.260919e-17, 3.261751e-17, 
    3.261191e-17, 3.261865e-17, 3.261742e-17, 3.262131e-17, 3.26202e-17, 
    3.262504e-17, 3.262182e-17, 3.262767e-17, 3.26243e-17, 3.26248e-17, 
    3.26217e-17, 3.260295e-17, 3.260627e-17, 3.260274e-17, 3.260322e-17, 
    3.260302e-17, 3.260028e-17, 3.259885e-17, 3.259607e-17, 3.259659e-17, 
    3.259866e-17, 3.260344e-17, 3.260185e-17, 3.260597e-17, 3.260588e-17, 
    3.261042e-17, 3.260837e-17, 3.261607e-17, 3.261389e-17, 3.262024e-17, 
    3.261863e-17, 3.262016e-17, 3.26197e-17, 3.262016e-17, 3.261781e-17, 
    3.261881e-17, 3.261676e-17, 3.260874e-17, 3.261107e-17, 3.260409e-17, 
    3.25998e-17, 3.259712e-17, 3.259517e-17, 3.259544e-17, 3.259596e-17, 
    3.259867e-17, 3.260128e-17, 3.260325e-17, 3.260456e-17, 3.260586e-17, 
    3.260963e-17, 3.261177e-17, 3.261648e-17, 3.261568e-17, 3.261707e-17, 
    3.261847e-17, 3.262076e-17, 3.262039e-17, 3.262139e-17, 3.261707e-17, 
    3.261992e-17, 3.261522e-17, 3.26165e-17, 3.260599e-17, 3.260229e-17, 
    3.260053e-17, 3.259915e-17, 3.259565e-17, 3.259806e-17, 3.25971e-17, 
    3.259942e-17, 3.260087e-17, 3.260016e-17, 3.26046e-17, 3.260286e-17, 
    3.26119e-17, 3.260801e-17, 3.261831e-17, 3.261585e-17, 3.261891e-17, 
    3.261736e-17, 3.262e-17, 3.261762e-17, 3.262178e-17, 3.262266e-17, 
    3.262205e-17, 3.262446e-17, 3.261749e-17, 3.262013e-17, 3.260013e-17, 
    3.260025e-17, 3.26008e-17, 3.259836e-17, 3.259822e-17, 3.259605e-17, 
    3.2598e-17, 3.259881e-17, 3.260097e-17, 3.26022e-17, 3.260339e-17, 
    3.260601e-17, 3.26089e-17, 3.261301e-17, 3.261601e-17, 3.261801e-17, 
    3.26168e-17, 3.261786e-17, 3.261666e-17, 3.261611e-17, 3.262231e-17, 
    3.261881e-17, 3.262411e-17, 3.262382e-17, 3.26214e-17, 3.262386e-17, 
    3.260033e-17, 3.259967e-17, 3.259731e-17, 3.259915e-17, 3.259582e-17, 
    3.259766e-17, 3.25987e-17, 3.260285e-17, 3.260382e-17, 3.260465e-17, 
    3.260633e-17, 3.260847e-17, 3.261221e-17, 3.261552e-17, 3.261857e-17, 
    3.261835e-17, 3.261842e-17, 3.261908e-17, 3.261742e-17, 3.261936e-17, 
    3.261966e-17, 3.261883e-17, 3.262378e-17, 3.262237e-17, 3.262382e-17, 
    3.26229e-17, 3.259989e-17, 3.260101e-17, 3.26004e-17, 3.260154e-17, 
    3.260072e-17, 3.260429e-17, 3.260536e-17, 3.261045e-17, 3.260842e-17, 
    3.261171e-17, 3.260877e-17, 3.260928e-17, 3.261173e-17, 3.260895e-17, 
    3.261529e-17, 3.26109e-17, 3.261911e-17, 3.261462e-17, 3.261938e-17, 
    3.261855e-17, 3.261995e-17, 3.262118e-17, 3.262277e-17, 3.262563e-17, 
    3.262498e-17, 3.262741e-17, 3.260271e-17, 3.260414e-17, 3.260406e-17, 
    3.260559e-17, 3.260672e-17, 3.260922e-17, 3.261317e-17, 3.26117e-17, 
    3.261446e-17, 3.2615e-17, 3.261083e-17, 3.261335e-17, 3.260514e-17, 
    3.260642e-17, 3.260569e-17, 3.260279e-17, 3.261198e-17, 3.260723e-17, 
    3.261605e-17, 3.261348e-17, 3.2621e-17, 3.261721e-17, 3.262461e-17, 
    3.262767e-17, 3.263075e-17, 3.263413e-17, 3.260497e-17, 3.260399e-17, 
    3.260579e-17, 3.26082e-17, 3.261056e-17, 3.261363e-17, 3.261397e-17, 
    3.261453e-17, 3.261604e-17, 3.26173e-17, 3.261467e-17, 3.261761e-17, 
    3.260663e-17, 3.261241e-17, 3.260358e-17, 3.260618e-17, 3.260808e-17, 
    3.260729e-17, 3.261154e-17, 3.261253e-17, 3.261654e-17, 3.261449e-17, 
    3.262687e-17, 3.262138e-17, 3.263685e-17, 3.263249e-17, 3.260364e-17, 
    3.260499e-17, 3.260964e-17, 3.260743e-17, 3.261386e-17, 3.261542e-17, 
    3.261673e-17, 3.261834e-17, 3.261854e-17, 3.26195e-17, 3.261793e-17, 
    3.261946e-17, 3.261363e-17, 3.261624e-17, 3.260916e-17, 3.261085e-17, 
    3.261009e-17, 3.260922e-17, 3.26119e-17, 3.26147e-17, 3.261482e-17, 
    3.261571e-17, 3.261809e-17, 3.261389e-17, 3.262746e-17, 3.261894e-17, 
    3.260646e-17, 3.260898e-17, 3.260942e-17, 3.260843e-17, 3.261526e-17, 
    3.261277e-17, 3.261949e-17, 3.261769e-17, 3.262066e-17, 3.261918e-17, 
    3.261895e-17, 3.261706e-17, 3.261587e-17, 3.261288e-17, 3.261046e-17, 
    3.260858e-17, 3.260902e-17, 3.261109e-17, 3.261488e-17, 3.261853e-17, 
    3.261772e-17, 3.262044e-17, 3.261339e-17, 3.26163e-17, 3.261515e-17, 
    3.261817e-17, 3.261165e-17, 3.261699e-17, 3.261026e-17, 3.261086e-17, 
    3.261272e-17, 3.261645e-17, 3.261738e-17, 3.261825e-17, 3.261773e-17, 
    3.261499e-17, 3.261458e-17, 3.26127e-17, 3.261214e-17, 3.261074e-17, 
    3.260953e-17, 3.261061e-17, 3.261173e-17, 3.261502e-17, 3.261796e-17, 
    3.262118e-17, 3.2622e-17, 3.262561e-17, 3.262258e-17, 3.262749e-17, 
    3.262317e-17, 3.263073e-17, 3.26174e-17, 3.262318e-17, 3.261283e-17, 
    3.261396e-17, 3.261593e-17, 3.262061e-17, 3.261815e-17, 3.262106e-17, 
    3.261457e-17, 3.261113e-17, 3.261032e-17, 3.260868e-17, 3.261036e-17, 
    3.261023e-17, 3.261183e-17, 3.261132e-17, 3.261513e-17, 3.261308e-17, 
    3.261893e-17, 3.262105e-17, 3.262713e-17, 3.263083e-17, 3.263472e-17, 
    3.26364e-17, 3.263691e-17, 3.263713e-17 ;

 MEG_ethanol =
  1.676205e-18, 1.676468e-18, 1.676418e-18, 1.676627e-18, 1.676513e-18, 
    1.676648e-18, 1.676261e-18, 1.676476e-18, 1.67634e-18, 1.676232e-18, 
    1.677027e-18, 1.676637e-18, 1.677455e-18, 1.677202e-18, 1.677845e-18, 
    1.677412e-18, 1.677933e-18, 1.677838e-18, 1.678138e-18, 1.678052e-18, 
    1.678426e-18, 1.678178e-18, 1.678629e-18, 1.67837e-18, 1.678408e-18, 
    1.678169e-18, 1.67672e-18, 1.676977e-18, 1.676704e-18, 1.676741e-18, 
    1.676726e-18, 1.676514e-18, 1.676403e-18, 1.676189e-18, 1.676229e-18, 
    1.676388e-18, 1.676758e-18, 1.676635e-18, 1.676953e-18, 1.676946e-18, 
    1.677297e-18, 1.677139e-18, 1.677733e-18, 1.677565e-18, 1.678056e-18, 
    1.677932e-18, 1.678049e-18, 1.678014e-18, 1.67805e-18, 1.677868e-18, 
    1.677945e-18, 1.677787e-18, 1.677167e-18, 1.677348e-18, 1.676808e-18, 
    1.676476e-18, 1.676269e-18, 1.676119e-18, 1.67614e-18, 1.676179e-18, 
    1.676389e-18, 1.676591e-18, 1.676743e-18, 1.676845e-18, 1.676945e-18, 
    1.677236e-18, 1.677402e-18, 1.677765e-18, 1.677704e-18, 1.677811e-18, 
    1.677919e-18, 1.678096e-18, 1.678068e-18, 1.678145e-18, 1.677811e-18, 
    1.678031e-18, 1.677668e-18, 1.677767e-18, 1.676955e-18, 1.676669e-18, 
    1.676533e-18, 1.676427e-18, 1.676156e-18, 1.676342e-18, 1.676268e-18, 
    1.676448e-18, 1.676559e-18, 1.676505e-18, 1.676847e-18, 1.676713e-18, 
    1.677412e-18, 1.677111e-18, 1.677907e-18, 1.677717e-18, 1.677953e-18, 
    1.677833e-18, 1.678037e-18, 1.677854e-18, 1.678175e-18, 1.678242e-18, 
    1.678196e-18, 1.678382e-18, 1.677843e-18, 1.678048e-18, 1.676502e-18, 
    1.676511e-18, 1.676554e-18, 1.676365e-18, 1.676355e-18, 1.676187e-18, 
    1.676338e-18, 1.6764e-18, 1.676567e-18, 1.676662e-18, 1.676754e-18, 
    1.676956e-18, 1.67718e-18, 1.677497e-18, 1.677729e-18, 1.677883e-18, 
    1.67779e-18, 1.677872e-18, 1.677779e-18, 1.677737e-18, 1.678216e-18, 
    1.677945e-18, 1.678355e-18, 1.678333e-18, 1.678146e-18, 1.678335e-18, 
    1.676517e-18, 1.676466e-18, 1.676284e-18, 1.676427e-18, 1.676169e-18, 
    1.676311e-18, 1.676391e-18, 1.676712e-18, 1.676787e-18, 1.676851e-18, 
    1.676981e-18, 1.677147e-18, 1.677436e-18, 1.677691e-18, 1.677926e-18, 
    1.67791e-18, 1.677915e-18, 1.677966e-18, 1.677838e-18, 1.677987e-18, 
    1.678011e-18, 1.677947e-18, 1.67833e-18, 1.67822e-18, 1.678332e-18, 
    1.678261e-18, 1.676484e-18, 1.67657e-18, 1.676523e-18, 1.676611e-18, 
    1.676548e-18, 1.676824e-18, 1.676906e-18, 1.677299e-18, 1.677142e-18, 
    1.677397e-18, 1.67717e-18, 1.677209e-18, 1.677398e-18, 1.677183e-18, 
    1.677673e-18, 1.677334e-18, 1.677968e-18, 1.677622e-18, 1.67799e-18, 
    1.677925e-18, 1.678033e-18, 1.678128e-18, 1.678251e-18, 1.678472e-18, 
    1.678422e-18, 1.67861e-18, 1.676701e-18, 1.676812e-18, 1.676806e-18, 
    1.676924e-18, 1.677011e-18, 1.677204e-18, 1.67751e-18, 1.677396e-18, 
    1.677609e-18, 1.677651e-18, 1.677329e-18, 1.677523e-18, 1.676889e-18, 
    1.676988e-18, 1.676931e-18, 1.676708e-18, 1.677418e-18, 1.677051e-18, 
    1.677732e-18, 1.677533e-18, 1.678114e-18, 1.677822e-18, 1.678393e-18, 
    1.678629e-18, 1.678868e-18, 1.679129e-18, 1.676876e-18, 1.676801e-18, 
    1.676939e-18, 1.677125e-18, 1.677308e-18, 1.677545e-18, 1.677571e-18, 
    1.677615e-18, 1.677732e-18, 1.677828e-18, 1.677625e-18, 1.677853e-18, 
    1.677004e-18, 1.677451e-18, 1.676769e-18, 1.67697e-18, 1.677116e-18, 
    1.677055e-18, 1.677384e-18, 1.67746e-18, 1.67777e-18, 1.677612e-18, 
    1.678568e-18, 1.678144e-18, 1.679339e-18, 1.679002e-18, 1.676773e-18, 
    1.676878e-18, 1.677237e-18, 1.677066e-18, 1.677563e-18, 1.677683e-18, 
    1.677785e-18, 1.677909e-18, 1.677925e-18, 1.677999e-18, 1.677877e-18, 
    1.677995e-18, 1.677545e-18, 1.677747e-18, 1.6772e-18, 1.677331e-18, 
    1.677271e-18, 1.677204e-18, 1.677412e-18, 1.677628e-18, 1.677638e-18, 
    1.677706e-18, 1.677889e-18, 1.677565e-18, 1.678613e-18, 1.677956e-18, 
    1.676991e-18, 1.677185e-18, 1.67722e-18, 1.677143e-18, 1.677671e-18, 
    1.677479e-18, 1.677998e-18, 1.677859e-18, 1.678088e-18, 1.677974e-18, 
    1.677956e-18, 1.677811e-18, 1.677718e-18, 1.677487e-18, 1.6773e-18, 
    1.677155e-18, 1.677189e-18, 1.677349e-18, 1.677642e-18, 1.677924e-18, 
    1.677861e-18, 1.678071e-18, 1.677526e-18, 1.677752e-18, 1.677663e-18, 
    1.677896e-18, 1.677392e-18, 1.677805e-18, 1.677285e-18, 1.677331e-18, 
    1.677475e-18, 1.677763e-18, 1.677835e-18, 1.677902e-18, 1.677862e-18, 
    1.67765e-18, 1.677618e-18, 1.677473e-18, 1.67743e-18, 1.677321e-18, 
    1.677229e-18, 1.677312e-18, 1.677399e-18, 1.677653e-18, 1.677879e-18, 
    1.678129e-18, 1.678192e-18, 1.678471e-18, 1.678236e-18, 1.678616e-18, 
    1.678282e-18, 1.678866e-18, 1.677836e-18, 1.678283e-18, 1.677484e-18, 
    1.677571e-18, 1.677723e-18, 1.678084e-18, 1.677895e-18, 1.678119e-18, 
    1.677617e-18, 1.677352e-18, 1.67729e-18, 1.677163e-18, 1.677292e-18, 
    1.677282e-18, 1.677406e-18, 1.677366e-18, 1.677661e-18, 1.677503e-18, 
    1.677955e-18, 1.678118e-18, 1.678588e-18, 1.678874e-18, 1.679174e-18, 
    1.679304e-18, 1.679344e-18, 1.67936e-18 ;

 MEG_formaldehyde =
  3.352411e-19, 3.352936e-19, 3.352836e-19, 3.353254e-19, 3.353026e-19, 
    3.353297e-19, 3.352521e-19, 3.352952e-19, 3.35268e-19, 3.352464e-19, 
    3.354054e-19, 3.353274e-19, 3.354909e-19, 3.354403e-19, 3.35569e-19, 
    3.354825e-19, 3.355866e-19, 3.355675e-19, 3.356276e-19, 3.356104e-19, 
    3.356853e-19, 3.356355e-19, 3.357259e-19, 3.35674e-19, 3.356817e-19, 
    3.356337e-19, 3.353441e-19, 3.353953e-19, 3.353408e-19, 3.353481e-19, 
    3.353451e-19, 3.353027e-19, 3.352807e-19, 3.352377e-19, 3.352457e-19, 
    3.352777e-19, 3.353515e-19, 3.353271e-19, 3.353906e-19, 3.353892e-19, 
    3.354594e-19, 3.354277e-19, 3.355467e-19, 3.35513e-19, 3.356112e-19, 
    3.355863e-19, 3.356098e-19, 3.356028e-19, 3.356099e-19, 3.355735e-19, 
    3.35589e-19, 3.355574e-19, 3.354334e-19, 3.354695e-19, 3.353616e-19, 
    3.352953e-19, 3.352538e-19, 3.352237e-19, 3.35228e-19, 3.352359e-19, 
    3.352778e-19, 3.353182e-19, 3.353487e-19, 3.353689e-19, 3.35389e-19, 
    3.354472e-19, 3.354804e-19, 3.35553e-19, 3.355407e-19, 3.355622e-19, 
    3.355839e-19, 3.356192e-19, 3.356135e-19, 3.356289e-19, 3.355622e-19, 
    3.356062e-19, 3.355335e-19, 3.355533e-19, 3.35391e-19, 3.353338e-19, 
    3.353066e-19, 3.352854e-19, 3.352312e-19, 3.352684e-19, 3.352536e-19, 
    3.352895e-19, 3.353118e-19, 3.353009e-19, 3.353694e-19, 3.353427e-19, 
    3.354823e-19, 3.354221e-19, 3.355813e-19, 3.355433e-19, 3.355906e-19, 
    3.355666e-19, 3.356074e-19, 3.355707e-19, 3.356349e-19, 3.356485e-19, 
    3.356391e-19, 3.356763e-19, 3.355686e-19, 3.356095e-19, 3.353005e-19, 
    3.353022e-19, 3.353108e-19, 3.35273e-19, 3.352709e-19, 3.352374e-19, 
    3.352675e-19, 3.352801e-19, 3.353134e-19, 3.353324e-19, 3.353508e-19, 
    3.353913e-19, 3.354359e-19, 3.354994e-19, 3.355457e-19, 3.355767e-19, 
    3.355579e-19, 3.355744e-19, 3.355558e-19, 3.355473e-19, 3.356432e-19, 
    3.35589e-19, 3.35671e-19, 3.356665e-19, 3.356291e-19, 3.35667e-19, 
    3.353035e-19, 3.352933e-19, 3.352567e-19, 3.352853e-19, 3.352338e-19, 
    3.352622e-19, 3.352783e-19, 3.353425e-19, 3.353574e-19, 3.353702e-19, 
    3.353963e-19, 3.354293e-19, 3.354872e-19, 3.355382e-19, 3.355853e-19, 
    3.355819e-19, 3.355831e-19, 3.355932e-19, 3.355676e-19, 3.355975e-19, 
    3.356022e-19, 3.355894e-19, 3.356659e-19, 3.356441e-19, 3.356664e-19, 
    3.356523e-19, 3.352967e-19, 3.35314e-19, 3.353046e-19, 3.353221e-19, 
    3.353095e-19, 3.353647e-19, 3.353813e-19, 3.354599e-19, 3.354285e-19, 
    3.354794e-19, 3.354339e-19, 3.354418e-19, 3.354796e-19, 3.354366e-19, 
    3.355347e-19, 3.354668e-19, 3.355936e-19, 3.355244e-19, 3.355979e-19, 
    3.355851e-19, 3.356067e-19, 3.356256e-19, 3.356501e-19, 3.356944e-19, 
    3.356843e-19, 3.35722e-19, 3.353402e-19, 3.353624e-19, 3.353611e-19, 
    3.353849e-19, 3.354022e-19, 3.354408e-19, 3.35502e-19, 3.354792e-19, 
    3.355218e-19, 3.355301e-19, 3.354658e-19, 3.355046e-19, 3.353778e-19, 
    3.353976e-19, 3.353863e-19, 3.353416e-19, 3.354835e-19, 3.354102e-19, 
    3.355464e-19, 3.355067e-19, 3.356228e-19, 3.355643e-19, 3.356786e-19, 
    3.357259e-19, 3.357735e-19, 3.358257e-19, 3.353753e-19, 3.353601e-19, 
    3.353878e-19, 3.354251e-19, 3.354615e-19, 3.35509e-19, 3.355142e-19, 
    3.355229e-19, 3.355463e-19, 3.355657e-19, 3.35525e-19, 3.355706e-19, 
    3.354009e-19, 3.354902e-19, 3.353538e-19, 3.353939e-19, 3.354232e-19, 
    3.35411e-19, 3.354767e-19, 3.35492e-19, 3.35554e-19, 3.355223e-19, 
    3.357136e-19, 3.356287e-19, 3.358678e-19, 3.358003e-19, 3.353546e-19, 
    3.353755e-19, 3.354473e-19, 3.354133e-19, 3.355125e-19, 3.355367e-19, 
    3.35557e-19, 3.355818e-19, 3.35585e-19, 3.355998e-19, 3.355754e-19, 
    3.35599e-19, 3.355091e-19, 3.355494e-19, 3.354399e-19, 3.354661e-19, 
    3.354543e-19, 3.354408e-19, 3.354823e-19, 3.355255e-19, 3.355275e-19, 
    3.355412e-19, 3.355779e-19, 3.355129e-19, 3.357227e-19, 3.355911e-19, 
    3.353982e-19, 3.354371e-19, 3.354439e-19, 3.354286e-19, 3.355342e-19, 
    3.354958e-19, 3.355996e-19, 3.355717e-19, 3.356176e-19, 3.355947e-19, 
    3.355913e-19, 3.355621e-19, 3.355437e-19, 3.354973e-19, 3.3546e-19, 
    3.35431e-19, 3.354378e-19, 3.354697e-19, 3.355284e-19, 3.355848e-19, 
    3.355723e-19, 3.356141e-19, 3.355053e-19, 3.355503e-19, 3.355325e-19, 
    3.355791e-19, 3.354783e-19, 3.355609e-19, 3.354569e-19, 3.354662e-19, 
    3.35495e-19, 3.355527e-19, 3.35567e-19, 3.355804e-19, 3.355724e-19, 
    3.355301e-19, 3.355236e-19, 3.354946e-19, 3.354861e-19, 3.354643e-19, 
    3.354458e-19, 3.354624e-19, 3.354797e-19, 3.355305e-19, 3.355759e-19, 
    3.356257e-19, 3.356384e-19, 3.356941e-19, 3.356473e-19, 3.357232e-19, 
    3.356564e-19, 3.357732e-19, 3.355673e-19, 3.356566e-19, 3.354967e-19, 
    3.355141e-19, 3.355446e-19, 3.356168e-19, 3.355789e-19, 3.356237e-19, 
    3.355235e-19, 3.354703e-19, 3.354579e-19, 3.354325e-19, 3.354585e-19, 
    3.354564e-19, 3.354812e-19, 3.354733e-19, 3.355322e-19, 3.355006e-19, 
    3.355909e-19, 3.356236e-19, 3.357176e-19, 3.357748e-19, 3.358347e-19, 
    3.358607e-19, 3.358687e-19, 3.35872e-19 ;

 MEG_isoprene =
  2.29442e-19, 2.294858e-19, 2.294775e-19, 2.295123e-19, 2.294933e-19, 
    2.295159e-19, 2.294512e-19, 2.294872e-19, 2.294645e-19, 2.294465e-19, 
    2.29579e-19, 2.29514e-19, 2.296503e-19, 2.296081e-19, 2.297152e-19, 
    2.296432e-19, 2.2973e-19, 2.29714e-19, 2.297641e-19, 2.297498e-19, 
    2.298121e-19, 2.297707e-19, 2.298459e-19, 2.298027e-19, 2.298091e-19, 
    2.297692e-19, 2.295279e-19, 2.295706e-19, 2.295251e-19, 2.295313e-19, 
    2.295287e-19, 2.294934e-19, 2.29475e-19, 2.294392e-19, 2.294459e-19, 
    2.294725e-19, 2.295341e-19, 2.295137e-19, 2.295667e-19, 2.295655e-19, 
    2.29624e-19, 2.295976e-19, 2.296967e-19, 2.296687e-19, 2.297504e-19, 
    2.297297e-19, 2.297493e-19, 2.297434e-19, 2.297493e-19, 2.29719e-19, 
    2.29732e-19, 2.297056e-19, 2.296024e-19, 2.296324e-19, 2.295424e-19, 
    2.294872e-19, 2.294527e-19, 2.294275e-19, 2.294311e-19, 2.294377e-19, 
    2.294726e-19, 2.295063e-19, 2.295317e-19, 2.295486e-19, 2.295653e-19, 
    2.296138e-19, 2.296414e-19, 2.297019e-19, 2.296917e-19, 2.297096e-19, 
    2.297276e-19, 2.297571e-19, 2.297523e-19, 2.297652e-19, 2.297096e-19, 
    2.297462e-19, 2.296857e-19, 2.297022e-19, 2.29567e-19, 2.295193e-19, 
    2.294966e-19, 2.294789e-19, 2.294338e-19, 2.294648e-19, 2.294525e-19, 
    2.294824e-19, 2.29501e-19, 2.294919e-19, 2.29549e-19, 2.295267e-19, 
    2.296431e-19, 2.295929e-19, 2.297256e-19, 2.296939e-19, 2.297333e-19, 
    2.297133e-19, 2.297473e-19, 2.297167e-19, 2.297701e-19, 2.297815e-19, 
    2.297737e-19, 2.298046e-19, 2.297149e-19, 2.29749e-19, 2.294915e-19, 
    2.29493e-19, 2.295001e-19, 2.294686e-19, 2.294669e-19, 2.294389e-19, 
    2.29464e-19, 2.294745e-19, 2.295023e-19, 2.295182e-19, 2.295335e-19, 
    2.295672e-19, 2.296044e-19, 2.296573e-19, 2.296959e-19, 2.297216e-19, 
    2.29706e-19, 2.297198e-19, 2.297043e-19, 2.296972e-19, 2.29777e-19, 
    2.297319e-19, 2.298002e-19, 2.297965e-19, 2.297653e-19, 2.297969e-19, 
    2.29494e-19, 2.294855e-19, 2.294551e-19, 2.294789e-19, 2.294359e-19, 
    2.294596e-19, 2.29473e-19, 2.295265e-19, 2.29539e-19, 2.295496e-19, 
    2.295714e-19, 2.295989e-19, 2.296471e-19, 2.296896e-19, 2.297288e-19, 
    2.29726e-19, 2.29727e-19, 2.297355e-19, 2.297141e-19, 2.29739e-19, 
    2.297429e-19, 2.297323e-19, 2.29796e-19, 2.297778e-19, 2.297964e-19, 
    2.297846e-19, 2.294884e-19, 2.295028e-19, 2.29495e-19, 2.295096e-19, 
    2.294991e-19, 2.295451e-19, 2.295589e-19, 2.296244e-19, 2.295982e-19, 
    2.296407e-19, 2.296027e-19, 2.296093e-19, 2.296408e-19, 2.29605e-19, 
    2.296867e-19, 2.296302e-19, 2.297358e-19, 2.296781e-19, 2.297393e-19, 
    2.297287e-19, 2.297466e-19, 2.297624e-19, 2.297828e-19, 2.298197e-19, 
    2.298113e-19, 2.298427e-19, 2.295247e-19, 2.295432e-19, 2.295421e-19, 
    2.295619e-19, 2.295764e-19, 2.296085e-19, 2.296595e-19, 2.296405e-19, 
    2.29676e-19, 2.296829e-19, 2.296293e-19, 2.296617e-19, 2.29556e-19, 
    2.295725e-19, 2.29563e-19, 2.295258e-19, 2.296441e-19, 2.29583e-19, 
    2.296964e-19, 2.296634e-19, 2.297601e-19, 2.297114e-19, 2.298065e-19, 
    2.298459e-19, 2.298856e-19, 2.29929e-19, 2.295539e-19, 2.295412e-19, 
    2.295644e-19, 2.295954e-19, 2.296257e-19, 2.296653e-19, 2.296696e-19, 
    2.296769e-19, 2.296964e-19, 2.297125e-19, 2.296787e-19, 2.297166e-19, 
    2.295752e-19, 2.296496e-19, 2.29536e-19, 2.295694e-19, 2.295938e-19, 
    2.295836e-19, 2.296384e-19, 2.296511e-19, 2.297028e-19, 2.296764e-19, 
    2.298357e-19, 2.29765e-19, 2.29964e-19, 2.299078e-19, 2.295367e-19, 
    2.295541e-19, 2.296139e-19, 2.295855e-19, 2.296682e-19, 2.296884e-19, 
    2.297052e-19, 2.297259e-19, 2.297286e-19, 2.297409e-19, 2.297206e-19, 
    2.297403e-19, 2.296654e-19, 2.296989e-19, 2.296077e-19, 2.296296e-19, 
    2.296197e-19, 2.296085e-19, 2.296431e-19, 2.296791e-19, 2.296807e-19, 
    2.296921e-19, 2.297227e-19, 2.296686e-19, 2.298432e-19, 2.297337e-19, 
    2.29573e-19, 2.296054e-19, 2.296111e-19, 2.295983e-19, 2.296863e-19, 
    2.296543e-19, 2.297407e-19, 2.297175e-19, 2.297558e-19, 2.297367e-19, 
    2.297338e-19, 2.297095e-19, 2.296942e-19, 2.296556e-19, 2.296245e-19, 
    2.296003e-19, 2.29606e-19, 2.296326e-19, 2.296815e-19, 2.297284e-19, 
    2.29718e-19, 2.297529e-19, 2.296622e-19, 2.296997e-19, 2.296849e-19, 
    2.297237e-19, 2.296397e-19, 2.297085e-19, 2.296219e-19, 2.296297e-19, 
    2.296537e-19, 2.297017e-19, 2.297136e-19, 2.297248e-19, 2.297181e-19, 
    2.296829e-19, 2.296775e-19, 2.296533e-19, 2.296462e-19, 2.29628e-19, 
    2.296126e-19, 2.296265e-19, 2.296409e-19, 2.296832e-19, 2.29721e-19, 
    2.297625e-19, 2.29773e-19, 2.298195e-19, 2.297805e-19, 2.298437e-19, 
    2.297881e-19, 2.298853e-19, 2.297138e-19, 2.297882e-19, 2.29655e-19, 
    2.296696e-19, 2.296949e-19, 2.297551e-19, 2.297235e-19, 2.297609e-19, 
    2.296773e-19, 2.296331e-19, 2.296227e-19, 2.296016e-19, 2.296232e-19, 
    2.296215e-19, 2.296421e-19, 2.296355e-19, 2.296847e-19, 2.296583e-19, 
    2.297335e-19, 2.297608e-19, 2.29839e-19, 2.298866e-19, 2.299365e-19, 
    2.299581e-19, 2.299648e-19, 2.299675e-19 ;

 MEG_methanol =
  5.79797e-17, 5.798538e-17, 5.79843e-17, 5.798882e-17, 5.798635e-17, 
    5.798929e-17, 5.79809e-17, 5.798556e-17, 5.798261e-17, 5.798028e-17, 
    5.799747e-17, 5.798904e-17, 5.800672e-17, 5.800125e-17, 5.801515e-17, 
    5.80058e-17, 5.801706e-17, 5.801499e-17, 5.802149e-17, 5.801963e-17, 
    5.802771e-17, 5.802234e-17, 5.803209e-17, 5.802649e-17, 5.802732e-17, 
    5.802215e-17, 5.799084e-17, 5.799639e-17, 5.799049e-17, 5.799128e-17, 
    5.799095e-17, 5.798637e-17, 5.798398e-17, 5.797935e-17, 5.798021e-17, 
    5.798366e-17, 5.799165e-17, 5.798901e-17, 5.799588e-17, 5.799572e-17, 
    5.800331e-17, 5.799989e-17, 5.801274e-17, 5.800911e-17, 5.801971e-17, 
    5.801703e-17, 5.801957e-17, 5.801881e-17, 5.801957e-17, 5.801564e-17, 
    5.801732e-17, 5.80139e-17, 5.80005e-17, 5.80044e-17, 5.799273e-17, 
    5.798557e-17, 5.798109e-17, 5.797782e-17, 5.797829e-17, 5.797914e-17, 
    5.798368e-17, 5.798804e-17, 5.799134e-17, 5.799353e-17, 5.79957e-17, 
    5.8002e-17, 5.800558e-17, 5.801342e-17, 5.80121e-17, 5.801441e-17, 
    5.801676e-17, 5.802058e-17, 5.801996e-17, 5.802162e-17, 5.801442e-17, 
    5.801917e-17, 5.801132e-17, 5.801345e-17, 5.799592e-17, 5.798974e-17, 
    5.798678e-17, 5.798449e-17, 5.797863e-17, 5.798266e-17, 5.798106e-17, 
    5.798494e-17, 5.798735e-17, 5.798617e-17, 5.799359e-17, 5.799069e-17, 
    5.800579e-17, 5.799928e-17, 5.801649e-17, 5.801238e-17, 5.801749e-17, 
    5.801489e-17, 5.80193e-17, 5.801534e-17, 5.802227e-17, 5.802374e-17, 
    5.802273e-17, 5.802675e-17, 5.801511e-17, 5.801953e-17, 5.798612e-17, 
    5.798631e-17, 5.798724e-17, 5.798316e-17, 5.798293e-17, 5.79793e-17, 
    5.798256e-17, 5.798392e-17, 5.798752e-17, 5.798958e-17, 5.799157e-17, 
    5.799594e-17, 5.800077e-17, 5.800764e-17, 5.801264e-17, 5.801598e-17, 
    5.801395e-17, 5.801574e-17, 5.801373e-17, 5.801281e-17, 5.802317e-17, 
    5.801731e-17, 5.802616e-17, 5.802569e-17, 5.802165e-17, 5.802574e-17, 
    5.798645e-17, 5.798535e-17, 5.79814e-17, 5.798449e-17, 5.797891e-17, 
    5.798199e-17, 5.798373e-17, 5.799067e-17, 5.799228e-17, 5.799367e-17, 
    5.799648e-17, 5.800006e-17, 5.800631e-17, 5.801182e-17, 5.801691e-17, 
    5.801655e-17, 5.801667e-17, 5.801777e-17, 5.801499e-17, 5.801823e-17, 
    5.801874e-17, 5.801736e-17, 5.802562e-17, 5.802327e-17, 5.802568e-17, 
    5.802415e-17, 5.798572e-17, 5.798759e-17, 5.798657e-17, 5.798847e-17, 
    5.798711e-17, 5.799308e-17, 5.799486e-17, 5.800336e-17, 5.799997e-17, 
    5.800548e-17, 5.800055e-17, 5.800141e-17, 5.80055e-17, 5.800085e-17, 
    5.801145e-17, 5.800411e-17, 5.801781e-17, 5.801033e-17, 5.801828e-17, 
    5.801689e-17, 5.801922e-17, 5.802127e-17, 5.802392e-17, 5.802871e-17, 
    5.802761e-17, 5.803168e-17, 5.799042e-17, 5.799283e-17, 5.799269e-17, 
    5.799525e-17, 5.799713e-17, 5.80013e-17, 5.800791e-17, 5.800544e-17, 
    5.801005e-17, 5.801095e-17, 5.8004e-17, 5.80082e-17, 5.799449e-17, 
    5.799662e-17, 5.799541e-17, 5.799058e-17, 5.800591e-17, 5.799799e-17, 
    5.801271e-17, 5.800842e-17, 5.802097e-17, 5.801465e-17, 5.802699e-17, 
    5.80321e-17, 5.803724e-17, 5.804288e-17, 5.799422e-17, 5.799257e-17, 
    5.799558e-17, 5.79996e-17, 5.800354e-17, 5.800867e-17, 5.800923e-17, 
    5.801018e-17, 5.80127e-17, 5.80148e-17, 5.80104e-17, 5.801532e-17, 
    5.799698e-17, 5.800664e-17, 5.799189e-17, 5.799623e-17, 5.799939e-17, 
    5.799808e-17, 5.800519e-17, 5.800683e-17, 5.801353e-17, 5.801011e-17, 
    5.803078e-17, 5.80216e-17, 5.804742e-17, 5.804013e-17, 5.799199e-17, 
    5.799424e-17, 5.8002e-17, 5.799832e-17, 5.800905e-17, 5.801167e-17, 
    5.801385e-17, 5.801654e-17, 5.801687e-17, 5.801847e-17, 5.801585e-17, 
    5.80184e-17, 5.800868e-17, 5.801303e-17, 5.80012e-17, 5.800404e-17, 
    5.800276e-17, 5.80013e-17, 5.800579e-17, 5.801045e-17, 5.801067e-17, 
    5.801215e-17, 5.801611e-17, 5.80091e-17, 5.803175e-17, 5.801754e-17, 
    5.79967e-17, 5.80009e-17, 5.800163e-17, 5.799999e-17, 5.801139e-17, 
    5.800724e-17, 5.801845e-17, 5.801544e-17, 5.802041e-17, 5.801793e-17, 
    5.801756e-17, 5.801441e-17, 5.801242e-17, 5.800741e-17, 5.800337e-17, 
    5.800024e-17, 5.800098e-17, 5.800443e-17, 5.801077e-17, 5.801685e-17, 
    5.80155e-17, 5.802003e-17, 5.800826e-17, 5.801313e-17, 5.801122e-17, 
    5.801624e-17, 5.800536e-17, 5.801428e-17, 5.800304e-17, 5.800405e-17, 
    5.800716e-17, 5.801339e-17, 5.801494e-17, 5.801638e-17, 5.801552e-17, 
    5.801095e-17, 5.801025e-17, 5.800711e-17, 5.800619e-17, 5.800384e-17, 
    5.800183e-17, 5.800363e-17, 5.80055e-17, 5.8011e-17, 5.801589e-17, 
    5.802128e-17, 5.802265e-17, 5.802867e-17, 5.802361e-17, 5.80318e-17, 
    5.80246e-17, 5.803721e-17, 5.801497e-17, 5.802462e-17, 5.800734e-17, 
    5.800922e-17, 5.801251e-17, 5.802031e-17, 5.801622e-17, 5.802107e-17, 
    5.801024e-17, 5.800449e-17, 5.800315e-17, 5.800041e-17, 5.800321e-17, 
    5.800298e-17, 5.800566e-17, 5.800481e-17, 5.801118e-17, 5.800776e-17, 
    5.801752e-17, 5.802106e-17, 5.803121e-17, 5.803738e-17, 5.804385e-17, 
    5.804666e-17, 5.804752e-17, 5.804788e-17 ;

 MEG_pinene_a =
  4.795989e-17, 4.796509e-17, 4.79641e-17, 4.796825e-17, 4.796599e-17, 
    4.796868e-17, 4.796099e-17, 4.796526e-17, 4.796256e-17, 4.796042e-17, 
    4.797618e-17, 4.796845e-17, 4.798467e-17, 4.797965e-17, 4.79924e-17, 
    4.798382e-17, 4.799415e-17, 4.799226e-17, 4.799822e-17, 4.799652e-17, 
    4.800394e-17, 4.799901e-17, 4.800796e-17, 4.800282e-17, 4.800358e-17, 
    4.799883e-17, 4.79701e-17, 4.797519e-17, 4.796978e-17, 4.797051e-17, 
    4.797021e-17, 4.7966e-17, 4.796382e-17, 4.795956e-17, 4.796035e-17, 
    4.796352e-17, 4.797084e-17, 4.796842e-17, 4.797472e-17, 4.797458e-17, 
    4.798154e-17, 4.79784e-17, 4.799019e-17, 4.798686e-17, 4.799659e-17, 
    4.799412e-17, 4.799646e-17, 4.799576e-17, 4.799647e-17, 4.799286e-17, 
    4.79944e-17, 4.799126e-17, 4.797897e-17, 4.798254e-17, 4.797184e-17, 
    4.796526e-17, 4.796116e-17, 4.795817e-17, 4.795859e-17, 4.795938e-17, 
    4.796354e-17, 4.796754e-17, 4.797056e-17, 4.797256e-17, 4.797456e-17, 
    4.798033e-17, 4.798362e-17, 4.799082e-17, 4.79896e-17, 4.799173e-17, 
    4.799388e-17, 4.799739e-17, 4.799682e-17, 4.799835e-17, 4.799174e-17, 
    4.79961e-17, 4.798889e-17, 4.799085e-17, 4.797475e-17, 4.796909e-17, 
    4.796638e-17, 4.796428e-17, 4.795891e-17, 4.79626e-17, 4.796114e-17, 
    4.796469e-17, 4.79669e-17, 4.796582e-17, 4.797262e-17, 4.796996e-17, 
    4.798381e-17, 4.797784e-17, 4.799363e-17, 4.798986e-17, 4.799455e-17, 
    4.799217e-17, 4.799622e-17, 4.799258e-17, 4.799894e-17, 4.800029e-17, 
    4.799936e-17, 4.800305e-17, 4.799237e-17, 4.799642e-17, 4.796578e-17, 
    4.796595e-17, 4.79668e-17, 4.796306e-17, 4.796285e-17, 4.795952e-17, 
    4.796251e-17, 4.796376e-17, 4.796706e-17, 4.796895e-17, 4.797077e-17, 
    4.797478e-17, 4.797921e-17, 4.798551e-17, 4.79901e-17, 4.799316e-17, 
    4.799131e-17, 4.799295e-17, 4.79911e-17, 4.799026e-17, 4.799976e-17, 
    4.799439e-17, 4.800252e-17, 4.800208e-17, 4.799837e-17, 4.800213e-17, 
    4.796608e-17, 4.796507e-17, 4.796144e-17, 4.796428e-17, 4.795916e-17, 
    4.796198e-17, 4.796358e-17, 4.796994e-17, 4.797143e-17, 4.797269e-17, 
    4.797528e-17, 4.797856e-17, 4.798429e-17, 4.798935e-17, 4.799402e-17, 
    4.799369e-17, 4.79938e-17, 4.799481e-17, 4.799226e-17, 4.799523e-17, 
    4.79957e-17, 4.799443e-17, 4.800202e-17, 4.799985e-17, 4.800207e-17, 
    4.800067e-17, 4.79654e-17, 4.796713e-17, 4.796619e-17, 4.796793e-17, 
    4.796668e-17, 4.797215e-17, 4.797379e-17, 4.798159e-17, 4.797847e-17, 
    4.798353e-17, 4.797901e-17, 4.797979e-17, 4.798354e-17, 4.797928e-17, 
    4.7989e-17, 4.798228e-17, 4.799485e-17, 4.798798e-17, 4.799528e-17, 
    4.7994e-17, 4.799614e-17, 4.799803e-17, 4.800046e-17, 4.800485e-17, 
    4.800385e-17, 4.800758e-17, 4.796972e-17, 4.797192e-17, 4.797179e-17, 
    4.797415e-17, 4.797587e-17, 4.797969e-17, 4.798576e-17, 4.79835e-17, 
    4.798773e-17, 4.798855e-17, 4.798217e-17, 4.798602e-17, 4.797345e-17, 
    4.797541e-17, 4.797429e-17, 4.796986e-17, 4.798393e-17, 4.797666e-17, 
    4.799016e-17, 4.798623e-17, 4.799775e-17, 4.799194e-17, 4.800328e-17, 
    4.800796e-17, 4.801269e-17, 4.801787e-17, 4.79732e-17, 4.797169e-17, 
    4.797444e-17, 4.797813e-17, 4.798175e-17, 4.798646e-17, 4.798697e-17, 
    4.798784e-17, 4.799016e-17, 4.799208e-17, 4.798805e-17, 4.799257e-17, 
    4.797573e-17, 4.79846e-17, 4.797107e-17, 4.797505e-17, 4.797795e-17, 
    4.797674e-17, 4.798326e-17, 4.798477e-17, 4.799092e-17, 4.798778e-17, 
    4.800675e-17, 4.799833e-17, 4.802204e-17, 4.801535e-17, 4.797115e-17, 
    4.797322e-17, 4.798034e-17, 4.797697e-17, 4.798681e-17, 4.79892e-17, 
    4.799121e-17, 4.799367e-17, 4.799399e-17, 4.799546e-17, 4.799305e-17, 
    4.799539e-17, 4.798647e-17, 4.799046e-17, 4.797961e-17, 4.798221e-17, 
    4.798103e-17, 4.79797e-17, 4.798381e-17, 4.79881e-17, 4.798829e-17, 
    4.798965e-17, 4.799329e-17, 4.798685e-17, 4.800764e-17, 4.79946e-17, 
    4.797548e-17, 4.797932e-17, 4.798e-17, 4.797849e-17, 4.798896e-17, 
    4.798515e-17, 4.799544e-17, 4.799268e-17, 4.799723e-17, 4.799496e-17, 
    4.799462e-17, 4.799173e-17, 4.79899e-17, 4.79853e-17, 4.79816e-17, 
    4.797872e-17, 4.79794e-17, 4.798256e-17, 4.798838e-17, 4.799397e-17, 
    4.799273e-17, 4.799689e-17, 4.798609e-17, 4.799055e-17, 4.798879e-17, 
    4.799341e-17, 4.798342e-17, 4.79916e-17, 4.798129e-17, 4.798222e-17, 
    4.798507e-17, 4.799079e-17, 4.799221e-17, 4.799354e-17, 4.799274e-17, 
    4.798855e-17, 4.798791e-17, 4.798503e-17, 4.798418e-17, 4.798202e-17, 
    4.798019e-17, 4.798184e-17, 4.798355e-17, 4.79886e-17, 4.799309e-17, 
    4.799804e-17, 4.799929e-17, 4.800482e-17, 4.800017e-17, 4.800769e-17, 
    4.800108e-17, 4.801266e-17, 4.799223e-17, 4.80011e-17, 4.798524e-17, 
    4.798697e-17, 4.798999e-17, 4.799715e-17, 4.799339e-17, 4.799784e-17, 
    4.798789e-17, 4.798262e-17, 4.798139e-17, 4.797888e-17, 4.798145e-17, 
    4.798124e-17, 4.79837e-17, 4.798291e-17, 4.798876e-17, 4.798562e-17, 
    4.799458e-17, 4.799783e-17, 4.800715e-17, 4.801281e-17, 4.801876e-17, 
    4.802134e-17, 4.802213e-17, 4.802246e-17 ;

 MEG_thujene_a =
  1.210137e-18, 1.210263e-18, 1.210239e-18, 1.21034e-18, 1.210285e-18, 
    1.21035e-18, 1.210164e-18, 1.210267e-18, 1.210202e-18, 1.21015e-18, 
    1.210532e-18, 1.210345e-18, 1.210738e-18, 1.210616e-18, 1.210925e-18, 
    1.210717e-18, 1.210967e-18, 1.210921e-18, 1.211066e-18, 1.211025e-18, 
    1.211205e-18, 1.211085e-18, 1.211302e-18, 1.211177e-18, 1.211196e-18, 
    1.211081e-18, 1.210385e-18, 1.210508e-18, 1.210377e-18, 1.210395e-18, 
    1.210387e-18, 1.210285e-18, 1.210232e-18, 1.210129e-18, 1.210148e-18, 
    1.210225e-18, 1.210403e-18, 1.210344e-18, 1.210497e-18, 1.210493e-18, 
    1.210662e-18, 1.210586e-18, 1.210871e-18, 1.210791e-18, 1.211027e-18, 
    1.210967e-18, 1.211023e-18, 1.211006e-18, 1.211023e-18, 1.210936e-18, 
    1.210973e-18, 1.210897e-18, 1.210599e-18, 1.210686e-18, 1.210427e-18, 
    1.210267e-18, 1.210168e-18, 1.210096e-18, 1.210106e-18, 1.210125e-18, 
    1.210226e-18, 1.210323e-18, 1.210396e-18, 1.210444e-18, 1.210493e-18, 
    1.210633e-18, 1.210712e-18, 1.210887e-18, 1.210857e-18, 1.210909e-18, 
    1.210961e-18, 1.211046e-18, 1.211032e-18, 1.211069e-18, 1.210909e-18, 
    1.211015e-18, 1.21084e-18, 1.210887e-18, 1.210497e-18, 1.21036e-18, 
    1.210295e-18, 1.210244e-18, 1.210114e-18, 1.210203e-18, 1.210167e-18, 
    1.210254e-18, 1.210307e-18, 1.210281e-18, 1.210446e-18, 1.210381e-18, 
    1.210717e-18, 1.210572e-18, 1.210955e-18, 1.210863e-18, 1.210977e-18, 
    1.210919e-18, 1.211017e-18, 1.210929e-18, 1.211084e-18, 1.211116e-18, 
    1.211094e-18, 1.211183e-18, 1.210924e-18, 1.211022e-18, 1.21028e-18, 
    1.210284e-18, 1.210305e-18, 1.210214e-18, 1.210209e-18, 1.210128e-18, 
    1.210201e-18, 1.210231e-18, 1.210311e-18, 1.210357e-18, 1.210401e-18, 
    1.210498e-18, 1.210605e-18, 1.210758e-18, 1.210869e-18, 1.210944e-18, 
    1.210899e-18, 1.210938e-18, 1.210894e-18, 1.210873e-18, 1.211103e-18, 
    1.210973e-18, 1.21117e-18, 1.21116e-18, 1.21107e-18, 1.211161e-18, 
    1.210287e-18, 1.210263e-18, 1.210175e-18, 1.210244e-18, 1.21012e-18, 
    1.210188e-18, 1.210227e-18, 1.210381e-18, 1.210417e-18, 1.210448e-18, 
    1.21051e-18, 1.210589e-18, 1.210729e-18, 1.210851e-18, 1.210964e-18, 
    1.210956e-18, 1.210959e-18, 1.210983e-18, 1.210922e-18, 1.210994e-18, 
    1.211005e-18, 1.210974e-18, 1.211158e-18, 1.211106e-18, 1.211159e-18, 
    1.211125e-18, 1.210271e-18, 1.210313e-18, 1.21029e-18, 1.210332e-18, 
    1.210302e-18, 1.210434e-18, 1.210474e-18, 1.210663e-18, 1.210588e-18, 
    1.21071e-18, 1.210601e-18, 1.210619e-18, 1.21071e-18, 1.210607e-18, 
    1.210843e-18, 1.21068e-18, 1.210984e-18, 1.210818e-18, 1.210995e-18, 
    1.210964e-18, 1.211016e-18, 1.211061e-18, 1.21112e-18, 1.211227e-18, 
    1.211202e-18, 1.211293e-18, 1.210375e-18, 1.210429e-18, 1.210426e-18, 
    1.210483e-18, 1.210524e-18, 1.210617e-18, 1.210764e-18, 1.210709e-18, 
    1.210812e-18, 1.210832e-18, 1.210677e-18, 1.210771e-18, 1.210466e-18, 
    1.210513e-18, 1.210486e-18, 1.210379e-18, 1.21072e-18, 1.210544e-18, 
    1.210871e-18, 1.210775e-18, 1.211055e-18, 1.210914e-18, 1.211189e-18, 
    1.211302e-18, 1.211417e-18, 1.211542e-18, 1.21046e-18, 1.210423e-18, 
    1.21049e-18, 1.210579e-18, 1.210667e-18, 1.210781e-18, 1.210793e-18, 
    1.210814e-18, 1.210871e-18, 1.210917e-18, 1.21082e-18, 1.210929e-18, 
    1.210521e-18, 1.210736e-18, 1.210408e-18, 1.210504e-18, 1.210575e-18, 
    1.210546e-18, 1.210703e-18, 1.21074e-18, 1.210889e-18, 1.210813e-18, 
    1.211273e-18, 1.211069e-18, 1.211643e-18, 1.211481e-18, 1.21041e-18, 
    1.21046e-18, 1.210633e-18, 1.210551e-18, 1.210789e-18, 1.210848e-18, 
    1.210896e-18, 1.210956e-18, 1.210963e-18, 1.210999e-18, 1.210941e-18, 
    1.210997e-18, 1.210781e-18, 1.210878e-18, 1.210615e-18, 1.210678e-18, 
    1.21065e-18, 1.210617e-18, 1.210717e-18, 1.210821e-18, 1.210825e-18, 
    1.210858e-18, 1.210946e-18, 1.21079e-18, 1.211294e-18, 1.210978e-18, 
    1.210515e-18, 1.210608e-18, 1.210625e-18, 1.210588e-18, 1.210842e-18, 
    1.210749e-18, 1.210999e-18, 1.210932e-18, 1.211042e-18, 1.210987e-18, 
    1.210979e-18, 1.210909e-18, 1.210864e-18, 1.210753e-18, 1.210663e-18, 
    1.210594e-18, 1.21061e-18, 1.210687e-18, 1.210828e-18, 1.210963e-18, 
    1.210933e-18, 1.211034e-18, 1.210772e-18, 1.21088e-18, 1.210838e-18, 
    1.210949e-18, 1.210707e-18, 1.210906e-18, 1.210656e-18, 1.210678e-18, 
    1.210747e-18, 1.210886e-18, 1.21092e-18, 1.210953e-18, 1.210933e-18, 
    1.210832e-18, 1.210816e-18, 1.210746e-18, 1.210726e-18, 1.210674e-18, 
    1.210629e-18, 1.210669e-18, 1.210711e-18, 1.210833e-18, 1.210942e-18, 
    1.211061e-18, 1.211092e-18, 1.211226e-18, 1.211113e-18, 1.211296e-18, 
    1.211135e-18, 1.211416e-18, 1.210921e-18, 1.211136e-18, 1.210751e-18, 
    1.210793e-18, 1.210866e-18, 1.21104e-18, 1.210949e-18, 1.211057e-18, 
    1.210816e-18, 1.210688e-18, 1.210658e-18, 1.210597e-18, 1.21066e-18, 
    1.210655e-18, 1.210714e-18, 1.210695e-18, 1.210837e-18, 1.210761e-18, 
    1.210978e-18, 1.211056e-18, 1.211282e-18, 1.21142e-18, 1.211564e-18, 
    1.211626e-18, 1.211645e-18, 1.211653e-18 ;

 MR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 M_LITR1C_TO_LEACHING =
  -8.240992e-27, 2.334972e-25, 1.922918e-25, -3.021727e-25, -4.669934e-26, 
    -2.060268e-25, 1.950388e-25, -2.637143e-25, -3.735953e-25, -9.065174e-26, 
    1.483394e-25, -3.076667e-25, -8.241066e-26, -3.763423e-25, 2.362442e-25, 
    -3.323899e-25, -2.170149e-25, -1.895446e-25, -3.681012e-25, 
    -4.944636e-26, -1.20869e-25, -3.186548e-25, -1.758095e-25, -4.065596e-25, 
    4.505122e-25, 1.895448e-25, -7.691661e-26, -7.966364e-26, -3.598602e-25, 
    3.296438e-26, 1.813037e-25, -2.774494e-25, -1.071339e-25, 6.043463e-26, 
    -7.691661e-26, -6.455508e-25, -6.318148e-26, -2.884375e-25, 
    -2.087738e-25, -1.318571e-25, -5.246816e-25, -1.648207e-26, 1.703156e-25, 
    3.598603e-25, -1.538333e-25, 3.516192e-25, -2.197619e-25, -3.763423e-25, 
    -2.087738e-25, 2.362442e-25, -6.675269e-25, 2.801966e-25, -5.768744e-26, 
    -1.758095e-25, 1.428454e-25, -1.23616e-25, -2.417381e-25, 1.620745e-25, 
    -2.829435e-25, -8.241066e-26, 1.922918e-25, -9.065174e-26, 4.889705e-25, 
    8.241083e-26, -9.339876e-26, 2.747026e-25, 7.142273e-26, 1.318573e-25, 
    9.614595e-26, -1.098802e-26, -3.37884e-25, -4.120529e-26, -2.801964e-25, 
    -1.648214e-25, 8.241157e-27, -2.582203e-25, -2.939316e-25, -2.3075e-25, 
    -2.142679e-25, 1.538335e-25, -1.730625e-25, 2.499793e-25, 1.483394e-25, 
    8.241157e-27, 1.730626e-25, -1.813036e-25, 1.840507e-25, 2.334972e-25, 
    -1.648207e-26, 3.049198e-25, -6.592851e-26, -3.571124e-26, 4.66995e-26, 
    -4.56006e-25, -4.889703e-25, -4.120529e-26, -2.142679e-25, 3.57114e-26, 
    1.153751e-25, 1.0164e-25, 6.592867e-26, 2.334972e-25, 5.494132e-27, 
    2.774496e-25, 8.241157e-27, 7.691677e-26, -4.944636e-26, -1.016398e-25, 
    -8.543246e-25, -5.164406e-25, 2.08774e-25, -1.510863e-25, -1.15375e-25, 
    -3.104137e-25, -2.884375e-25, -4.807293e-25, -1.758095e-25, 4.697413e-25, 
    2.856907e-25, 3.653544e-25, -4.50512e-25, -5.494041e-26, -4.779822e-25, 
    7.691677e-26, -3.516191e-25, -2.197619e-25, -2.197612e-26, 1.758097e-25, 
    1.373521e-26, 2.472323e-25, -6.867554e-26, -1.318571e-25, -2.774494e-25, 
    -3.873304e-25, -2.609673e-25, -4.120536e-25, 6.592867e-26, -3.351369e-25, 
    4.972116e-25, -1.23616e-25, 4.230419e-25, 2.747107e-27, -5.493967e-27, 
    -1.318571e-25, -1.23616e-25, 5.658872e-25, -4.120536e-25, -2.774494e-25, 
    2.280031e-25, 2.554734e-25, -2.197619e-25, -1.620744e-25, 6.757682e-25, 
    6.53792e-25, 6.043463e-26, -3.351369e-25, -1.400982e-25, -1.098809e-25, 
    -2.417381e-25, 1.318573e-25, 1.098811e-25, 2.11521e-25, -5.494041e-26, 
    -4.752352e-25, 7.142273e-26, 4.834764e-25, 1.867978e-25, 3.543663e-25, 
    4.120538e-25, -4.58753e-25, 1.620745e-25, -1.373512e-25, 3.296438e-26, 
    -4.669934e-26, 1.840507e-25, -9.614578e-26, 8.241157e-27, -4.038125e-25, 
    -2.554732e-25, -4.312828e-25, 1.428454e-25, -1.867976e-25, 7.416975e-26, 
    1.291103e-25, -2.994256e-25, -2.664613e-25, -4.669934e-26, -4.120529e-26, 
    1.785567e-25, -1.318571e-25, 2.280031e-25, 1.263632e-25, 1.263632e-25, 
    -8.515768e-26, -2.36244e-25, -3.323899e-25, 3.461252e-25, 8.25776e-32, 
    1.620745e-25, 4.395248e-26, 1.098811e-25, -3.571131e-25, 1.318573e-25, 
    -2.032798e-25, -7.142256e-26, 6.86757e-26, -9.614578e-26, -1.510863e-25, 
    -5.494041e-26, 1.977859e-25, -1.620744e-25, -1.950387e-25, -1.428452e-25, 
    -4.230417e-25, -2.911845e-25, 6.318165e-26, 3.735955e-25, 1.785567e-25, 
    1.922926e-26, 3.021735e-26, 2.747107e-27, 5.76876e-26, -1.922916e-25, 
    -7.691661e-26, -2.939316e-25, -1.538333e-25, -7.004912e-25, 2.08774e-25, 
    -4.175477e-25, 4.257889e-25, 8.515785e-26, 2.527264e-25, 1.730626e-25, 
    2.060269e-25, -4.148007e-25, -2.472321e-25, 6.86757e-26, 1.373521e-26, 
    -2.966786e-25, -1.23616e-25, -4.422709e-25, -9.065174e-26, 1.181221e-25, 
    -3.214018e-25, 3.488722e-25, 2.334972e-25, -2.472321e-25, 8.241157e-27, 
    -1.098809e-25, -1.648207e-26, 2.747033e-26, -3.296429e-25, 9.889298e-26, 
    1.620745e-25, -4.285358e-25, 2.334972e-25, 2.362442e-25, 4.944653e-26, 
    -7.691661e-26, -2.225089e-25, 5.603931e-25, 1.813037e-25, 1.593275e-25, 
    2.362442e-25, -2.527262e-25, -1.23616e-25, -6.510448e-25, -2.994256e-25, 
    -2.417381e-25, 1.620745e-25, -3.104137e-25, 2.719555e-25, 1.181221e-25, 
    -2.25256e-25, 2.334972e-25, -2.774494e-25, -4.53259e-25, -3.241488e-25, 
    8.241083e-26, -1.263631e-25, -2.774494e-25, 7.142273e-26, 6.620331e-25, 
    -2.25256e-25, -1.400982e-25, 1.400983e-25, -1.098809e-25, -3.43378e-25, 
    6.180807e-25, -7.966364e-26, 5.109467e-25, -1.346041e-25, -2.499792e-25, 
    -9.889281e-26, 4.065598e-25, -2.994256e-25, 1.373521e-26, -8.240992e-27, 
    7.416975e-26, -3.214018e-25, -6.455508e-25, -2.939316e-25, -3.021727e-25, 
    -2.746942e-27, 3.653544e-25, 5.548991e-25, -2.747024e-25, -2.197619e-25, 
    -9.889281e-26, -1.950387e-25, 1.620745e-25, 9.06519e-26, -2.36244e-25, 
    -1.840506e-25, -3.131607e-25, 8.790487e-26, -3.40631e-25, 5.76876e-26, 
    -1.648214e-25, 8.515785e-26, 3.021735e-26, 1.373513e-25, -5.576459e-25, 
    -2.472321e-25, -3.214018e-25, 1.373513e-25, 3.433782e-25, 4.889705e-25, 
    -3.818364e-25, 8.790487e-26, -2.747016e-26, 1.04387e-25, 2.472323e-25, 
    -2.472321e-25, 2.005329e-25, 4.450181e-25, -2.554732e-25, 8.257433e-32 ;

 M_LITR2C_TO_LEACHING =
  -5.494044e-26, -3.296424e-26, 7.14227e-26, -2.74702e-26, -1.703155e-25, 
    -1.730625e-25, -2.032798e-25, 1.593275e-25, -4.669937e-26, -6.592854e-26, 
    6.867567e-26, 4.669947e-26, -2.197614e-26, 4.395245e-26, 1.428453e-25, 
    -1.071339e-25, -2.527262e-25, 4.395245e-26, 3.021733e-26, -1.785566e-25, 
    -6.592854e-26, 1.346043e-25, 2.19762e-25, -5.768747e-26, -7.142259e-26, 
    1.098815e-26, 8.241128e-27, -2.966786e-25, -3.021722e-26, -3.845829e-26, 
    -7.416961e-26, 6.318163e-26, -1.318571e-25, -1.400982e-25, -5.219342e-26, 
    -2.142679e-25, 8.790485e-26, -1.510863e-25, 3.021733e-26, -1.758095e-25, 
    -1.648209e-26, 5.494103e-27, -1.813036e-25, -1.15375e-25, -9.339879e-26, 
    -1.895447e-25, 3.24149e-25, -8.515771e-26, 2.774496e-25, -1.922912e-26, 
    9.339889e-26, -9.889284e-26, 5.494103e-27, -3.268959e-25, 2.307501e-25, 
    -7.142259e-26, 9.339889e-26, 1.208691e-25, -7.142259e-26, -2.74702e-26, 
    7.691675e-26, -1.400982e-25, -5.768747e-26, -2.472317e-26, -4.038126e-25, 
    -5.219342e-26, -3.021722e-26, -1.15375e-25, -1.867976e-25, -1.043869e-25, 
    -8.241021e-27, 1.922918e-25, -1.373507e-26, 3.021733e-26, -2.25256e-25, 
    -1.565804e-25, 1.04387e-25, -2.637143e-25, 1.510864e-25, -5.494044e-26, 
    -2.746971e-27, 5.351492e-32, -1.236161e-25, 2.939317e-25, -4.944639e-26, 
    -4.669937e-26, 9.065187e-26, 6.867567e-26, -8.241069e-26, 9.889295e-26, 
    -5.219342e-26, 4.120543e-26, 8.790485e-26, 9.614592e-26, -1.648209e-26, 
    1.840507e-25, -6.592854e-26, 4.120543e-26, -6.867557e-26, -1.428452e-25, 
    1.813037e-25, -1.867976e-25, 2.14268e-25, 1.483394e-25, 1.620745e-25, 
    1.758096e-25, -1.043869e-25, 3.296435e-26, -7.142259e-26, 3.84584e-26, 
    -1.20869e-25, 3.433782e-25, -1.758095e-25, -1.593274e-25, -2.142679e-25, 
    -1.12628e-25, -7.691664e-26, -1.565804e-25, -9.889284e-26, 1.483394e-25, 
    1.593275e-25, -2.197614e-26, -3.653542e-25, 2.609674e-25, -1.18122e-25, 
    -1.785566e-25, -1.977857e-25, -1.648209e-26, 7.14227e-26, 9.614592e-26, 
    -2.774495e-25, 1.153751e-25, -1.428452e-25, -4.340298e-25, -2.966786e-25, 
    -6.867557e-26, -6.043449e-26, -9.339879e-26, 4.230418e-25, -4.395234e-26, 
    -2.746971e-27, 1.64822e-26, 1.373518e-26, -1.098809e-25, 1.181221e-25, 
    -1.346042e-25, 8.24108e-26, -2.197619e-25, -1.593274e-25, -1.291101e-25, 
    -2.746971e-27, -7.142259e-26, -1.648209e-26, 6.592865e-26, -3.159078e-25, 
    -2.087738e-25, -8.515771e-26, -2.746971e-27, 4.395245e-26, 1.263632e-25, 
    2.747078e-27, 1.291102e-25, -1.730625e-25, -1.455923e-25, -2.472317e-26, 
    2.499793e-25, -2.829435e-25, -1.098805e-26, -2.032798e-25, 2.14268e-25, 
    -4.615001e-25, -2.25256e-25, -3.296424e-26, -2.472317e-26, 7.691675e-26, 
    -1.20869e-25, 1.675686e-25, 1.098815e-26, 2.060269e-25, -1.593274e-25, 
    -2.115208e-25, 2.19762e-25, 2.14268e-25, -1.510863e-25, -4.120532e-26, 
    1.236162e-25, -2.225089e-25, -2.417381e-25, -1.648209e-26, 5.494055e-26, 
    1.09881e-25, -7.691664e-26, -2.087738e-25, -5.219342e-26, 1.373513e-25, 
    -1.373507e-26, -1.593274e-25, 5.494103e-27, -2.74702e-26, 2.252561e-25, 
    -5.493996e-27, 1.785567e-25, 2.747078e-27, -1.813036e-25, 1.483394e-25, 
    -1.922912e-26, 1.922923e-26, -3.681013e-25, -2.994256e-25, -7.691664e-26, 
    -6.318152e-26, -8.790474e-26, 2.005329e-25, 1.483394e-25, -3.296424e-26, 
    -7.691664e-26, -8.241021e-27, -9.889284e-26, -2.417381e-25, 
    -1.758095e-25, -9.889284e-26, -1.565804e-25, -2.939316e-25, 1.263632e-25, 
    -1.236161e-25, -5.219342e-26, 1.758096e-25, -7.691664e-26, 6.867567e-26, 
    1.09881e-25, -1.703155e-25, 5.351456e-32, 2.417382e-25, -2.417381e-25, 
    -2.472322e-25, -1.867976e-25, -9.339879e-26, -4.944639e-26, 1.208691e-25, 
    -3.241489e-25, -1.730625e-25, 1.64822e-26, -1.977857e-25, 1.730626e-25, 
    1.07134e-25, 2.74703e-26, 4.395245e-26, 7.14227e-26, -7.416961e-26, 
    7.691675e-26, -3.735953e-25, 3.571138e-26, -8.241069e-26, 7.691675e-26, 
    4.94465e-26, -2.746971e-27, 1.675686e-25, -2.74702e-26, -1.758095e-25, 
    -1.016399e-25, -2.197619e-25, -3.845829e-26, -2.060268e-25, 
    -7.416961e-26, 1.64822e-26, -6.867557e-26, -2.554732e-25, -4.944639e-26, 
    2.582204e-25, 1.620745e-25, 3.571138e-26, -2.74702e-26, -3.021722e-26, 
    -1.263631e-25, -2.142679e-25, 1.840507e-25, 1.593275e-25, -2.417381e-25, 
    2.856906e-25, 1.181221e-25, -5.494044e-26, -9.889284e-26, -2.582203e-25, 
    -5.493996e-27, 1.593275e-25, -1.318571e-25, -1.867976e-25, -5.768747e-26, 
    -3.186548e-25, 5.494103e-27, 7.14227e-26, 4.669947e-26, -5.493996e-27, 
    1.291102e-25, -1.373507e-26, 3.296435e-26, -6.043449e-26, 1.565805e-25, 
    -1.867976e-25, 1.593275e-25, 5.768757e-26, 6.592865e-26, 2.747078e-27, 
    2.005329e-25, 2.966787e-25, -3.681013e-25, -7.691664e-26, -1.483393e-25, 
    2.19762e-25, 1.0164e-25, -1.620744e-25, 5.494055e-26, 2.472328e-26, 
    -2.637143e-25, 4.94465e-26, 5.351469e-32, 2.472323e-25, -9.889284e-26, 
    -3.845829e-26, 2.911847e-25, 9.065187e-26, -1.922912e-26, -2.527262e-25, 
    3.021733e-26, 2.14268e-25, 2.582204e-25, 6.592865e-26, -1.648214e-25, 
    1.785567e-25, -1.675685e-25, -2.197614e-26, -3.296424e-26, 1.098815e-26, 
    3.626073e-25, 3.84584e-26, -9.889284e-26, -9.889284e-26, -3.845829e-26 ;

 M_LITR3C_TO_LEACHING =
  -1.648212e-26, -3.983183e-26, 2.472325e-26, 7.004916e-26, -8.10372e-26, 
    -8.790477e-26, 1.92292e-26, -1.167485e-25, -4.395237e-26, -4.395237e-26, 
    -1.304836e-25, -8.378423e-26, 6.180808e-26, -1.098807e-26, -6.043452e-26, 
    -1.648212e-26, 8.241101e-27, 2.747028e-26, -7.829018e-26, -6.592857e-26, 
    -3.296427e-26, -5.768749e-26, -1.030134e-25, -1.112545e-25, -2.47232e-26, 
    -4.395237e-26, -5.906101e-26, 5.768755e-26, 7.279618e-26, 7.416969e-26, 
    -1.030134e-25, -2.47232e-26, 7.966375e-26, -7.554316e-26, -8.241071e-26, 
    2.884379e-26, -1.785563e-26, -1.304836e-25, -1.455923e-25, 1.002664e-25, 
    3.296432e-26, -6.043452e-26, 4.12054e-26, 2.884379e-26, -3.296427e-26, 
    4.669945e-26, -9.61456e-27, 3.296432e-26, -8.515774e-26, -3.159076e-26, 
    -6.455506e-26, 1.236161e-25, -2.747022e-26, -2.28003e-25, 2.334974e-26, 
    -1.620744e-25, -1.565804e-25, -9.614584e-26, 1.648217e-26, 2.197622e-26, 
    -6.180803e-26, -3.57113e-26, -7.142262e-26, 5.21935e-26, -8.378423e-26, 
    -5.356696e-26, 7.966375e-26, -1.030134e-25, -6.592857e-26, -9.20253e-26, 
    -1.593274e-25, -1.854241e-25, -1.785563e-26, 8.241101e-27, 1.181221e-25, 
    -4.120511e-27, 6.592862e-26, -6.318154e-26, 2.197622e-26, -1.098807e-26, 
    -2.197617e-26, -9.751935e-26, -1.66195e-25, -1.057604e-25, 6.867589e-27, 
    9.339887e-26, -2.197617e-26, -1.112545e-25, -1.208691e-25, -6.867535e-27, 
    -6.180803e-26, -8.378423e-26, -3.433778e-26, 6.592862e-26, -2.197617e-26, 
    -7.966369e-26, -2.746998e-27, 4.395242e-26, 6.31816e-26, -6.455506e-26, 
    -6.867535e-27, 1.373513e-25, 2.197622e-26, 2.884379e-26, 1.648217e-26, 
    1.744361e-25, 2.334974e-26, -1.565804e-25, -1.455923e-25, 1.304837e-25, 
    -1.922915e-26, -4.395237e-26, 3.433784e-26, 4.120564e-27, -2.211355e-25, 
    -1.12628e-25, -3.983183e-26, 4.257891e-26, -6.455506e-26, -6.455506e-26, 
    1.442188e-25, -3.433778e-26, -4.669939e-26, 1.552069e-25, -1.785563e-26, 
    -1.37351e-26, -1.222426e-25, 3.433784e-26, 1.373515e-26, -1.524598e-25, 
    -1.167485e-25, -1.057604e-25, 1.92292e-26, -4.120511e-27, -1.208691e-25, 
    1.318572e-25, -4.944642e-26, 1.648217e-26, -2.609671e-26, -6.592857e-26, 
    -9.477233e-26, -6.043452e-26, 3.571135e-26, -8.241047e-27, 1.648217e-26, 
    4.257891e-26, -7.416964e-26, -6.455506e-26, -1.442188e-25, -5.768749e-26, 
    2.675729e-32, 6.043457e-26, 3.159081e-26, 5.631404e-26, -5.768749e-26, 
    6.592862e-26, 1.552069e-25, 2.675744e-32, -6.867535e-27, 1.648215e-25, 
    -5.631398e-26, -4.944642e-26, -1.236161e-25, 1.785569e-26, -1.785563e-26, 
    2.197622e-26, -3.57113e-26, -4.395237e-26, 4.257891e-26, 7.004916e-26, 
    7.966375e-26, 3.02173e-26, -8.515774e-26, -6.867535e-27, 1.236164e-26, 
    6.455511e-26, -1.37351e-26, 1.332307e-25, -5.768749e-26, -2.747022e-26, 
    -6.867559e-26, -3.296427e-26, 9.065185e-26, 4.12054e-26, -7.966369e-26, 
    5.906106e-26, 7.142267e-26, -1.758096e-25, -4.532588e-26, -6.318154e-26, 
    7.829024e-26, 1.648217e-26, -7.966369e-26, -7.829018e-26, -2.197617e-26, 
    6.31816e-26, -1.510861e-26, 8.515779e-26, -1.922915e-26, -8.378423e-26, 
    1.208691e-25, 3.708486e-26, 1.085075e-25, -2.334968e-26, 1.181221e-25, 
    8.103726e-26, 3.433784e-26, -1.703155e-25, 3.296432e-26, 5.768755e-26, 
    -1.922915e-26, -1.703155e-25, 6.867565e-26, 3.845837e-26, 8.241077e-26, 
    -1.648212e-26, -1.922915e-26, -2.47232e-26, 1.455923e-25, 4.12054e-26, 
    9.75194e-26, -7.142262e-26, -3.159076e-26, 2.060271e-26, -2.747022e-26, 
    2.675739e-32, -8.241047e-27, -6.592857e-26, 7.966375e-26, -5.219344e-26, 
    -7.279613e-26, 4.395242e-26, -7.829018e-26, -3.296427e-26, -1.043869e-25, 
    1.373539e-27, 7.554321e-26, 7.691672e-26, -1.648215e-25, -8.241047e-27, 
    -9.61456e-27, -8.241047e-27, -1.37351e-26, 3.983189e-26, 8.653131e-26, 
    -5.768749e-26, -3.159076e-26, 1.236164e-26, 6.867589e-27, -7.00491e-26, 
    2.472325e-26, -1.538334e-25, -1.318572e-25, 3.983189e-26, -3.57113e-26, 
    2.472325e-26, 7.142267e-26, 2.609676e-26, -6.867559e-26, 3.845837e-26, 
    1.483394e-25, 2.609676e-26, 3.02173e-26, -8.241047e-27, -5.494023e-27, 
    -1.208691e-25, 2.884379e-26, -2.747022e-26, 5.494052e-26, 5.494076e-27, 
    2.472325e-26, -1.016399e-25, -1.799301e-25, 6.592862e-26, -1.043869e-25, 
    -1.881712e-25, 1.09881e-25, -5.768749e-26, -1.071339e-25, -5.768749e-26, 
    8.927833e-26, 3.708486e-26, 7.966375e-26, -6.180803e-26, 9.889292e-26, 
    1.263632e-25, -6.867535e-27, 2.197622e-26, 3.983189e-26, -1.593274e-25, 
    1.236161e-25, -6.043452e-26, -3.296427e-26, -6.043452e-26, 5.768755e-26, 
    6.043457e-26, -1.840506e-25, 1.909182e-25, 8.241101e-27, -1.098807e-26, 
    8.241101e-27, -9.889287e-26, -1.15375e-25, 5.494076e-27, -1.922915e-26, 
    2.747028e-26, -1.236158e-26, 5.906106e-26, -5.081993e-26, 1.167486e-25, 
    2.472325e-26, -6.043452e-26, -5.494023e-27, 8.790482e-26, -7.966369e-26, 
    -5.906101e-26, 4.532594e-26, -2.197617e-26, -1.318572e-25, -2.060266e-26, 
    4.944647e-26, 3.433784e-26, 1.92292e-26, 8.103726e-26, -1.098807e-26, 
    3.296432e-26, -9.889287e-26, 9.065185e-26, -2.334968e-26, 9.202536e-26, 
    -1.12628e-25, -9.339881e-26, -5.494047e-26, -3.433778e-26, -1.318572e-25, 
    2.472325e-26, 2.472325e-26, -3.021725e-26 ;

 M_SOIL1C_TO_LEACHING =
  -5.117639e-22, -1.429219e-21, 4.171381e-20, -4.010526e-21, 1.646285e-20, 
    1.943773e-20, 2.413334e-20, -1.059138e-20, -3.189486e-20, 4.076046e-20, 
    2.408386e-20, 3.096355e-20, 4.254542e-21, 2.105639e-20, -2.665529e-20, 
    2.948881e-20, -7.255447e-21, 2.095712e-20, -1.418857e-20, 1.411308e-20, 
    -2.657641e-20, 1.699491e-21, -2.98309e-21, 4.437741e-21, -1.199117e-20, 
    4.143052e-20, 9.485607e-21, 1.851095e-20, 3.393957e-20, -3.205035e-20, 
    -5.615712e-20, 1.00163e-20, -2.188421e-20, -3.511552e-22, -9.067112e-22, 
    -6.905981e-21, -3.59436e-21, -1.81434e-20, -3.356042e-20, 1.019357e-20, 
    2.014192e-21, 3.766141e-20, 1.075492e-21, 6.534758e-21, -3.624156e-20, 
    -5.077785e-22, -1.198723e-20, -1.050487e-20, -7.419696e-21, 
    -2.724307e-20, 3.407499e-20, 3.756446e-20, 2.317147e-20, 2.062515e-21, 
    -1.338363e-20, 9.187905e-21, 2.134447e-20, -1.395337e-20, 4.458269e-20, 
    -1.488406e-20, -2.597787e-20, -4.784256e-20, -3.9214e-22, 8.341127e-21, 
    4.424538e-20, 6.279579e-22, 5.354724e-20, 3.130309e-20, -1.571221e-20, 
    -1.553324e-20, -1.868313e-20, 4.55792e-21, 2.000518e-20, 8.145461e-21, 
    1.567318e-20, -4.380631e-21, 3.321437e-20, 1.807469e-20, 2.544466e-20, 
    -1.865731e-21, 3.064236e-20, 1.206354e-20, 4.21362e-20, -1.475431e-20, 
    -2.999215e-21, 2.185087e-20, -9.79012e-21, 9.791238e-21, 1.76181e-20, 
    -3.987635e-21, 1.684793e-20, 1.585638e-20, 8.940519e-21, 7.707805e-21, 
    6.129327e-21, -1.585951e-20, -2.935034e-21, -2.914616e-20, -9.969644e-21, 
    7.011667e-22, -3.214761e-20, -3.116088e-20, -4.80217e-21, 1.247887e-20, 
    -2.687183e-20, -2.407933e-20, -3.412787e-20, 3.575045e-20, 1.834979e-20, 
    5.195184e-21, -1.440824e-20, 2.710711e-20, 3.573575e-20, 7.083244e-21, 
    -1.025972e-20, -2.140528e-20, -6.873184e-21, -5.7171e-20, -1.97397e-20, 
    -7.113552e-22, -7.898931e-21, 1.36019e-20, 2.917499e-20, 1.010084e-20, 
    -2.310472e-21, -1.098381e-20, 1.182915e-20, 2.894427e-20, 1.138387e-20, 
    3.091492e-20, -1.972388e-20, 5.315111e-20, -8.68295e-21, 1.859266e-20, 
    -7.09371e-21, -2.101221e-21, -1.044011e-20, 4.136605e-20, -2.525068e-20, 
    -2.517985e-21, -2.116523e-20, 3.532998e-21, 1.729692e-20, -6.007458e-21, 
    6.236886e-22, -1.509783e-21, -1.763477e-20, -1.104093e-20, -2.909497e-20, 
    -8.788661e-21, -4.197423e-20, 2.844668e-20, 4.290158e-20, -2.405672e-20, 
    2.583426e-20, -1.208758e-20, 9.226375e-21, 5.00009e-21, 2.055169e-20, 
    6.708935e-21, -4.134673e-21, -3.395795e-20, -1.291826e-20, -2.338692e-20, 
    -2.212708e-20, -1.975497e-20, -4.362253e-21, 4.420976e-20, 3.672542e-22, 
    1.793815e-20, -4.785698e-20, -4.89917e-21, -2.376154e-20, -1.63226e-20, 
    -5.104082e-20, 2.253026e-20, 2.964347e-20, 2.079684e-20, -4.377807e-21, 
    -8.46836e-21, 4.418792e-21, 2.45105e-20, 1.021591e-20, 5.641322e-21, 
    1.462734e-20, 1.636786e-20, 6.691675e-21, -3.183564e-21, -3.187784e-21, 
    -6.768869e-21, 3.225138e-21, -2.434934e-20, 2.589646e-20, 1.443029e-20, 
    3.354912e-20, 6.49717e-21, 4.535737e-20, -1.392957e-20, -6.367113e-21, 
    -6.160622e-22, -1.582501e-20, 2.471636e-21, 6.926065e-21, 2.343355e-20, 
    -1.707439e-20, -1.509274e-20, 2.086326e-20, -9.68013e-21, 3.44875e-20, 
    2.574834e-21, -1.260443e-20, 2.635589e-20, -4.664487e-21, 1.306779e-21, 
    -6.538727e-21, 2.064841e-20, 7.118597e-21, -1.183765e-20, 2.144344e-20, 
    -3.564943e-21, 2.302192e-20, 4.507831e-20, 1.849938e-20, -2.182625e-20, 
    1.789261e-20, -2.114403e-20, 2.024041e-20, 1.935039e-20, 3.98596e-21, 
    1.31754e-21, 2.788488e-20, -1.548601e-20, -3.71316e-20, 1.690532e-20, 
    1.664946e-20, -2.29343e-20, -2.608727e-20, -5.728966e-21, 1.006579e-20, 
    1.284899e-20, 2.807603e-20, -6.768297e-21, 1.606188e-21, 8.155078e-21, 
    -1.6015e-20, -2.001988e-20, -4.481396e-20, -2.951681e-20, -1.646821e-20, 
    -3.762862e-21, -1.394069e-22, 1.729804e-20, 1.645466e-20, 2.449291e-21, 
    7.573234e-21, -8.772284e-21, -3.075546e-20, 1.84626e-20, -3.4401e-20, 
    5.459559e-20, 1.917253e-20, 1.293775e-20, 2.576583e-20, -5.249208e-21, 
    2.648903e-20, 1.888528e-20, -9.384116e-21, -1.486458e-20, -9.472054e-21, 
    2.207591e-20, -2.810598e-20, 4.784653e-20, 3.698911e-20, -3.981754e-20, 
    2.102693e-21, 2.607992e-20, -1.610435e-20, 2.498266e-20, 2.303519e-20, 
    -2.254785e-21, 5.999637e-22, -1.004456e-20, 1.926697e-20, -1.650357e-20, 
    -9.810546e-22, 1.597202e-20, 4.513512e-21, 3.579882e-20, -9.480065e-22, 
    5.945272e-21, -6.926327e-21, -8.052168e-21, -4.750163e-21, 8.550068e-21, 
    -8.145461e-21, 1.372461e-20, -1.583999e-20, -2.243526e-20, -3.671598e-20, 
    1.503762e-20, -2.298594e-21, -9.150031e-21, -4.0491e-20, 5.974662e-21, 
    4.024165e-20, 3.579908e-20, 1.045311e-20, 4.543532e-22, 1.340566e-20, 
    -7.012575e-21, -1.948838e-20, 2.787443e-20, 1.197676e-20, -1.368814e-20, 
    3.071362e-20, 1.416622e-20, -3.480973e-21, 4.573114e-20, 3.382958e-20, 
    2.590547e-20, -2.651026e-20, 1.435735e-20, 2.453567e-20, 2.812946e-20, 
    1.485836e-20, -1.824575e-20, -4.970117e-21, -1.469124e-20, -4.310801e-21, 
    1.400845e-20, -1.957657e-20, 3.944632e-20, 3.459918e-20, 3.557941e-20, 
    -2.006549e-21, -1.054049e-20, 9.894157e-21, -8.477121e-21 ;

 M_SOIL2C_TO_LEACHING =
  -1.154532e-20, 5.034276e-20, -5.961387e-21, -4.406062e-21, 4.280093e-20, 
    -1.905266e-20, -2.195094e-20, 4.186507e-20, 1.432852e-20, 8.489545e-21, 
    -1.303219e-20, -1.185603e-20, 1.436131e-20, -2.106061e-20, 3.693311e-21, 
    -2.335752e-20, -4.748436e-20, 2.116607e-20, -1.429459e-20, 5.967045e-21, 
    -1.779311e-20, -2.748155e-21, -2.289215e-20, -1.282607e-20, 
    -8.299008e-21, -3.699531e-21, -1.389395e-20, -1.817336e-20, 2.091653e-21, 
    -3.707363e-20, 2.146182e-20, -1.727822e-20, 1.223741e-20, 1.214894e-20, 
    1.811059e-20, -2.070889e-20, 4.814066e-21, -2.665529e-20, -4.586748e-21, 
    -1.720728e-20, -1.435255e-20, -1.587279e-20, 4.72559e-20, 3.274926e-20, 
    5.595523e-20, -1.808176e-20, -2.090398e-20, -8.298142e-21, 2.339317e-21, 
    1.783241e-20, 7.512227e-22, -2.385654e-20, 3.329411e-20, -3.011083e-20, 
    -1.361348e-21, 7.398778e-21, -1.324735e-20, -4.037101e-21, -1.066376e-20, 
    4.809526e-21, 9.389481e-21, 3.166387e-20, -2.593349e-20, -2.27587e-20, 
    1.260894e-20, -1.806933e-20, -4.308539e-21, -3.352371e-21, 3.40494e-21, 
    2.710314e-20, 3.083264e-20, -9.364621e-21, -4.684009e-21, 1.034507e-21, 
    -1.015795e-20, 3.702071e-21, -3.141337e-20, -1.005023e-20, 4.251718e-21, 
    -2.465554e-20, 1.478393e-21, -6.19576e-21, -1.28133e-21, -1.969615e-20, 
    -1.958872e-20, -1.238614e-20, -2.131735e-20, -2.973791e-20, 2.639516e-20, 
    9.182964e-22, 4.665986e-23, 2.564453e-20, -7.392167e-20, -2.453804e-21, 
    9.980112e-21, -2.007333e-20, -5.506472e-21, -5.310531e-20, 3.489465e-20, 
    3.965809e-20, 3.815564e-20, -2.429223e-21, 3.802898e-20, 6.378362e-22, 
    6.124046e-22, -2.019151e-20, 1.681571e-20, 2.159017e-20, 2.974667e-20, 
    5.654051e-21, 3.624835e-20, 2.443784e-20, -1.48558e-20, -2.319805e-21, 
    -2.294078e-20, 2.33139e-21, -7.449952e-21, 2.626202e-20, -1.587167e-20, 
    2.45317e-20, 4.677779e-21, 5.682324e-20, 4.005474e-20, -1.748124e-21, 
    1.885814e-20, -2.066961e-20, -5.763469e-21, -1.298553e-20, 2.865762e-21, 
    -1.758591e-21, 2.143862e-20, -3.153579e-20, 2.331963e-21, -6.675632e-22, 
    2.172841e-20, 4.231492e-20, -1.12753e-20, 3.812918e-21, -9.503985e-21, 
    3.245157e-20, -4.073923e-20, -2.03563e-20, -3.812061e-21, -1.309241e-20, 
    3.176367e-20, -1.775834e-21, 6.653231e-21, -5.077829e-21, -4.941844e-21, 
    1.041298e-20, 3.144702e-20, 5.325503e-21, -1.123261e-20, 2.841161e-20, 
    -2.75015e-20, 2.002101e-20, -3.851362e-21, -1.365139e-20, 5.698432e-21, 
    6.037169e-21, 6.06429e-21, -4.372442e-21, 3.012186e-20, 4.81601e-20, 
    -2.312315e-20, -4.304716e-20, -1.055662e-20, -4.731302e-20, 
    -1.145039e-22, -2.195122e-20, -1.163888e-20, -6.111512e-21, 7.102472e-21, 
    -8.734401e-21, -1.437288e-20, 3.345157e-20, 3.242639e-20, 8.640537e-21, 
    -1.905323e-20, 1.994654e-21, 2.087176e-20, -3.269103e-20, -2.63457e-20, 
    1.86803e-20, 2.516925e-20, 2.722698e-20, 1.832519e-20, -1.270569e-21, 
    2.448051e-20, 9.250889e-22, 2.335866e-20, 2.647041e-20, -9.507953e-21, 
    1.875779e-20, -1.503026e-20, 2.054606e-20, 3.578807e-21, 1.973753e-21, 
    -2.545057e-20, -3.457375e-20, -1.227391e-20, -7.075333e-21, 3.372611e-20, 
    6.456447e-21, 1.957996e-20, 9.039042e-22, 2.264899e-20, -2.356304e-20, 
    1.674105e-20, 1.157301e-20, 1.858984e-20, 1.563497e-21, 7.432137e-21, 
    1.752027e-20, -2.305959e-21, -4.868609e-22, -3.257614e-21, -5.306964e-22, 
    4.418262e-20, -9.175747e-21, 1.006011e-20, -1.425781e-20, 2.226503e-21, 
    -1.389338e-20, 3.297432e-20, 1.867973e-20, 2.318688e-21, 5.746798e-21, 
    -1.096513e-20, 2.506521e-20, -4.653978e-20, 1.447525e-20, -6.149672e-21, 
    3.735524e-20, -6.578878e-21, -1.233554e-20, -2.070832e-20, 2.493629e-20, 
    2.892336e-20, 1.916265e-20, -1.065754e-20, 1.69551e-20, -2.658151e-20, 
    2.604405e-20, 6.076437e-21, -5.273002e-22, -4.140299e-21, -5.23674e-21, 
    1.773294e-21, -1.684988e-20, -2.522834e-20, 1.519902e-20, 1.080794e-20, 
    3.105034e-20, -2.653032e-20, 1.142092e-20, 1.542155e-20, 3.379744e-21, 
    -3.194603e-21, -3.413068e-20, -1.292343e-21, 4.543484e-21, -1.888924e-20, 
    -1.586291e-20, -3.467699e-21, 4.244091e-21, 5.244079e-21, -1.151338e-20, 
    -5.591266e-21, 5.290738e-21, -2.9864e-20, -1.12736e-20, -5.768554e-21, 
    3.511941e-20, 3.518641e-20, 1.099257e-20, 4.440565e-21, -1.344187e-20, 
    -2.346326e-20, 1.349559e-20, -2.748709e-20, -2.929825e-20, -1.002789e-20, 
    -6.31366e-21, 6.459533e-21, -6.750492e-21, -4.052153e-20, 1.716176e-20, 
    1.146021e-20, 1.522365e-20, -8.527461e-21, 1.369546e-20, 1.767407e-20, 
    1.344243e-20, 5.314491e-20, -5.033741e-21, 2.670704e-20, 2.587128e-20, 
    -1.739249e-20, -9.762453e-22, -1.532599e-20, -2.768869e-20, 1.26604e-20, 
    -2.063255e-20, -1.38097e-20, 1.014239e-20, 3.021855e-20, 3.496361e-20, 
    -2.331257e-20, 1.210482e-20, -1.920703e-20, 3.724924e-20, -1.495589e-20, 
    4.385099e-20, 1.372402e-20, 1.410007e-20, -2.730503e-20, -1.42974e-20, 
    -2.595187e-20, 1.75152e-21, -7.927197e-21, 2.988176e-21, -6.72475e-21, 
    -1.008585e-20, 2.529224e-20, 3.797643e-21, -1.828843e-20, 1.399575e-20, 
    -7.668788e-21, 1.385976e-20, 1.998869e-22, 1.364232e-20, -2.417573e-20, 
    1.023457e-20, -1.096825e-20, -2.103941e-20, -2.31548e-20, 1.085911e-20 ;

 M_SOIL3C_TO_LEACHING =
  1.871481e-20, -1.851548e-20, 1.624768e-20, -1.195895e-20, -3.522268e-21, 
    1.453746e-20, -1.78013e-20, 1.301267e-20, 8.913926e-21, 6.904292e-21, 
    1.953924e-20, 2.310363e-20, -3.556753e-20, 1.829607e-20, -4.813266e-20, 
    5.457839e-21, -5.909079e-21, 1.448373e-20, 1.035473e-20, -2.445705e-20, 
    1.423605e-20, 1.743656e-20, 1.702577e-20, 1.137565e-20, 1.277262e-20, 
    -1.937159e-20, -1.034088e-20, 2.654836e-21, 4.646226e-20, 7.917025e-21, 
    -4.064453e-20, -3.837899e-20, -2.13159e-20, 2.363614e-21, -7.218404e-21, 
    2.485826e-20, 3.725535e-21, 1.474163e-21, -1.082321e-20, -2.272844e-20, 
    -2.163231e-20, -1.994213e-20, -1.964441e-20, 4.360301e-20, -1.331577e-20, 
    1.952708e-20, 3.146594e-20, -4.67812e-20, -1.20972e-20, 2.946281e-20, 
    -1.083425e-20, -2.931663e-20, 3.437412e-20, -4.453015e-21, 8.8128e-22, 
    -5.468573e-21, -6.707507e-21, -2.057771e-20, -1.390243e-20, 1.321344e-20, 
    -7.398206e-21, -1.565309e-20, -2.426509e-20, 1.130274e-20, -1.099088e-20, 
    -1.291061e-20, 3.720484e-20, 1.221455e-20, -6.619863e-21, -1.524029e-22, 
    -2.697026e-20, -4.551597e-20, -1.539046e-20, 4.721718e-20, 2.733719e-21, 
    1.235334e-20, -1.942585e-20, 2.412202e-20, -1.207091e-20, -3.339957e-20, 
    -2.369877e-20, -3.740542e-21, 4.673662e-22, -8.657208e-21, 1.512638e-20, 
    2.418773e-21, 9.954663e-21, -5.748682e-20, 2.346944e-21, 3.072124e-20, 
    -4.28207e-20, -1.332396e-20, 1.102924e-21, 2.818826e-20, 5.788067e-21, 
    3.386436e-20, 1.028859e-21, -2.650798e-20, -1.804586e-20, 5.1457e-21, 
    8.589909e-21, -1.941428e-20, -1.477269e-20, -2.942888e-20, -1.313567e-20, 
    -3.072833e-20, 3.194546e-20, -1.566921e-20, 6.442011e-21, -5.346731e-21, 
    1.266945e-20, -1.57088e-20, -1.887483e-20, 3.16384e-20, -1.880388e-20, 
    2.703867e-20, -2.611244e-20, 1.469438e-20, 6.011426e-21, 1.062756e-20, 
    1.391401e-20, 8.995088e-21, 1.881284e-21, 2.568243e-20, 6.809282e-21, 
    4.082263e-20, -1.373537e-20, -5.859023e-21, 5.818584e-21, -1.137765e-20, 
    -5.790607e-21, 1.232338e-20, -1.19222e-20, 1.980106e-20, 1.035133e-20, 
    4.153796e-20, -1.835912e-20, 3.522968e-20, 1.191711e-20, -4.43794e-20, 
    -1.49381e-20, -1.165811e-20, -4.136052e-21, -9.745739e-21, -4.625192e-21, 
    -2.454443e-20, -8.459306e-21, 6.671298e-21, -4.949488e-21, -6.172018e-21, 
    -1.320637e-20, -5.386066e-22, 2.730895e-21, -3.29322e-20, 7.284013e-21, 
    1.839165e-21, -2.453764e-20, 1.383741e-20, -2.632197e-20, -1.695054e-20, 
    -2.426112e-20, -7.209904e-21, -3.926763e-20, 1.022298e-20, 5.764596e-20, 
    3.809345e-20, -3.373262e-21, -3.79411e-22, -2.691511e-20, -1.126485e-20, 
    3.092396e-20, 3.659969e-21, 1.700767e-20, 2.733979e-20, -1.239464e-20, 
    -3.608494e-20, -1.10576e-20, 6.139794e-21, 2.486787e-20, -8.934366e-22, 
    -5.067639e-20, -1.258999e-20, -1.072087e-20, 5.250326e-21, 3.890095e-21, 
    3.047018e-20, -2.037066e-21, 2.560832e-20, -7.278338e-21, -2.299649e-20, 
    2.510932e-21, -4.119381e-21, 1.260555e-20, -1.169967e-20, -1.41812e-20, 
    1.534919e-20, 4.86133e-20, -2.458062e-20, -4.866448e-20, 6.360041e-21, 
    -1.575947e-21, 2.869093e-20, 3.581264e-20, 4.211278e-21, 4.738031e-20, 
    1.11964e-22, -1.877926e-20, -1.001913e-20, -1.178721e-21, 8.136727e-21, 
    2.163745e-21, -5.085193e-21, -2.773645e-20, -2.056216e-20, -3.064807e-21, 
    3.034746e-20, 3.122931e-20, 1.311138e-20, -4.932245e-21, 1.520102e-20, 
    -1.080597e-20, 1.875182e-20, 7.427051e-21, -1.255606e-20, 1.326846e-21, 
    -9.148609e-21, -2.072558e-20, 1.435481e-20, 2.563943e-20, 1.007087e-20, 
    6.805314e-21, -8.001173e-22, 5.17341e-21, 9.226921e-21, -2.659254e-20, 
    6.019615e-21, -1.044802e-20, -5.397246e-20, 1.022861e-20, 3.386836e-20, 
    7.522606e-21, -1.440484e-20, 6.519777e-21, -4.562625e-20, -7.635992e-21, 
    3.663004e-20, 5.737465e-21, 1.267114e-20, -3.152164e-21, -2.819395e-21, 
    4.763438e-21, 2.492384e-20, -2.152627e-20, 6.722488e-21, -1.140761e-20, 
    -2.318502e-20, -3.092142e-20, 1.273966e-21, 2.896018e-21, 3.729782e-21, 
    2.531572e-20, 1.364799e-20, -1.760393e-20, -8.875792e-21, 3.254542e-20, 
    -1.424028e-20, 3.275548e-20, -4.356578e-21, -2.173181e-20, 2.300976e-20, 
    -2.316159e-20, 2.632253e-20, 5.355403e-20, -2.837656e-20, -1.212094e-20, 
    -1.781118e-20, 8.846937e-21, 2.998418e-20, 1.435255e-20, 1.667461e-20, 
    -6.339974e-21, -1.329626e-20, 1.859294e-20, -1.868791e-22, -1.059817e-20, 
    -4.666498e-20, 1.664465e-20, -3.218948e-20, -1.636162e-20, 3.012948e-20, 
    9.783334e-23, -1.661551e-20, 5.488919e-21, -4.913211e-20, -1.337062e-20, 
    -2.54992e-20, -2.691908e-20, 1.497963e-20, -2.093509e-20, 2.798757e-21, 
    -2.339872e-21, -1.016134e-20, -3.913136e-20, 7.887608e-21, 4.457236e-21, 
    -8.227991e-23, 9.995093e-21, -1.373024e-20, -1.325728e-21, -8.786147e-21, 
    4.137538e-20, -2.664168e-21, 1.184893e-21, 1.807979e-20, -1.092584e-20, 
    2.30697e-20, -7.681517e-21, 8.244315e-22, 5.963077e-21, -1.565623e-20, 
    -1.086139e-20, -5.648686e-21, -1.854718e-21, -2.458005e-20, 2.370407e-21, 
    -7.506503e-22, -1.619311e-20, -4.774645e-20, 2.794992e-20, 5.408188e-20, 
    -2.795754e-20, 5.05158e-20, 2.432981e-20, -2.483959e-20, 2.260858e-20, 
    -3.145438e-20, 2.175416e-20, -3.913758e-20 ;

 NBP =
  -6.191209e-08, -6.218511e-08, -6.213204e-08, -6.235225e-08, -6.22301e-08, 
    -6.237429e-08, -6.196745e-08, -6.219594e-08, -6.205008e-08, 
    -6.193667e-08, -6.277961e-08, -6.236208e-08, -6.321343e-08, -6.29471e-08, 
    -6.361618e-08, -6.317198e-08, -6.370576e-08, -6.360339e-08, 
    -6.391155e-08, -6.382326e-08, -6.421742e-08, -6.39523e-08, -6.442178e-08, 
    -6.415411e-08, -6.419598e-08, -6.394355e-08, -6.244612e-08, 
    -6.272763e-08, -6.242944e-08, -6.246958e-08, -6.245157e-08, 
    -6.223262e-08, -6.212228e-08, -6.189123e-08, -6.193318e-08, 
    -6.210288e-08, -6.248763e-08, -6.235703e-08, -6.26862e-08, -6.267877e-08, 
    -6.304526e-08, -6.288002e-08, -6.349605e-08, -6.332096e-08, 
    -6.382695e-08, -6.369969e-08, -6.382097e-08, -6.37842e-08, -6.382145e-08, 
    -6.363481e-08, -6.371478e-08, -6.355055e-08, -6.291096e-08, 
    -6.309892e-08, -6.253835e-08, -6.220129e-08, -6.197747e-08, 
    -6.181863e-08, -6.184109e-08, -6.188389e-08, -6.210387e-08, 
    -6.231072e-08, -6.246836e-08, -6.25738e-08, -6.267771e-08, -6.299219e-08, 
    -6.315867e-08, -6.353144e-08, -6.346419e-08, -6.357814e-08, 
    -6.368703e-08, -6.386984e-08, -6.383975e-08, -6.392029e-08, 
    -6.357515e-08, -6.380452e-08, -6.342587e-08, -6.352943e-08, -6.27059e-08, 
    -6.239227e-08, -6.225892e-08, -6.214224e-08, -6.185834e-08, 
    -6.205439e-08, -6.19771e-08, -6.216099e-08, -6.227782e-08, -6.222004e-08, 
    -6.257669e-08, -6.243803e-08, -6.316854e-08, -6.285387e-08, 
    -6.367434e-08, -6.347799e-08, -6.372139e-08, -6.359719e-08, 
    -6.381001e-08, -6.361848e-08, -6.395027e-08, -6.402251e-08, 
    -6.397314e-08, -6.41628e-08, -6.360786e-08, -6.382096e-08, -6.221842e-08, 
    -6.222784e-08, -6.227175e-08, -6.207874e-08, -6.206693e-08, 
    -6.189008e-08, -6.204745e-08, -6.211446e-08, -6.22846e-08, -6.238523e-08, 
    -6.248089e-08, -6.269123e-08, -6.292615e-08, -6.325467e-08, 
    -6.349072e-08, -6.364895e-08, -6.355192e-08, -6.363758e-08, 
    -6.354183e-08, -6.349695e-08, -6.399544e-08, -6.371552e-08, 
    -6.413553e-08, -6.411229e-08, -6.39222e-08, -6.411491e-08, -6.223446e-08, 
    -6.218023e-08, -6.199193e-08, -6.213929e-08, -6.187082e-08, 
    -6.202109e-08, -6.210749e-08, -6.244091e-08, -6.251418e-08, 
    -6.258211e-08, -6.271628e-08, -6.288847e-08, -6.319055e-08, -6.34534e-08, 
    -6.369337e-08, -6.367579e-08, -6.368198e-08, -6.373558e-08, -6.36028e-08, 
    -6.375738e-08, -6.378333e-08, -6.371549e-08, -6.410917e-08, -6.39967e-08, 
    -6.411179e-08, -6.403856e-08, -6.219786e-08, -6.228911e-08, -6.22398e-08, 
    -6.233252e-08, -6.22672e-08, -6.255767e-08, -6.264477e-08, -6.305234e-08, 
    -6.288508e-08, -6.315129e-08, -6.291213e-08, -6.29545e-08, -6.315996e-08, 
    -6.292505e-08, -6.34389e-08, -6.30905e-08, -6.373767e-08, -6.338972e-08, 
    -6.375947e-08, -6.369233e-08, -6.38035e-08, -6.390305e-08, -6.402831e-08, 
    -6.425942e-08, -6.420591e-08, -6.43992e-08, -6.242516e-08, -6.254352e-08, 
    -6.25331e-08, -6.265698e-08, -6.27486e-08, -6.294718e-08, -6.326568e-08, 
    -6.314591e-08, -6.33658e-08, -6.340995e-08, -6.307588e-08, -6.328098e-08, 
    -6.262274e-08, -6.272907e-08, -6.266577e-08, -6.243449e-08, 
    -6.317349e-08, -6.279422e-08, -6.349462e-08, -6.328914e-08, 
    -6.388886e-08, -6.359058e-08, -6.417645e-08, -6.442689e-08, 
    -6.466265e-08, -6.493813e-08, -6.260812e-08, -6.25277e-08, -6.267172e-08, 
    -6.287096e-08, -6.305586e-08, -6.330166e-08, -6.332682e-08, 
    -6.337287e-08, -6.349217e-08, -6.359246e-08, -6.338743e-08, 
    -6.361761e-08, -6.275372e-08, -6.320642e-08, -6.249729e-08, -6.27108e-08, 
    -6.285921e-08, -6.279412e-08, -6.313223e-08, -6.321191e-08, 
    -6.353574e-08, -6.336835e-08, -6.436507e-08, -6.392407e-08, 
    -6.514793e-08, -6.480587e-08, -6.249959e-08, -6.260785e-08, 
    -6.298463e-08, -6.280536e-08, -6.331808e-08, -6.344429e-08, -6.35469e-08, 
    -6.367805e-08, -6.369222e-08, -6.376993e-08, -6.364259e-08, 
    -6.376491e-08, -6.330219e-08, -6.350896e-08, -6.294157e-08, 
    -6.307966e-08, -6.301614e-08, -6.294646e-08, -6.316152e-08, 
    -6.339064e-08, -6.339556e-08, -6.346902e-08, -6.367603e-08, 
    -6.332016e-08, -6.442196e-08, -6.374147e-08, -6.27259e-08, -6.293441e-08, 
    -6.296421e-08, -6.288344e-08, -6.343164e-08, -6.3233e-08, -6.376804e-08, 
    -6.362344e-08, -6.386038e-08, -6.374263e-08, -6.372531e-08, 
    -6.357409e-08, -6.347994e-08, -6.32421e-08, -6.304859e-08, -6.289515e-08, 
    -6.293084e-08, -6.309938e-08, -6.340467e-08, -6.36935e-08, -6.363022e-08, 
    -6.384236e-08, -6.32809e-08, -6.351632e-08, -6.342533e-08, -6.36626e-08, 
    -6.314273e-08, -6.358538e-08, -6.302958e-08, -6.307831e-08, 
    -6.322905e-08, -6.353228e-08, -6.359939e-08, -6.367102e-08, 
    -6.362682e-08, -6.341242e-08, -6.33773e-08, -6.322539e-08, -6.318344e-08, 
    -6.30677e-08, -6.297188e-08, -6.305942e-08, -6.315137e-08, -6.341251e-08, 
    -6.364786e-08, -6.390447e-08, -6.396727e-08, -6.426707e-08, -6.4023e-08, 
    -6.442575e-08, -6.40833e-08, -6.467612e-08, -6.361105e-08, -6.407326e-08, 
    -6.323592e-08, -6.332613e-08, -6.348927e-08, -6.386351e-08, 
    -6.366148e-08, -6.389776e-08, -6.337593e-08, -6.310519e-08, 
    -6.303516e-08, -6.290448e-08, -6.303815e-08, -6.302728e-08, 
    -6.315518e-08, -6.311409e-08, -6.342119e-08, -6.325622e-08, 
    -6.372487e-08, -6.38959e-08, -6.437893e-08, -6.467506e-08, -6.497654e-08, 
    -6.510964e-08, -6.515015e-08, -6.516709e-08 ;

 NDEPLOY =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NDEP_TO_SMINN =
  3.989144e-10, 3.989147e-10, 3.989121e-10, 3.989123e-10, 3.989108e-10, 
    3.989089e-10, 3.989084e-10, 3.989066e-10, 3.98906e-10, 3.989042e-10, 
    3.989026e-10, 3.989029e-10, 3.989014e-10, 3.988995e-10, 3.988979e-10, 
    3.988982e-10, 3.988966e-10, 3.988948e-10, 3.988943e-10, 3.988924e-10, 
    3.988909e-10, 3.988911e-10, 3.988885e-10, 3.988888e-10, 3.988872e-10, 
    3.988854e-10, 3.989112e-10, 3.989115e-10, 3.989089e-10, 3.989092e-10, 
    3.989076e-10, 3.989057e-10, 3.989052e-10, 3.989034e-10, 3.989018e-10, 
    3.989021e-10, 3.989005e-10, 3.988987e-10, 3.988971e-10, 3.988974e-10, 
    3.988947e-10, 3.98895e-10, 3.988934e-10, 3.988916e-10, 3.988911e-10, 
    3.988892e-10, 3.988887e-10, 3.988869e-10, 3.988853e-10, 3.988856e-10, 
    3.98883e-10, 3.988832e-10, 3.989091e-10, 3.989072e-10, 3.989067e-10, 
    3.989049e-10, 3.989033e-10, 3.989036e-10, 3.98901e-10, 3.989012e-10, 
    3.988997e-10, 3.988978e-10, 3.988973e-10, 3.988955e-10, 3.988939e-10, 
    3.988942e-10, 3.988926e-10, 3.988908e-10, 3.988903e-10, 3.988884e-10, 
    3.988879e-10, 3.98886e-10, 3.988855e-10, 3.988837e-10, 3.988821e-10, 
    3.988824e-10, 3.988798e-10, 3.9888e-10, 3.989059e-10, 3.98904e-10, 
    3.989035e-10, 3.989017e-10, 3.989001e-10, 3.989004e-10, 3.988988e-10, 
    3.98897e-10, 3.988965e-10, 3.988946e-10, 3.988941e-10, 3.988923e-10, 
    3.988907e-10, 3.98891e-10, 3.988894e-10, 3.988876e-10, 3.98886e-10, 
    3.988863e-10, 3.988836e-10, 3.988839e-10, 3.988813e-10, 3.988816e-10, 
    3.988789e-10, 3.988792e-10, 3.988766e-10, 3.988768e-10, 3.989017e-10, 
    3.989019e-10, 3.989004e-10, 3.988985e-10, 3.98898e-10, 3.988962e-10, 
    3.988946e-10, 3.988949e-10, 3.988933e-10, 3.988914e-10, 3.988899e-10, 
    3.988901e-10, 3.988886e-10, 3.988867e-10, 3.988862e-10, 3.988844e-10, 
    3.988839e-10, 3.98882e-10, 3.988815e-10, 3.988797e-10, 3.988781e-10, 
    3.988784e-10, 3.988757e-10, 3.98876e-10, 3.988744e-10, 3.988726e-10, 
    3.988995e-10, 3.988977e-10, 3.988972e-10, 3.988953e-10, 3.988938e-10, 
    3.98894e-10, 3.988924e-10, 3.988906e-10, 3.98889e-10, 3.988893e-10, 
    3.988878e-10, 3.988859e-10, 3.988854e-10, 3.988835e-10, 3.98883e-10, 
    3.988812e-10, 3.988807e-10, 3.988788e-10, 3.988783e-10, 3.988765e-10, 
    3.988749e-10, 3.988752e-10, 3.988725e-10, 3.988728e-10, 3.988712e-10, 
    3.988694e-10, 3.988963e-10, 3.988945e-10, 3.988929e-10, 3.988932e-10, 
    3.988906e-10, 3.988908e-10, 3.988893e-10, 3.988874e-10, 3.988858e-10, 
    3.988861e-10, 3.988835e-10, 3.988838e-10, 3.988822e-10, 3.988803e-10, 
    3.988798e-10, 3.98878e-10, 3.988775e-10, 3.988756e-10, 3.988751e-10, 
    3.988733e-10, 3.988717e-10, 3.98872e-10, 3.988694e-10, 3.988696e-10, 
    3.98867e-10, 3.988673e-10, 3.988931e-10, 3.988913e-10, 3.988908e-10, 
    3.988889e-10, 3.988874e-10, 3.988876e-10, 3.988861e-10, 3.988842e-10, 
    3.988826e-10, 3.988829e-10, 3.988803e-10, 3.988806e-10, 3.98879e-10, 
    3.988772e-10, 3.988767e-10, 3.988748e-10, 3.988743e-10, 3.988724e-10, 
    3.988719e-10, 3.988701e-10, 3.988685e-10, 3.988688e-10, 3.988662e-10, 
    3.988664e-10, 3.988649e-10, 3.98863e-10, 3.988899e-10, 3.988881e-10, 
    3.988865e-10, 3.988868e-10, 3.988842e-10, 3.988845e-10, 3.988829e-10, 
    3.98881e-10, 3.988795e-10, 3.988797e-10, 3.988782e-10, 3.988763e-10, 
    3.988758e-10, 3.98874e-10, 3.988724e-10, 3.988727e-10, 3.9887e-10, 
    3.988703e-10, 3.988687e-10, 3.988669e-10, 3.988653e-10, 3.988656e-10, 
    3.98863e-10, 3.988632e-10, 3.988606e-10, 3.988609e-10, 3.988868e-10, 
    3.988849e-10, 3.988833e-10, 3.988836e-10, 3.98881e-10, 3.988813e-10, 
    3.988786e-10, 3.988789e-10, 3.988763e-10, 3.988765e-10, 3.988739e-10, 
    3.988742e-10, 3.988716e-10, 3.988719e-10, 3.988703e-10, 3.988684e-10, 
    3.988679e-10, 3.988661e-10, 3.988645e-10, 3.988648e-10, 3.988632e-10, 
    3.988614e-10, 3.988609e-10, 3.98859e-10, 3.988585e-10, 3.988566e-10, 
    3.988836e-10, 3.988817e-10, 3.988802e-10, 3.988804e-10, 3.988778e-10, 
    3.988781e-10, 3.988765e-10, 3.988747e-10, 3.988731e-10, 3.988734e-10, 
    3.988707e-10, 3.98871e-10, 3.988684e-10, 3.988687e-10, 3.98866e-10, 
    3.988663e-10, 3.988637e-10, 3.988639e-10, 3.988613e-10, 3.988616e-10, 
    3.9886e-10, 3.988582e-10, 3.988566e-10, 3.988569e-10, 3.988542e-10, 
    3.988545e-10, 3.988793e-10, 3.988796e-10, 3.98878e-10, 3.988762e-10, 
    3.988746e-10, 3.988749e-10, 3.988722e-10, 3.988725e-10, 3.988699e-10, 
    3.988702e-10, 3.988686e-10, 3.988667e-10, 3.988652e-10, 3.988655e-10, 
    3.988628e-10, 3.988631e-10, 3.988605e-10, 3.988607e-10, 3.988592e-10, 
    3.988573e-10, 3.988568e-10, 3.98855e-10, 3.988545e-10, 3.988526e-10, 
    3.988521e-10, 3.988503e-10, 3.988761e-10, 3.988764e-10, 3.988748e-10, 
    3.98873e-10, 3.988725e-10, 3.988706e-10, 3.98869e-10, 3.988693e-10, 
    3.988678e-10, 3.988659e-10, 3.988644e-10, 3.988646e-10, 3.98862e-10, 
    3.988623e-10, 3.988607e-10, 3.988589e-10, 3.988573e-10, 3.988576e-10, 
    3.988549e-10, 3.988552e-10, 3.988536e-10, 3.988518e-10, 3.988513e-10, 
    3.988494e-10, 3.988489e-10, 3.988476e-10 ;

 NEE =
  6.191209e-08, 6.218511e-08, 6.213204e-08, 6.235225e-08, 6.22301e-08, 
    6.237429e-08, 6.196745e-08, 6.219594e-08, 6.205008e-08, 6.193667e-08, 
    6.277961e-08, 6.236208e-08, 6.321343e-08, 6.29471e-08, 6.361618e-08, 
    6.317198e-08, 6.370576e-08, 6.360339e-08, 6.391155e-08, 6.382326e-08, 
    6.421742e-08, 6.39523e-08, 6.442178e-08, 6.415411e-08, 6.419598e-08, 
    6.394355e-08, 6.244612e-08, 6.272763e-08, 6.242944e-08, 6.246958e-08, 
    6.245157e-08, 6.223262e-08, 6.212228e-08, 6.189123e-08, 6.193318e-08, 
    6.210288e-08, 6.248763e-08, 6.235703e-08, 6.26862e-08, 6.267877e-08, 
    6.304526e-08, 6.288002e-08, 6.349605e-08, 6.332096e-08, 6.382695e-08, 
    6.369969e-08, 6.382097e-08, 6.37842e-08, 6.382145e-08, 6.363481e-08, 
    6.371478e-08, 6.355055e-08, 6.291096e-08, 6.309892e-08, 6.253835e-08, 
    6.220129e-08, 6.197747e-08, 6.181863e-08, 6.184109e-08, 6.188389e-08, 
    6.210387e-08, 6.231072e-08, 6.246836e-08, 6.25738e-08, 6.267771e-08, 
    6.299219e-08, 6.315867e-08, 6.353144e-08, 6.346419e-08, 6.357814e-08, 
    6.368703e-08, 6.386984e-08, 6.383975e-08, 6.392029e-08, 6.357515e-08, 
    6.380452e-08, 6.342587e-08, 6.352943e-08, 6.27059e-08, 6.239227e-08, 
    6.225892e-08, 6.214224e-08, 6.185834e-08, 6.205439e-08, 6.19771e-08, 
    6.216099e-08, 6.227782e-08, 6.222004e-08, 6.257669e-08, 6.243803e-08, 
    6.316854e-08, 6.285387e-08, 6.367434e-08, 6.347799e-08, 6.372139e-08, 
    6.359719e-08, 6.381001e-08, 6.361848e-08, 6.395027e-08, 6.402251e-08, 
    6.397314e-08, 6.41628e-08, 6.360786e-08, 6.382096e-08, 6.221842e-08, 
    6.222784e-08, 6.227175e-08, 6.207874e-08, 6.206693e-08, 6.189008e-08, 
    6.204745e-08, 6.211446e-08, 6.22846e-08, 6.238523e-08, 6.248089e-08, 
    6.269123e-08, 6.292615e-08, 6.325467e-08, 6.349072e-08, 6.364895e-08, 
    6.355192e-08, 6.363758e-08, 6.354183e-08, 6.349695e-08, 6.399544e-08, 
    6.371552e-08, 6.413553e-08, 6.411229e-08, 6.39222e-08, 6.411491e-08, 
    6.223446e-08, 6.218023e-08, 6.199193e-08, 6.213929e-08, 6.187082e-08, 
    6.202109e-08, 6.210749e-08, 6.244091e-08, 6.251418e-08, 6.258211e-08, 
    6.271628e-08, 6.288847e-08, 6.319055e-08, 6.34534e-08, 6.369337e-08, 
    6.367579e-08, 6.368198e-08, 6.373558e-08, 6.36028e-08, 6.375738e-08, 
    6.378333e-08, 6.371549e-08, 6.410917e-08, 6.39967e-08, 6.411179e-08, 
    6.403856e-08, 6.219786e-08, 6.228911e-08, 6.22398e-08, 6.233252e-08, 
    6.22672e-08, 6.255767e-08, 6.264477e-08, 6.305234e-08, 6.288508e-08, 
    6.315129e-08, 6.291213e-08, 6.29545e-08, 6.315996e-08, 6.292505e-08, 
    6.34389e-08, 6.30905e-08, 6.373767e-08, 6.338972e-08, 6.375947e-08, 
    6.369233e-08, 6.38035e-08, 6.390305e-08, 6.402831e-08, 6.425942e-08, 
    6.420591e-08, 6.43992e-08, 6.242516e-08, 6.254352e-08, 6.25331e-08, 
    6.265698e-08, 6.27486e-08, 6.294718e-08, 6.326568e-08, 6.314591e-08, 
    6.33658e-08, 6.340995e-08, 6.307588e-08, 6.328098e-08, 6.262274e-08, 
    6.272907e-08, 6.266577e-08, 6.243449e-08, 6.317349e-08, 6.279422e-08, 
    6.349462e-08, 6.328914e-08, 6.388886e-08, 6.359058e-08, 6.417645e-08, 
    6.442689e-08, 6.466265e-08, 6.493813e-08, 6.260812e-08, 6.25277e-08, 
    6.267172e-08, 6.287096e-08, 6.305586e-08, 6.330166e-08, 6.332682e-08, 
    6.337287e-08, 6.349217e-08, 6.359246e-08, 6.338743e-08, 6.361761e-08, 
    6.275372e-08, 6.320642e-08, 6.249729e-08, 6.27108e-08, 6.285921e-08, 
    6.279412e-08, 6.313223e-08, 6.321191e-08, 6.353574e-08, 6.336835e-08, 
    6.436507e-08, 6.392407e-08, 6.514793e-08, 6.480587e-08, 6.249959e-08, 
    6.260785e-08, 6.298463e-08, 6.280536e-08, 6.331808e-08, 6.344429e-08, 
    6.35469e-08, 6.367805e-08, 6.369222e-08, 6.376993e-08, 6.364259e-08, 
    6.376491e-08, 6.330219e-08, 6.350896e-08, 6.294157e-08, 6.307966e-08, 
    6.301614e-08, 6.294646e-08, 6.316152e-08, 6.339064e-08, 6.339556e-08, 
    6.346902e-08, 6.367603e-08, 6.332016e-08, 6.442196e-08, 6.374147e-08, 
    6.27259e-08, 6.293441e-08, 6.296421e-08, 6.288344e-08, 6.343164e-08, 
    6.3233e-08, 6.376804e-08, 6.362344e-08, 6.386038e-08, 6.374263e-08, 
    6.372531e-08, 6.357409e-08, 6.347994e-08, 6.32421e-08, 6.304859e-08, 
    6.289515e-08, 6.293084e-08, 6.309938e-08, 6.340467e-08, 6.36935e-08, 
    6.363022e-08, 6.384236e-08, 6.32809e-08, 6.351632e-08, 6.342533e-08, 
    6.36626e-08, 6.314273e-08, 6.358538e-08, 6.302958e-08, 6.307831e-08, 
    6.322905e-08, 6.353228e-08, 6.359939e-08, 6.367102e-08, 6.362682e-08, 
    6.341242e-08, 6.33773e-08, 6.322539e-08, 6.318344e-08, 6.30677e-08, 
    6.297188e-08, 6.305942e-08, 6.315137e-08, 6.341251e-08, 6.364786e-08, 
    6.390447e-08, 6.396727e-08, 6.426707e-08, 6.4023e-08, 6.442575e-08, 
    6.40833e-08, 6.467612e-08, 6.361105e-08, 6.407326e-08, 6.323592e-08, 
    6.332613e-08, 6.348927e-08, 6.386351e-08, 6.366148e-08, 6.389776e-08, 
    6.337593e-08, 6.310519e-08, 6.303516e-08, 6.290448e-08, 6.303815e-08, 
    6.302728e-08, 6.315518e-08, 6.311409e-08, 6.342119e-08, 6.325622e-08, 
    6.372487e-08, 6.38959e-08, 6.437893e-08, 6.467506e-08, 6.497654e-08, 
    6.510964e-08, 6.515015e-08, 6.516709e-08 ;

 NEM =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NEP =
  -6.191209e-08, -6.218511e-08, -6.213204e-08, -6.235225e-08, -6.22301e-08, 
    -6.237429e-08, -6.196745e-08, -6.219594e-08, -6.205008e-08, 
    -6.193667e-08, -6.277961e-08, -6.236208e-08, -6.321343e-08, -6.29471e-08, 
    -6.361618e-08, -6.317198e-08, -6.370576e-08, -6.360339e-08, 
    -6.391155e-08, -6.382326e-08, -6.421742e-08, -6.39523e-08, -6.442178e-08, 
    -6.415411e-08, -6.419598e-08, -6.394355e-08, -6.244612e-08, 
    -6.272763e-08, -6.242944e-08, -6.246958e-08, -6.245157e-08, 
    -6.223262e-08, -6.212228e-08, -6.189123e-08, -6.193318e-08, 
    -6.210288e-08, -6.248763e-08, -6.235703e-08, -6.26862e-08, -6.267877e-08, 
    -6.304526e-08, -6.288002e-08, -6.349605e-08, -6.332096e-08, 
    -6.382695e-08, -6.369969e-08, -6.382097e-08, -6.37842e-08, -6.382145e-08, 
    -6.363481e-08, -6.371478e-08, -6.355055e-08, -6.291096e-08, 
    -6.309892e-08, -6.253835e-08, -6.220129e-08, -6.197747e-08, 
    -6.181863e-08, -6.184109e-08, -6.188389e-08, -6.210387e-08, 
    -6.231072e-08, -6.246836e-08, -6.25738e-08, -6.267771e-08, -6.299219e-08, 
    -6.315867e-08, -6.353144e-08, -6.346419e-08, -6.357814e-08, 
    -6.368703e-08, -6.386984e-08, -6.383975e-08, -6.392029e-08, 
    -6.357515e-08, -6.380452e-08, -6.342587e-08, -6.352943e-08, -6.27059e-08, 
    -6.239227e-08, -6.225892e-08, -6.214224e-08, -6.185834e-08, 
    -6.205439e-08, -6.19771e-08, -6.216099e-08, -6.227782e-08, -6.222004e-08, 
    -6.257669e-08, -6.243803e-08, -6.316854e-08, -6.285387e-08, 
    -6.367434e-08, -6.347799e-08, -6.372139e-08, -6.359719e-08, 
    -6.381001e-08, -6.361848e-08, -6.395027e-08, -6.402251e-08, 
    -6.397314e-08, -6.41628e-08, -6.360786e-08, -6.382096e-08, -6.221842e-08, 
    -6.222784e-08, -6.227175e-08, -6.207874e-08, -6.206693e-08, 
    -6.189008e-08, -6.204745e-08, -6.211446e-08, -6.22846e-08, -6.238523e-08, 
    -6.248089e-08, -6.269123e-08, -6.292615e-08, -6.325467e-08, 
    -6.349072e-08, -6.364895e-08, -6.355192e-08, -6.363758e-08, 
    -6.354183e-08, -6.349695e-08, -6.399544e-08, -6.371552e-08, 
    -6.413553e-08, -6.411229e-08, -6.39222e-08, -6.411491e-08, -6.223446e-08, 
    -6.218023e-08, -6.199193e-08, -6.213929e-08, -6.187082e-08, 
    -6.202109e-08, -6.210749e-08, -6.244091e-08, -6.251418e-08, 
    -6.258211e-08, -6.271628e-08, -6.288847e-08, -6.319055e-08, -6.34534e-08, 
    -6.369337e-08, -6.367579e-08, -6.368198e-08, -6.373558e-08, -6.36028e-08, 
    -6.375738e-08, -6.378333e-08, -6.371549e-08, -6.410917e-08, -6.39967e-08, 
    -6.411179e-08, -6.403856e-08, -6.219786e-08, -6.228911e-08, -6.22398e-08, 
    -6.233252e-08, -6.22672e-08, -6.255767e-08, -6.264477e-08, -6.305234e-08, 
    -6.288508e-08, -6.315129e-08, -6.291213e-08, -6.29545e-08, -6.315996e-08, 
    -6.292505e-08, -6.34389e-08, -6.30905e-08, -6.373767e-08, -6.338972e-08, 
    -6.375947e-08, -6.369233e-08, -6.38035e-08, -6.390305e-08, -6.402831e-08, 
    -6.425942e-08, -6.420591e-08, -6.43992e-08, -6.242516e-08, -6.254352e-08, 
    -6.25331e-08, -6.265698e-08, -6.27486e-08, -6.294718e-08, -6.326568e-08, 
    -6.314591e-08, -6.33658e-08, -6.340995e-08, -6.307588e-08, -6.328098e-08, 
    -6.262274e-08, -6.272907e-08, -6.266577e-08, -6.243449e-08, 
    -6.317349e-08, -6.279422e-08, -6.349462e-08, -6.328914e-08, 
    -6.388886e-08, -6.359058e-08, -6.417645e-08, -6.442689e-08, 
    -6.466265e-08, -6.493813e-08, -6.260812e-08, -6.25277e-08, -6.267172e-08, 
    -6.287096e-08, -6.305586e-08, -6.330166e-08, -6.332682e-08, 
    -6.337287e-08, -6.349217e-08, -6.359246e-08, -6.338743e-08, 
    -6.361761e-08, -6.275372e-08, -6.320642e-08, -6.249729e-08, -6.27108e-08, 
    -6.285921e-08, -6.279412e-08, -6.313223e-08, -6.321191e-08, 
    -6.353574e-08, -6.336835e-08, -6.436507e-08, -6.392407e-08, 
    -6.514793e-08, -6.480587e-08, -6.249959e-08, -6.260785e-08, 
    -6.298463e-08, -6.280536e-08, -6.331808e-08, -6.344429e-08, -6.35469e-08, 
    -6.367805e-08, -6.369222e-08, -6.376993e-08, -6.364259e-08, 
    -6.376491e-08, -6.330219e-08, -6.350896e-08, -6.294157e-08, 
    -6.307966e-08, -6.301614e-08, -6.294646e-08, -6.316152e-08, 
    -6.339064e-08, -6.339556e-08, -6.346902e-08, -6.367603e-08, 
    -6.332016e-08, -6.442196e-08, -6.374147e-08, -6.27259e-08, -6.293441e-08, 
    -6.296421e-08, -6.288344e-08, -6.343164e-08, -6.3233e-08, -6.376804e-08, 
    -6.362344e-08, -6.386038e-08, -6.374263e-08, -6.372531e-08, 
    -6.357409e-08, -6.347994e-08, -6.32421e-08, -6.304859e-08, -6.289515e-08, 
    -6.293084e-08, -6.309938e-08, -6.340467e-08, -6.36935e-08, -6.363022e-08, 
    -6.384236e-08, -6.32809e-08, -6.351632e-08, -6.342533e-08, -6.36626e-08, 
    -6.314273e-08, -6.358538e-08, -6.302958e-08, -6.307831e-08, 
    -6.322905e-08, -6.353228e-08, -6.359939e-08, -6.367102e-08, 
    -6.362682e-08, -6.341242e-08, -6.33773e-08, -6.322539e-08, -6.318344e-08, 
    -6.30677e-08, -6.297188e-08, -6.305942e-08, -6.315137e-08, -6.341251e-08, 
    -6.364786e-08, -6.390447e-08, -6.396727e-08, -6.426707e-08, -6.4023e-08, 
    -6.442575e-08, -6.40833e-08, -6.467612e-08, -6.361105e-08, -6.407326e-08, 
    -6.323592e-08, -6.332613e-08, -6.348927e-08, -6.386351e-08, 
    -6.366148e-08, -6.389776e-08, -6.337593e-08, -6.310519e-08, 
    -6.303516e-08, -6.290448e-08, -6.303815e-08, -6.302728e-08, 
    -6.315518e-08, -6.311409e-08, -6.342119e-08, -6.325622e-08, 
    -6.372487e-08, -6.38959e-08, -6.437893e-08, -6.467506e-08, -6.497654e-08, 
    -6.510964e-08, -6.515015e-08, -6.516709e-08 ;

 NET_NMIN =
  8.721912e-09, 8.760372e-09, 8.752895e-09, 8.783916e-09, 8.766709e-09, 
    8.787021e-09, 8.729709e-09, 8.761898e-09, 8.74135e-09, 8.725375e-09, 
    8.844117e-09, 8.7853e-09, 8.905227e-09, 8.86771e-09, 8.96196e-09, 
    8.899388e-09, 8.974578e-09, 8.960157e-09, 9.003568e-09, 8.991131e-09, 
    9.046653e-09, 9.009307e-09, 9.07544e-09, 9.037736e-09, 9.043633e-09, 
    9.008075e-09, 8.797138e-09, 8.836794e-09, 8.794789e-09, 8.800443e-09, 
    8.797906e-09, 8.767064e-09, 8.75152e-09, 8.718974e-09, 8.724882e-09, 
    8.748787e-09, 8.802986e-09, 8.784589e-09, 8.830959e-09, 8.829912e-09, 
    8.881537e-09, 8.85826e-09, 8.945038e-09, 8.920374e-09, 8.99165e-09, 
    8.973724e-09, 8.990808e-09, 8.985627e-09, 8.990875e-09, 8.964585e-09, 
    8.975849e-09, 8.952716e-09, 8.862619e-09, 8.889096e-09, 8.81013e-09, 
    8.762651e-09, 8.731121e-09, 8.708747e-09, 8.711909e-09, 8.717939e-09, 
    8.748928e-09, 8.778065e-09, 8.800272e-09, 8.815125e-09, 8.829762e-09, 
    8.874061e-09, 8.897513e-09, 8.950024e-09, 8.940549e-09, 8.956602e-09, 
    8.971941e-09, 8.997691e-09, 8.993453e-09, 9.004798e-09, 8.95618e-09, 
    8.988491e-09, 8.935151e-09, 8.94974e-09, 8.833734e-09, 8.789552e-09, 
    8.770768e-09, 8.754332e-09, 8.714341e-09, 8.741957e-09, 8.731071e-09, 
    8.756973e-09, 8.773431e-09, 8.765292e-09, 8.815531e-09, 8.795999e-09, 
    8.898903e-09, 8.854577e-09, 8.970152e-09, 8.942494e-09, 8.976781e-09, 
    8.959286e-09, 8.989263e-09, 8.962283e-09, 9.009021e-09, 9.019197e-09, 
    9.012243e-09, 9.03896e-09, 8.960788e-09, 8.990807e-09, 8.765063e-09, 
    8.76639e-09, 8.772576e-09, 8.745387e-09, 8.743724e-09, 8.718811e-09, 
    8.740979e-09, 8.750419e-09, 8.774386e-09, 8.788561e-09, 8.802036e-09, 
    8.831667e-09, 8.864759e-09, 8.911036e-09, 8.944287e-09, 8.966575e-09, 
    8.952909e-09, 8.964975e-09, 8.951486e-09, 8.945165e-09, 9.015384e-09, 
    8.975953e-09, 9.035118e-09, 9.031844e-09, 9.005068e-09, 9.032212e-09, 
    8.767323e-09, 8.759684e-09, 8.733159e-09, 8.753917e-09, 8.716098e-09, 
    8.737266e-09, 8.749438e-09, 8.796405e-09, 8.806727e-09, 8.816295e-09, 
    8.835196e-09, 8.859451e-09, 8.902004e-09, 8.93903e-09, 8.972833e-09, 
    8.970357e-09, 8.971228e-09, 8.978779e-09, 8.960074e-09, 8.98185e-09, 
    8.985505e-09, 8.97595e-09, 9.031405e-09, 9.015562e-09, 9.031774e-09, 
    9.021458e-09, 8.762167e-09, 8.775022e-09, 8.768075e-09, 8.781137e-09, 
    8.771934e-09, 8.812853e-09, 8.825122e-09, 8.882535e-09, 8.858973e-09, 
    8.896474e-09, 8.862783e-09, 8.868752e-09, 8.897694e-09, 8.864604e-09, 
    8.936986e-09, 8.88791e-09, 8.979073e-09, 8.930059e-09, 8.982144e-09, 
    8.972687e-09, 8.988346e-09, 9.00237e-09, 9.020014e-09, 9.052569e-09, 
    9.045031e-09, 9.072258e-09, 8.794186e-09, 8.810859e-09, 8.809392e-09, 
    8.826842e-09, 8.839747e-09, 8.867721e-09, 8.912587e-09, 8.895715e-09, 
    8.92669e-09, 8.932909e-09, 8.88585e-09, 8.914742e-09, 8.822019e-09, 
    8.836997e-09, 8.82808e-09, 8.7955e-09, 8.899601e-09, 8.846174e-09, 
    8.944836e-09, 8.91589e-09, 9.00037e-09, 8.958354e-09, 9.040881e-09, 
    9.076159e-09, 9.10937e-09, 9.148176e-09, 8.81996e-09, 8.808631e-09, 
    8.828918e-09, 8.856984e-09, 8.883029e-09, 8.917656e-09, 8.9212e-09, 
    8.927686e-09, 8.94449e-09, 8.958619e-09, 8.929736e-09, 8.96216e-09, 
    8.840469e-09, 8.90424e-09, 8.804347e-09, 8.834423e-09, 8.85533e-09, 
    8.84616e-09, 8.893788e-09, 8.905013e-09, 8.95063e-09, 8.927048e-09, 
    9.067451e-09, 9.00533e-09, 9.177728e-09, 9.129545e-09, 8.804673e-09, 
    8.819922e-09, 8.872996e-09, 8.847743e-09, 8.919968e-09, 8.937747e-09, 
    8.952201e-09, 8.970676e-09, 8.972671e-09, 8.983618e-09, 8.96568e-09, 
    8.98291e-09, 8.91773e-09, 8.946857e-09, 8.866931e-09, 8.886382e-09, 
    8.877435e-09, 8.867619e-09, 8.897914e-09, 8.93019e-09, 8.930882e-09, 
    8.941231e-09, 8.970392e-09, 8.920261e-09, 9.075465e-09, 8.979608e-09, 
    8.836551e-09, 8.865922e-09, 8.870121e-09, 8.858742e-09, 8.935964e-09, 
    8.907983e-09, 8.983352e-09, 8.962981e-09, 8.996358e-09, 8.979772e-09, 
    8.977332e-09, 8.956031e-09, 8.942769e-09, 8.909265e-09, 8.882006e-09, 
    8.860392e-09, 8.865419e-09, 8.889161e-09, 8.932165e-09, 8.972851e-09, 
    8.963938e-09, 8.993822e-09, 8.914731e-09, 8.947893e-09, 8.935075e-09, 
    8.968499e-09, 8.895267e-09, 8.95762e-09, 8.879328e-09, 8.886193e-09, 
    8.907428e-09, 8.950141e-09, 8.959595e-09, 8.969685e-09, 8.963458e-09, 
    8.933257e-09, 8.928311e-09, 8.906912e-09, 8.901003e-09, 8.884698e-09, 
    8.8712e-09, 8.883533e-09, 8.896484e-09, 8.933271e-09, 8.966422e-09, 
    9.002568e-09, 9.011417e-09, 9.053647e-09, 9.019266e-09, 9.075999e-09, 
    9.027761e-09, 9.111268e-09, 8.961238e-09, 9.026346e-09, 8.908394e-09, 
    8.921101e-09, 8.944083e-09, 8.9968e-09, 8.968342e-09, 9.001624e-09, 
    8.928116e-09, 8.889979e-09, 8.880114e-09, 8.861706e-09, 8.880535e-09, 
    8.879004e-09, 8.897022e-09, 8.891232e-09, 8.934492e-09, 8.911255e-09, 
    8.97727e-09, 9.001362e-09, 9.069405e-09, 9.111118e-09, 9.153586e-09, 
    9.172334e-09, 9.178041e-09, 9.180426e-09 ;

 NFIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NFIX_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 NPP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 OCDEP =
  6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 6.047846e-14, 
    6.047846e-14, 6.047846e-14, 6.047846e-14 ;

 O_SCALAR =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 PARVEGLN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PBOT =
  100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 100154.5, 
    100154.5, 100154.5 ;

 PCH4 =
  0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 0.1702627, 
    0.1702627, 0.1702627 ;

 PCO2 =
  28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 28.51399, 
    28.51399, 28.51399 ;

 PCT_LANDUNIT =
  100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 
    100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PCT_NAT_PFT =
  13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 13.53654, 
    13.53654, 13.53654,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 14.28591, 
    14.28591, 14.28591,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 2.921148, 
    2.921148, 2.921148,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 13.53892, 
    13.53892, 13.53892,
  55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 55.71749, 
    55.71749, 55.71749,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_CTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_FIRE_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PFT_NTRUNC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PLANT_NDEMAND =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 POTENTIAL_IMMOB =
  5.00767e-14, 5.021391e-14, 5.018725e-14, 5.029783e-14, 5.023652e-14, 
    5.03089e-14, 5.010455e-14, 5.021933e-14, 5.014608e-14, 5.008909e-14, 
    5.051216e-14, 5.030277e-14, 5.072961e-14, 5.059623e-14, 5.093115e-14, 
    5.070883e-14, 5.097595e-14, 5.092479e-14, 5.107884e-14, 5.103473e-14, 
    5.123149e-14, 5.10992e-14, 5.133348e-14, 5.119994e-14, 5.122082e-14, 
    5.109482e-14, 5.034498e-14, 5.048609e-14, 5.03366e-14, 5.035673e-14, 
    5.034771e-14, 5.023776e-14, 5.01823e-14, 5.006624e-14, 5.008733e-14, 
    5.017259e-14, 5.036579e-14, 5.030026e-14, 5.046545e-14, 5.046172e-14, 
    5.064542e-14, 5.056262e-14, 5.08711e-14, 5.07835e-14, 5.103657e-14, 
    5.097296e-14, 5.103357e-14, 5.10152e-14, 5.103381e-14, 5.094051e-14, 
    5.098049e-14, 5.089838e-14, 5.057812e-14, 5.067229e-14, 5.039125e-14, 
    5.022198e-14, 5.010957e-14, 5.002974e-14, 5.004103e-14, 5.006253e-14, 
    5.017309e-14, 5.027701e-14, 5.035615e-14, 5.040906e-14, 5.046119e-14, 
    5.061875e-14, 5.070219e-14, 5.088879e-14, 5.085517e-14, 5.091215e-14, 
    5.096663e-14, 5.105799e-14, 5.104296e-14, 5.108319e-14, 5.091068e-14, 
    5.102534e-14, 5.083601e-14, 5.088781e-14, 5.047519e-14, 5.031795e-14, 
    5.025093e-14, 5.019237e-14, 5.00497e-14, 5.014823e-14, 5.010939e-14, 
    5.020181e-14, 5.026049e-14, 5.023147e-14, 5.041051e-14, 5.034092e-14, 
    5.070713e-14, 5.054949e-14, 5.096027e-14, 5.086208e-14, 5.098381e-14, 
    5.092171e-14, 5.102808e-14, 5.093235e-14, 5.109817e-14, 5.113424e-14, 
    5.110959e-14, 5.12043e-14, 5.092704e-14, 5.103356e-14, 5.023065e-14, 
    5.023538e-14, 5.025744e-14, 5.016046e-14, 5.015453e-14, 5.006566e-14, 
    5.014476e-14, 5.017841e-14, 5.02639e-14, 5.031441e-14, 5.036243e-14, 
    5.046796e-14, 5.058571e-14, 5.075028e-14, 5.086844e-14, 5.094759e-14, 
    5.089907e-14, 5.094191e-14, 5.089402e-14, 5.087157e-14, 5.112071e-14, 
    5.098085e-14, 5.119068e-14, 5.117909e-14, 5.108414e-14, 5.118039e-14, 
    5.023871e-14, 5.021148e-14, 5.011685e-14, 5.019091e-14, 5.005598e-14, 
    5.01315e-14, 5.017489e-14, 5.034234e-14, 5.037914e-14, 5.041322e-14, 
    5.048053e-14, 5.056685e-14, 5.071818e-14, 5.084976e-14, 5.09698e-14, 
    5.096101e-14, 5.096411e-14, 5.09909e-14, 5.092451e-14, 5.100179e-14, 
    5.101474e-14, 5.098085e-14, 5.117753e-14, 5.112137e-14, 5.117884e-14, 
    5.114228e-14, 5.022034e-14, 5.026616e-14, 5.024139e-14, 5.028795e-14, 
    5.025514e-14, 5.040092e-14, 5.044461e-14, 5.064893e-14, 5.056515e-14, 
    5.069851e-14, 5.057871e-14, 5.059994e-14, 5.070279e-14, 5.05852e-14, 
    5.084247e-14, 5.066803e-14, 5.099194e-14, 5.081783e-14, 5.100284e-14, 
    5.096928e-14, 5.102485e-14, 5.107458e-14, 5.113715e-14, 5.125249e-14, 
    5.12258e-14, 5.132223e-14, 5.033446e-14, 5.039384e-14, 5.038864e-14, 
    5.045079e-14, 5.049672e-14, 5.059628e-14, 5.075581e-14, 5.069585e-14, 
    5.080595e-14, 5.082803e-14, 5.066078e-14, 5.076346e-14, 5.043359e-14, 
    5.048689e-14, 5.045518e-14, 5.033913e-14, 5.070963e-14, 5.051957e-14, 
    5.087039e-14, 5.076756e-14, 5.106749e-14, 5.091836e-14, 5.12111e-14, 
    5.133598e-14, 5.145358e-14, 5.159071e-14, 5.042627e-14, 5.038593e-14, 
    5.045818e-14, 5.055804e-14, 5.065073e-14, 5.077382e-14, 5.078643e-14, 
    5.080947e-14, 5.086918e-14, 5.091934e-14, 5.081673e-14, 5.093192e-14, 
    5.049919e-14, 5.072613e-14, 5.037065e-14, 5.047773e-14, 5.055217e-14, 
    5.051955e-14, 5.0689e-14, 5.07289e-14, 5.089095e-14, 5.080722e-14, 
    5.130514e-14, 5.108504e-14, 5.169514e-14, 5.152488e-14, 5.037183e-14, 
    5.042615e-14, 5.061502e-14, 5.052519e-14, 5.078206e-14, 5.084521e-14, 
    5.089656e-14, 5.096212e-14, 5.096922e-14, 5.100806e-14, 5.094441e-14, 
    5.100556e-14, 5.077409e-14, 5.087757e-14, 5.059348e-14, 5.066265e-14, 
    5.063085e-14, 5.059593e-14, 5.070367e-14, 5.081833e-14, 5.082084e-14, 
    5.085757e-14, 5.096097e-14, 5.07831e-14, 5.133343e-14, 5.09937e-14, 
    5.048536e-14, 5.058984e-14, 5.060481e-14, 5.056434e-14, 5.083888e-14, 
    5.073945e-14, 5.100712e-14, 5.093483e-14, 5.105327e-14, 5.099442e-14, 
    5.098576e-14, 5.091016e-14, 5.086305e-14, 5.0744e-14, 5.064708e-14, 
    5.057022e-14, 5.05881e-14, 5.067253e-14, 5.082536e-14, 5.096984e-14, 
    5.09382e-14, 5.104427e-14, 5.076344e-14, 5.088123e-14, 5.08357e-14, 
    5.095441e-14, 5.069424e-14, 5.091566e-14, 5.063758e-14, 5.066199e-14, 
    5.073748e-14, 5.088918e-14, 5.092281e-14, 5.09586e-14, 5.093653e-14, 
    5.082924e-14, 5.081168e-14, 5.073565e-14, 5.071463e-14, 5.065668e-14, 
    5.060867e-14, 5.065253e-14, 5.069856e-14, 5.082931e-14, 5.094702e-14, 
    5.107528e-14, 5.110667e-14, 5.125624e-14, 5.113442e-14, 5.133531e-14, 
    5.116443e-14, 5.146017e-14, 5.092856e-14, 5.115951e-14, 5.074093e-14, 
    5.078609e-14, 5.086768e-14, 5.105478e-14, 5.095385e-14, 5.10719e-14, 
    5.0811e-14, 5.067541e-14, 5.064038e-14, 5.057488e-14, 5.064187e-14, 
    5.063643e-14, 5.07005e-14, 5.067992e-14, 5.083365e-14, 5.075109e-14, 
    5.098553e-14, 5.107098e-14, 5.131211e-14, 5.145971e-14, 5.160989e-14, 
    5.167611e-14, 5.169627e-14, 5.170469e-14 ;

 POT_F_DENIT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.605194e-45, 0, 4.551417e-42, 
    2.802597e-45, 1.913193e-41, 3.698027e-42, 4.768479e-40, 1.216804e-40, 
    4.618803e-38, 8.893803e-40, 8.562508e-37, 1.82806e-38, 3.377825e-38, 
    7.783162e-40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.403934e-43, 3.363116e-44, 1.288718e-40, 1.736209e-41, 1.174148e-40, 
    6.60418e-41, 1.182948e-40, 6.143292e-42, 2.207185e-41, 1.56525e-42, 0, 
    1.401298e-45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 
    1.146262e-42, 3.783506e-43, 2.455075e-42, 1.418815e-41, 2.508002e-40, 
    1.572887e-40, 5.453685e-40, 2.337366e-42, 9.083777e-41, 1.989844e-43, 
    1.108427e-42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.802597e-45, 0, 
    1.158313e-41, 4.750402e-43, 2.451432e-41, 3.343498e-42, 9.89597e-41, 
    4.718172e-42, 8.623619e-40, 2.577666e-39, 1.221582e-39, 2.076547e-38, 
    3.974082e-42, 1.174288e-40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.121039e-44, 5.857428e-43, 7.708543e-42, 1.600283e-42, 6.42075e-42, 
    1.356457e-42, 6.488012e-43, 1.713117e-39, 2.23367e-41, 1.389566e-38, 
    9.852799e-39, 5.616474e-40, 1.024267e-38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4.203895e-45, 3.152922e-43, 1.569594e-41, 1.185358e-41, 
    1.308673e-41, 3.069544e-41, 3.661593e-42, 4.331554e-41, 6.516038e-41, 
    2.232128e-41, 9.408437e-39, 1.745448e-39, 9.780899e-39, 3.279918e-39, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1.401298e-45, 0, 0, 2.802597e-45, 0, 
    2.480298e-43, 0, 3.1724e-41, 1.093013e-43, 4.476448e-41, 1.543811e-41, 
    8.93538e-41, 4.185454e-40, 2.811773e-39, 8.485865e-38, 3.902624e-38, 
    6.231172e-37, 0, 0, 0, 0, 0, 0, 1.261169e-44, 1.401298e-45, 7.286752e-44, 
    1.527415e-43, 0, 1.681558e-44, 0, 0, 0, 0, 2.802597e-45, 0, 6.249791e-43, 
    1.961818e-44, 3.363915e-40, 3.005785e-42, 2.536987e-38, 9.203849e-37, 
    2.340174e-35, 8.675964e-34, 0, 0, 0, 0, 0, 2.522337e-44, 3.783506e-44, 
    8.267661e-44, 5.997557e-43, 3.09687e-42, 1.050974e-43, 4.652311e-42, 0, 
    4.203895e-45, 0, 0, 0, 0, 1.401298e-45, 5.605194e-45, 1.228939e-42, 
    7.567012e-44, 3.850611e-37, 5.781982e-40, 1.20543e-32, 1.566253e-34, 0, 
    0, 0, 0, 3.222986e-44, 2.718519e-43, 1.474166e-42, 1.229499e-41, 
    1.541148e-41, 5.278831e-41, 6.960249e-42, 4.876519e-41, 2.522337e-44, 
    7.917336e-43, 0, 0, 0, 0, 2.802597e-45, 1.107026e-43, 1.205117e-43, 
    4.091792e-43, 1.193206e-41, 3.363116e-44, 8.600233e-37, 3.375868e-41, 0, 
    0, 0, 0, 2.200039e-43, 7.006492e-45, 5.123568e-41, 5.111937e-42, 
    2.165973e-40, 3.4315e-41, 2.608517e-41, 2.298129e-42, 4.904545e-43, 
    8.407791e-45, 0, 0, 0, 1.401298e-45, 1.401298e-43, 1.573378e-41, 
    5.706087e-42, 1.638048e-40, 1.681558e-44, 8.940284e-43, 1.975831e-43, 
    9.598894e-42, 1.401298e-45, 2.766163e-42, 0, 0, 7.006492e-45, 
    1.161676e-42, 3.465411e-42, 1.098618e-41, 5.399203e-42, 1.59748e-43, 
    8.82818e-44, 7.006492e-45, 2.802597e-45, 0, 0, 0, 1.401298e-45, 
    1.59748e-43, 7.578222e-42, 4.277912e-40, 1.117072e-39, 9.486179e-38, 
    2.598732e-39, 9.070593e-37, 6.421963e-39, 2.808711e-35, 4.191284e-42, 
    5.521899e-39, 8.407791e-45, 3.783506e-44, 5.717298e-43, 2.275709e-40, 
    9.427936e-42, 3.860339e-40, 8.68805e-44, 1.401298e-45, 0, 0, 0, 0, 
    1.401298e-45, 1.401298e-45, 1.849714e-43, 1.121039e-44, 2.590861e-41, 
    3.750631e-40, 4.682267e-37, 2.766208e-35, 1.414291e-33, 7.510774e-33, 
    1.238513e-32, 1.524886e-32 ;

 POT_F_NIT =
  3.831289e-11, 3.864309e-11, 3.857878e-11, 3.884595e-11, 3.869762e-11, 
    3.887273e-11, 3.83797e-11, 3.865619e-11, 3.847956e-11, 3.834253e-11, 
    3.936713e-11, 3.885786e-11, 3.98999e-11, 3.957237e-11, 4.039783e-11, 
    3.984882e-11, 4.050901e-11, 4.038195e-11, 4.076504e-11, 4.065509e-11, 
    4.114711e-11, 4.081582e-11, 4.140342e-11, 4.106787e-11, 4.112025e-11, 
    4.080489e-11, 3.896012e-11, 3.930356e-11, 3.89398e-11, 3.898867e-11, 
    3.896674e-11, 3.870066e-11, 3.856692e-11, 3.828768e-11, 3.833829e-11, 
    3.854343e-11, 3.901062e-11, 3.88517e-11, 3.925288e-11, 3.92438e-11, 
    3.96929e-11, 3.949007e-11, 4.024895e-11, 4.003249e-11, 4.065967e-11, 
    4.050145e-11, 4.065222e-11, 4.060646e-11, 4.06528e-11, 4.04209e-11, 
    4.052016e-11, 4.031641e-11, 3.952807e-11, 3.975893e-11, 3.907245e-11, 
    3.866267e-11, 3.839178e-11, 3.820015e-11, 3.822721e-11, 3.827882e-11, 
    3.854463e-11, 3.879543e-11, 3.898714e-11, 3.911564e-11, 3.924248e-11, 
    3.962769e-11, 3.983241e-11, 4.029277e-11, 4.02095e-11, 4.035063e-11, 
    4.048572e-11, 4.071304e-11, 4.067558e-11, 4.077588e-11, 4.034689e-11, 
    4.063172e-11, 4.016206e-11, 4.029023e-11, 3.927698e-11, 3.889456e-11, 
    3.873256e-11, 3.859109e-11, 3.824802e-11, 3.848476e-11, 3.839133e-11, 
    3.861378e-11, 3.875547e-11, 3.868536e-11, 3.911915e-11, 3.895019e-11, 
    3.984455e-11, 3.945801e-11, 4.046996e-11, 4.022658e-11, 4.052839e-11, 
    4.037424e-11, 4.063855e-11, 4.040062e-11, 4.081325e-11, 4.090338e-11, 
    4.084176e-11, 4.107871e-11, 4.038742e-11, 4.065216e-11, 3.868342e-11, 
    3.869485e-11, 3.874812e-11, 3.85142e-11, 3.849992e-11, 3.828626e-11, 
    3.847634e-11, 3.855742e-11, 3.876369e-11, 3.888595e-11, 3.900237e-11, 
    3.925899e-11, 3.954662e-11, 3.995068e-11, 4.024232e-11, 4.043842e-11, 
    4.031812e-11, 4.042431e-11, 4.030559e-11, 4.025001e-11, 4.086958e-11, 
    4.052106e-11, 4.104457e-11, 4.101551e-11, 4.077823e-11, 4.101878e-11, 
    3.870287e-11, 3.86371e-11, 3.840923e-11, 3.858749e-11, 3.826303e-11, 
    3.844446e-11, 3.854898e-11, 3.89537e-11, 3.904293e-11, 3.912575e-11, 
    3.92896e-11, 3.95004e-11, 3.987164e-11, 4.019613e-11, 4.049357e-11, 
    4.047173e-11, 4.047941e-11, 4.054599e-11, 4.038115e-11, 4.057308e-11, 
    4.060533e-11, 4.052102e-11, 4.101161e-11, 4.087113e-11, 4.101488e-11, 
    4.092338e-11, 3.865847e-11, 3.876918e-11, 3.870932e-11, 3.88219e-11, 
    3.874255e-11, 3.909595e-11, 3.920223e-11, 3.970157e-11, 3.949625e-11, 
    3.98233e-11, 3.95294e-11, 3.958139e-11, 3.983395e-11, 3.954524e-11, 
    4.017817e-11, 3.974846e-11, 4.054857e-11, 4.011736e-11, 4.057567e-11, 
    4.049224e-11, 4.063041e-11, 4.075435e-11, 4.091057e-11, 4.119964e-11, 
    4.11326e-11, 4.137497e-11, 3.893453e-11, 3.907869e-11, 3.9066e-11, 
    3.921714e-11, 3.932911e-11, 3.957241e-11, 3.996426e-11, 3.981666e-11, 
    4.008784e-11, 4.014239e-11, 3.973049e-11, 3.998311e-11, 3.917529e-11, 
    3.93052e-11, 3.922783e-11, 3.894582e-11, 3.985059e-11, 3.938488e-11, 
    4.024709e-11, 3.999313e-11, 4.073665e-11, 4.036597e-11, 4.109572e-11, 
    4.140975e-11, 4.17065e-11, 4.205463e-11, 3.91575e-11, 3.90594e-11, 
    3.923513e-11, 3.947893e-11, 3.970588e-11, 4.000865e-11, 4.003969e-11, 
    4.009656e-11, 4.024408e-11, 4.036834e-11, 4.011453e-11, 4.039951e-11, 
    3.933533e-11, 3.989115e-11, 3.902227e-11, 3.928284e-11, 3.946448e-11, 
    3.938476e-11, 3.979976e-11, 3.989789e-11, 4.029799e-11, 4.009091e-11, 
    4.13321e-11, 4.078051e-11, 4.232075e-11, 4.188729e-11, 3.902515e-11, 
    3.915714e-11, 3.961837e-11, 3.939856e-11, 4.002889e-11, 4.018485e-11, 
    4.031187e-11, 4.047454e-11, 4.049212e-11, 4.058868e-11, 4.04305e-11, 
    4.058242e-11, 4.000924e-11, 4.026485e-11, 3.956547e-11, 3.973508e-11, 
    3.9657e-11, 3.957144e-11, 3.98358e-11, 4.011846e-11, 4.012453e-11, 
    4.021538e-11, 4.047196e-11, 4.003137e-11, 4.140353e-11, 4.055322e-11, 
    3.930135e-11, 3.955673e-11, 3.959329e-11, 3.949421e-11, 4.016919e-11, 
    3.992392e-11, 4.058633e-11, 4.040673e-11, 4.07012e-11, 4.055473e-11, 
    4.053319e-11, 4.034554e-11, 4.022892e-11, 3.993511e-11, 3.969688e-11, 
    3.950852e-11, 3.955227e-11, 3.975932e-11, 4.013578e-11, 4.049364e-11, 
    4.04151e-11, 4.067872e-11, 3.998292e-11, 4.027391e-11, 4.016129e-11, 
    4.045525e-11, 3.981272e-11, 4.035956e-11, 3.967356e-11, 3.973346e-11, 
    3.991905e-11, 4.029374e-11, 4.03769e-11, 4.046577e-11, 4.041092e-11, 
    4.01454e-11, 4.010198e-11, 3.99145e-11, 3.986281e-11, 3.972037e-11, 
    3.960263e-11, 3.971019e-11, 3.982329e-11, 4.014548e-11, 4.043698e-11, 
    4.075606e-11, 4.083435e-11, 4.120916e-11, 4.090388e-11, 4.140826e-11, 
    4.09792e-11, 4.172343e-11, 4.039138e-11, 4.096674e-11, 3.992751e-11, 
    4.003879e-11, 4.024048e-11, 4.070509e-11, 4.045392e-11, 4.074775e-11, 
    4.010028e-11, 3.976648e-11, 3.968037e-11, 3.951995e-11, 3.968403e-11, 
    3.967067e-11, 3.982799e-11, 3.977739e-11, 4.015618e-11, 3.995248e-11, 
    4.053259e-11, 4.074538e-11, 4.134947e-11, 4.172209e-11, 4.210324e-11, 
    4.227207e-11, 4.232353e-11, 4.234505e-11 ;

 PROD100C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD100N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10C_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PROD10N_LOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_CLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PRODUCT_NLOSS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHA =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSHADE_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 PSNSUN_TO_CPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Q2M =
  0.0005857516, 0.0005857558, 0.000585755, 0.0005857584, 0.0005857565, 
    0.0005857587, 0.0005857525, 0.0005857559, 0.0005857538, 0.000585752, 
    0.0005857648, 0.0005857585, 0.0005857716, 0.0005857676, 0.0005857779, 
    0.0005857709, 0.0005857793, 0.0005857777, 0.0005857826, 0.0005857812, 
    0.0005857872, 0.0005857832, 0.0005857904, 0.0005857863, 0.0005857869, 
    0.000585783, 0.0005857599, 0.0005857639, 0.0005857596, 0.0005857602, 
    0.0005857599, 0.0005857566, 0.0005857548, 0.0005857513, 0.000585752, 
    0.0005857545, 0.0005857605, 0.0005857585, 0.0005857636, 0.0005857635, 
    0.0005857691, 0.0005857665, 0.0005857761, 0.0005857734, 0.0005857812, 
    0.0005857793, 0.0005857811, 0.0005857806, 0.0005857811, 0.0005857782, 
    0.0005857795, 0.0005857769, 0.000585767, 0.0005857699, 0.0005857613, 
    0.0005857559, 0.0005857526, 0.0005857502, 0.0005857506, 0.0005857512, 
    0.0005857545, 0.0005857578, 0.0005857602, 0.0005857619, 0.0005857634, 
    0.0005857681, 0.0005857708, 0.0005857766, 0.0005857756, 0.0005857773, 
    0.000585779, 0.0005857819, 0.0005857814, 0.0005857827, 0.0005857773, 
    0.0005857808, 0.000585775, 0.0005857766, 0.0005857636, 0.000585759, 
    0.0005857568, 0.0005857552, 0.0005857508, 0.0005857538, 0.0005857526, 
    0.0005857554, 0.0005857573, 0.0005857564, 0.0005857619, 0.0005857598, 
    0.0005857709, 0.0005857661, 0.0005857788, 0.0005857758, 0.0005857796, 
    0.0005857777, 0.0005857809, 0.000585778, 0.0005857832, 0.0005857843, 
    0.0005857835, 0.0005857865, 0.0005857778, 0.0005857811, 0.0005857563, 
    0.0005857565, 0.0005857572, 0.0005857542, 0.000585754, 0.0005857513, 
    0.0005857537, 0.0005857547, 0.0005857574, 0.0005857589, 0.0005857604, 
    0.0005857636, 0.0005857672, 0.0005857723, 0.000585776, 0.0005857784, 
    0.000585777, 0.0005857783, 0.0005857768, 0.0005857761, 0.0005857838, 
    0.0005857794, 0.0005857861, 0.0005857857, 0.0005857827, 0.0005857857, 
    0.0005857566, 0.0005857558, 0.0005857528, 0.0005857552, 0.000585751, 
    0.0005857533, 0.0005857546, 0.0005857597, 0.0005857609, 0.0005857619, 
    0.000585764, 0.0005857667, 0.0005857713, 0.0005857754, 0.0005857791, 
    0.0005857789, 0.000585779, 0.0005857798, 0.0005857777, 0.0005857801, 
    0.0005857805, 0.0005857795, 0.0005857857, 0.0005857839, 0.0005857857, 
    0.0005857846, 0.000585756, 0.0005857574, 0.0005857567, 0.0005857581, 
    0.0005857571, 0.0005857615, 0.0005857628, 0.0005857691, 0.0005857666, 
    0.0005857707, 0.000585767, 0.0005857677, 0.0005857707, 0.0005857673, 
    0.0005857751, 0.0005857697, 0.0005857798, 0.0005857743, 0.0005857802, 
    0.0005857791, 0.0005857809, 0.0005857824, 0.0005857844, 0.0005857879, 
    0.0005857871, 0.0005857901, 0.0005857595, 0.0005857613, 0.0005857612, 
    0.0005857631, 0.0005857645, 0.0005857676, 0.0005857725, 0.0005857706, 
    0.0005857741, 0.0005857747, 0.0005857696, 0.0005857727, 0.0005857626, 
    0.0005857641, 0.0005857632, 0.0005857596, 0.000585771, 0.0005857651, 
    0.0005857761, 0.0005857729, 0.0005857822, 0.0005857775, 0.0005857866, 
    0.0005857905, 0.0005857943, 0.0005857985, 0.0005857623, 0.0005857612, 
    0.0005857634, 0.0005857663, 0.0005857692, 0.000585773, 0.0005857734, 
    0.0005857741, 0.0005857761, 0.0005857776, 0.0005857743, 0.000585778, 
    0.0005857644, 0.0005857715, 0.0005857606, 0.0005857638, 0.0005857662, 
    0.0005857652, 0.0005857705, 0.0005857717, 0.0005857766, 0.0005857741, 
    0.0005857895, 0.0005857826, 0.0005858019, 0.0005857965, 0.0005857607, 
    0.0005857624, 0.0005857681, 0.0005857654, 0.0005857733, 0.0005857752, 
    0.0005857769, 0.0005857789, 0.0005857791, 0.0005857803, 0.0005857784, 
    0.0005857802, 0.000585773, 0.0005857763, 0.0005857675, 0.0005857696, 
    0.0005857687, 0.0005857676, 0.0005857709, 0.0005857744, 0.0005857745, 
    0.0005857756, 0.0005857786, 0.0005857734, 0.0005857902, 0.0005857796, 
    0.0005857642, 0.0005857673, 0.0005857678, 0.0005857666, 0.0005857751, 
    0.000585772, 0.0005857803, 0.0005857781, 0.0005857818, 0.0005857799, 
    0.0005857797, 0.0005857773, 0.0005857758, 0.0005857721, 0.0005857691, 
    0.0005857668, 0.0005857673, 0.0005857699, 0.0005857746, 0.0005857791, 
    0.0005857781, 0.0005857815, 0.0005857727, 0.0005857763, 0.0005857749, 
    0.0005857787, 0.0005857706, 0.0005857772, 0.0005857689, 0.0005857696, 
    0.0005857719, 0.0005857765, 0.0005857777, 0.0005857788, 0.0005857782, 
    0.0005857747, 0.0005857742, 0.0005857719, 0.0005857712, 0.0005857695, 
    0.000585768, 0.0005857693, 0.0005857707, 0.0005857748, 0.0005857784, 
    0.0005857824, 0.0005857834, 0.0005857879, 0.0005857841, 0.0005857903, 
    0.0005857849, 0.0005857943, 0.0005857777, 0.0005857849, 0.000585772, 
    0.0005857734, 0.0005857759, 0.0005857817, 0.0005857787, 0.0005857822, 
    0.0005857742, 0.0005857699, 0.000585769, 0.0005857669, 0.000585769, 
    0.0005857688, 0.0005857708, 0.0005857702, 0.0005857749, 0.0005857724, 
    0.0005857796, 0.0005857822, 0.0005857898, 0.0005857944, 0.0005857992, 
    0.0005858013, 0.000585802, 0.0005858022 ;

 QBOT =
  0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 0.0005799045, 
    0.0005799045, 0.0005799045, 0.0005799045 ;

 QCHARGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_PERCH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRAI_XS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QDRIP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLOOD =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_ICE_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QFLX_LIQ_DYNBAL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QH2OSFC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QINFL =
  -2.651793e-07, -2.653274e-07, -2.65299e-07, -2.654173e-07, -2.653522e-07, 
    -2.654292e-07, -2.6521e-07, -2.653327e-07, -2.652548e-07, -2.651935e-07, 
    -2.65644e-07, -2.654227e-07, -2.658788e-07, -2.657376e-07, -2.660931e-07, 
    -2.65856e-07, -2.66141e-07, -2.660877e-07, -2.662513e-07, -2.662046e-07, 
    -2.664099e-07, -2.662728e-07, -2.665182e-07, -2.66378e-07, -2.663994e-07, 
    -2.66268e-07, -2.654687e-07, -2.65616e-07, -2.654596e-07, -2.654808e-07, 
    -2.654716e-07, -2.653531e-07, -2.652922e-07, -2.651689e-07, 
    -2.651916e-07, -2.652827e-07, -2.654903e-07, -2.654209e-07, 
    -2.655983e-07, -2.655944e-07, -2.657902e-07, -2.65702e-07, -2.660307e-07, 
    -2.659379e-07, -2.662066e-07, -2.66139e-07, -2.662032e-07, -2.661839e-07, 
    -2.662034e-07, -2.661043e-07, -2.661467e-07, -2.660599e-07, 
    -2.657183e-07, -2.658186e-07, -2.65518e-07, -2.653342e-07, -2.652151e-07, 
    -2.651293e-07, -2.651415e-07, -2.651643e-07, -2.652832e-07, 
    -2.653959e-07, -2.654811e-07, -2.655378e-07, -2.655938e-07, 
    -2.657592e-07, -2.658495e-07, -2.660487e-07, -2.660141e-07, 
    -2.660737e-07, -2.661323e-07, -2.662289e-07, -2.662132e-07, 
    -2.662553e-07, -2.66073e-07, -2.661938e-07, -2.659941e-07, -2.660487e-07, 
    -2.656041e-07, -2.654399e-07, -2.653656e-07, -2.653042e-07, 
    -2.651507e-07, -2.652565e-07, -2.652147e-07, -2.653152e-07, 
    -2.653781e-07, -2.653472e-07, -2.655394e-07, -2.654646e-07, 
    -2.658549e-07, -2.656872e-07, -2.661255e-07, -2.660213e-07, 
    -2.661506e-07, -2.660849e-07, -2.66197e-07, -2.660962e-07, -2.662714e-07, 
    -2.663089e-07, -2.662831e-07, -2.663835e-07, -2.660904e-07, 
    -2.662027e-07, -2.653461e-07, -2.653511e-07, -2.65375e-07, -2.652696e-07, 
    -2.652635e-07, -2.651681e-07, -2.652534e-07, -2.652893e-07, 
    -2.653821e-07, -2.65436e-07, -2.654875e-07, -2.656006e-07, -2.657257e-07, 
    -2.659015e-07, -2.66028e-07, -2.661124e-07, -2.66061e-07, -2.661063e-07, 
    -2.660555e-07, -2.660318e-07, -2.662945e-07, -2.661468e-07, 
    -2.663691e-07, -2.66357e-07, -2.662561e-07, -2.663583e-07, -2.653547e-07, 
    -2.653257e-07, -2.652232e-07, -2.653034e-07, -2.651577e-07, 
    -2.652387e-07, -2.652849e-07, -2.654651e-07, -2.655057e-07, 
    -2.655418e-07, -2.656143e-07, -2.657065e-07, -2.658675e-07, 
    -2.660077e-07, -2.661359e-07, -2.661266e-07, -2.661299e-07, 
    -2.661579e-07, -2.660877e-07, -2.661695e-07, -2.661828e-07, 
    -2.661474e-07, -2.663553e-07, -2.662961e-07, -2.663567e-07, 
    -2.663183e-07, -2.653352e-07, -2.653843e-07, -2.653577e-07, 
    -2.654074e-07, -2.65372e-07, -2.655276e-07, -2.655741e-07, -2.657928e-07, 
    -2.657044e-07, -2.658463e-07, -2.657193e-07, -2.657415e-07, 
    -2.658488e-07, -2.657265e-07, -2.65999e-07, -2.658126e-07, -2.66159e-07, 
    -2.659717e-07, -2.661706e-07, -2.661354e-07, -2.661942e-07, 
    -2.662463e-07, -2.663127e-07, -2.664333e-07, -2.664056e-07, 
    -2.665071e-07, -2.654577e-07, -2.655206e-07, -2.65516e-07, -2.655824e-07, 
    -2.656313e-07, -2.657382e-07, -2.65908e-07, -2.658445e-07, -2.659619e-07, 
    -2.659851e-07, -2.658073e-07, -2.659157e-07, -2.655634e-07, 
    -2.656195e-07, -2.655868e-07, -2.654621e-07, -2.658579e-07, 
    -2.656546e-07, -2.660299e-07, -2.659207e-07, -2.662388e-07, -2.6608e-07, 
    -2.663901e-07, -2.665195e-07, -2.666451e-07, -2.667863e-07, 
    -2.655559e-07, -2.655131e-07, -2.655906e-07, -2.656959e-07, -2.65796e-07, 
    -2.659272e-07, -2.659411e-07, -2.659653e-07, -2.660292e-07, 
    -2.660823e-07, -2.659721e-07, -2.660958e-07, -2.656307e-07, 
    -2.658759e-07, -2.654961e-07, -2.656095e-07, -2.656901e-07, 
    -2.656557e-07, -2.658375e-07, -2.658799e-07, -2.660513e-07, 
    -2.659633e-07, -2.664868e-07, -2.66256e-07, -2.668965e-07, -2.667181e-07, 
    -2.654979e-07, -2.655562e-07, -2.657573e-07, -2.656619e-07, 
    -2.659364e-07, -2.660033e-07, -2.660583e-07, -2.66127e-07, -2.661351e-07, 
    -2.661759e-07, -2.66109e-07, -2.661737e-07, -2.659275e-07, -2.660378e-07, 
    -2.657355e-07, -2.658088e-07, -2.657754e-07, -2.65738e-07, -2.65853e-07, 
    -2.659736e-07, -2.659777e-07, -2.66016e-07, -2.66121e-07, -2.659376e-07, 
    -2.665137e-07, -2.661564e-07, -2.656196e-07, -2.657296e-07, 
    -2.657471e-07, -2.657042e-07, -2.659965e-07, -2.658907e-07, 
    -2.661752e-07, -2.660988e-07, -2.662242e-07, -2.661618e-07, 
    -2.661526e-07, -2.660726e-07, -2.660223e-07, -2.658953e-07, -2.65792e-07, 
    -2.657106e-07, -2.657297e-07, -2.65819e-07, -2.659813e-07, -2.661352e-07, 
    -2.661014e-07, -2.662147e-07, -2.659165e-07, -2.660411e-07, 
    -2.659925e-07, -2.661193e-07, -2.658425e-07, -2.660738e-07, 
    -2.657826e-07, -2.658086e-07, -2.658886e-07, -2.660485e-07, -2.66086e-07, 
    -2.661233e-07, -2.661006e-07, -2.659857e-07, -2.659675e-07, -2.65887e-07, 
    -2.65864e-07, -2.65803e-07, -2.657517e-07, -2.657982e-07, -2.658467e-07, 
    -2.659864e-07, -2.66111e-07, -2.662468e-07, -2.662806e-07, -2.664348e-07, 
    -2.663073e-07, -2.665154e-07, -2.663354e-07, -2.666479e-07, 
    -2.660894e-07, -2.663332e-07, -2.658928e-07, -2.659408e-07, -2.66026e-07, 
    -2.662238e-07, -2.661187e-07, -2.662423e-07, -2.659669e-07, 
    -2.658214e-07, -2.657855e-07, -2.657153e-07, -2.657871e-07, 
    -2.657813e-07, -2.658497e-07, -2.658279e-07, -2.65991e-07, -2.659035e-07, 
    -2.661519e-07, -2.662417e-07, -2.664959e-07, -2.666499e-07, 
    -2.668083e-07, -2.668773e-07, -2.668984e-07, -2.669071e-07 ;

 QINTR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QIRRIG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QOVER_LAG =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRGWL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF_R =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QRUNOFF_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 QSNOMELT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSNWCPICE_NODYNLNDUSE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QSOIL =
  8.802504e-06, 8.828126e-06, 8.823152e-06, 8.843814e-06, 8.832363e-06, 
    8.845886e-06, 8.807713e-06, 8.82913e-06, 8.815465e-06, 8.804832e-06, 
    8.883915e-06, 8.84474e-06, 8.924839e-06, 8.899776e-06, 8.962832e-06, 
    8.920915e-06, 8.971299e-06, 8.96166e-06, 8.990775e-06, 8.982433e-06, 
    9.019629e-06, 8.994627e-06, 9.038992e-06, 9.013676e-06, 9.017621e-06, 
    8.993797e-06, 8.852654e-06, 8.879021e-06, 8.851084e-06, 8.854844e-06, 
    8.853165e-06, 8.832587e-06, 8.8222e-06, 8.800572e-06, 8.804504e-06, 
    8.820403e-06, 8.856536e-06, 8.844288e-06, 8.875239e-06, 8.87454e-06, 
    8.909024e-06, 8.893469e-06, 8.95153e-06, 8.935023e-06, 8.982783e-06, 
    8.970757e-06, 8.982211e-06, 8.978743e-06, 8.982256e-06, 8.964625e-06, 
    8.972175e-06, 8.956678e-06, 8.896375e-06, 8.914071e-06, 8.861314e-06, 
    8.829596e-06, 8.808645e-06, 8.793761e-06, 8.795864e-06, 8.799868e-06, 
    8.820496e-06, 8.839938e-06, 8.854755e-06, 8.864665e-06, 8.874439e-06, 
    8.903958e-06, 8.919677e-06, 8.95485e-06, 8.948531e-06, 8.959261e-06, 
    8.969563e-06, 8.986824e-06, 8.983987e-06, 8.991587e-06, 8.959002e-06, 
    8.980642e-06, 8.944925e-06, 8.954685e-06, 8.87697e-06, 8.847598e-06, 
    8.835016e-06, 8.824103e-06, 8.797479e-06, 8.815855e-06, 8.808607e-06, 
    8.825881e-06, 8.836847e-06, 8.831428e-06, 8.864936e-06, 8.851899e-06, 
    8.92061e-06, 8.890989e-06, 8.968362e-06, 8.949831e-06, 8.97281e-06, 
    8.961088e-06, 8.981166e-06, 8.963096e-06, 8.994426e-06, 9.001238e-06, 
    8.99658e-06, 9.014522e-06, 8.962091e-06, 8.982199e-06, 8.831271e-06, 
    8.832153e-06, 8.836281e-06, 8.818138e-06, 8.817035e-06, 8.800458e-06, 
    8.815219e-06, 8.821497e-06, 8.837493e-06, 8.846935e-06, 8.855924e-06, 
    8.875699e-06, 8.897788e-06, 8.928746e-06, 8.951029e-06, 8.965972e-06, 
    8.956818e-06, 8.964899e-06, 8.95586e-06, 8.95163e-06, 8.998677e-06, 
    8.972238e-06, 9.01194e-06, 9.009746e-06, 8.991762e-06, 9.009994e-06, 
    8.832775e-06, 8.827691e-06, 8.810006e-06, 8.823846e-06, 8.798655e-06, 
    8.812736e-06, 8.820827e-06, 8.852144e-06, 8.85906e-06, 8.865435e-06, 
    8.878063e-06, 8.894265e-06, 8.922705e-06, 8.947496e-06, 8.970168e-06, 
    8.968508e-06, 8.969091e-06, 8.974145e-06, 8.961611e-06, 8.976205e-06, 
    8.978643e-06, 8.97225e-06, 9.009452e-06, 8.99882e-06, 9.0097e-06, 
    9.00278e-06, 8.829346e-06, 8.837909e-06, 8.83328e-06, 8.841978e-06, 
    8.83584e-06, 8.863111e-06, 8.871293e-06, 8.90966e-06, 8.893939e-06, 
    8.919e-06, 8.896493e-06, 8.900472e-06, 8.919764e-06, 8.897718e-06, 
    8.946105e-06, 8.913242e-06, 8.974342e-06, 8.941437e-06, 8.976403e-06, 
    8.97007e-06, 8.980568e-06, 8.98996e-06, 9.001806e-06, 9.023637e-06, 
    9.018585e-06, 9.036874e-06, 8.85069e-06, 8.861795e-06, 8.860841e-06, 
    8.872484e-06, 8.881094e-06, 8.899799e-06, 8.929798e-06, 8.918521e-06, 
    8.939255e-06, 8.943411e-06, 8.911926e-06, 8.93123e-06, 8.869248e-06, 
    8.879226e-06, 8.873301e-06, 8.851553e-06, 8.921086e-06, 8.885359e-06, 
    8.951393e-06, 8.932015e-06, 8.988618e-06, 8.960428e-06, 9.015799e-06, 
    9.039441e-06, 9.061824e-06, 9.087871e-06, 8.867883e-06, 8.860334e-06, 
    8.873875e-06, 8.892585e-06, 8.910025e-06, 8.933192e-06, 8.935577e-06, 
    8.939913e-06, 8.951177e-06, 8.960639e-06, 8.941261e-06, 8.963014e-06, 
    8.881493e-06, 8.9242e-06, 8.857457e-06, 8.877501e-06, 8.891492e-06, 
    8.885378e-06, 8.917238e-06, 8.924744e-06, 8.955262e-06, 8.939495e-06, 
    9.033583e-06, 8.991911e-06, 9.107802e-06, 9.075351e-06, 8.85769e-06, 
    8.867869e-06, 8.903301e-06, 8.886439e-06, 8.934752e-06, 8.946648e-06, 
    8.956343e-06, 8.968703e-06, 8.970055e-06, 8.977385e-06, 8.965372e-06, 
    8.976919e-06, 8.933242e-06, 8.952755e-06, 8.899277e-06, 8.912269e-06, 
    8.9063e-06, 8.899736e-06, 8.919996e-06, 8.941559e-06, 8.942059e-06, 
    8.94897e-06, 8.968388e-06, 8.934949e-06, 9.038895e-06, 8.974584e-06, 
    8.878972e-06, 8.898552e-06, 8.901397e-06, 8.8938e-06, 8.945453e-06, 
    8.926721e-06, 8.977211e-06, 8.963564e-06, 8.985939e-06, 8.974815e-06, 
    8.973177e-06, 8.958906e-06, 8.950014e-06, 8.927572e-06, 8.909337e-06, 
    8.894907e-06, 8.898265e-06, 8.914119e-06, 8.942888e-06, 8.970161e-06, 
    8.964178e-06, 8.984238e-06, 8.931244e-06, 8.953432e-06, 8.944841e-06, 
    8.967255e-06, 8.918212e-06, 8.959852e-06, 8.907567e-06, 8.912154e-06, 
    8.926349e-06, 8.954912e-06, 8.961293e-06, 8.968038e-06, 8.963884e-06, 
    8.943626e-06, 8.940326e-06, 8.926014e-06, 8.922045e-06, 8.911158e-06, 
    8.902131e-06, 8.910369e-06, 8.919015e-06, 8.943651e-06, 8.96585e-06, 
    8.990089e-06, 8.996039e-06, 9.024297e-06, 9.001238e-06, 9.039245e-06, 
    9.006848e-06, 9.062994e-06, 8.962324e-06, 9.005974e-06, 8.927009e-06, 
    8.935514e-06, 8.950862e-06, 8.986183e-06, 8.967149e-06, 8.98943e-06, 
    8.940199e-06, 8.914648e-06, 8.908089e-06, 8.895777e-06, 8.908371e-06, 
    8.907347e-06, 8.919401e-06, 8.915529e-06, 8.944469e-06, 8.928921e-06, 
    8.973125e-06, 8.989264e-06, 9.034942e-06, 9.062957e-06, 9.091566e-06, 
    9.104185e-06, 9.10803e-06, 9.109635e-06 ;

 QVEGE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 QVEGT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RAIN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RETRANSN =
  4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 4.331019e-07, 
    4.331019e-07, 4.331019e-07, 4.331019e-07 ;

 RETRANSN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 RH2M =
  81.68652, 81.68572, 81.68587, 81.68524, 81.68559, 81.68517, 81.68635, 
    81.6857, 81.68611, 81.68644, 81.68403, 81.68521, 81.68273, 81.6835, 
    81.68156, 81.68286, 81.68129, 81.68158, 81.68067, 81.68093, 81.6798, 
    81.68055, 81.67919, 81.67997, 81.67986, 81.68058, 81.68496, 81.68418, 
    81.68501, 81.68489, 81.68494, 81.68559, 81.68591, 81.68657, 81.68645, 
    81.68596, 81.68484, 81.68521, 81.68425, 81.68427, 81.68321, 81.68369, 
    81.68189, 81.6824, 81.68092, 81.6813, 81.68094, 81.68105, 81.68094, 
    81.68149, 81.68125, 81.68173, 81.6836, 81.68306, 81.68469, 81.68569, 
    81.68633, 81.68678, 81.68671, 81.68659, 81.68596, 81.68535, 81.68488, 
    81.68458, 81.68427, 81.6834, 81.68289, 81.6818, 81.68198, 81.68166, 
    81.68133, 81.6808, 81.68089, 81.68065, 81.68166, 81.68099, 81.68209, 
    81.68179, 81.68425, 81.68511, 81.68552, 81.68584, 81.68667, 81.6861, 
    81.68633, 81.68578, 81.68545, 81.68561, 81.68457, 81.68497, 81.68286, 
    81.68378, 81.68137, 81.68195, 81.68123, 81.68159, 81.68098, 81.68153, 
    81.68056, 81.68036, 81.6805, 81.67994, 81.68156, 81.68095, 81.68562, 
    81.68559, 81.68546, 81.68604, 81.68607, 81.68657, 81.68612, 81.68593, 
    81.68542, 81.68513, 81.68485, 81.68424, 81.68356, 81.68261, 81.68191, 
    81.68144, 81.68172, 81.68147, 81.68176, 81.68188, 81.68044, 81.68125, 
    81.68002, 81.68008, 81.68065, 81.68008, 81.68557, 81.68572, 81.68628, 
    81.68584, 81.68663, 81.6862, 81.68595, 81.68498, 81.68475, 81.68456, 
    81.68417, 81.68367, 81.68279, 81.68202, 81.68131, 81.68136, 81.68134, 
    81.68119, 81.68158, 81.68113, 81.68105, 81.68125, 81.68009, 81.68042, 
    81.68008, 81.6803, 81.68568, 81.68541, 81.68555, 81.68529, 81.68548, 
    81.68465, 81.68439, 81.6832, 81.68368, 81.68291, 81.68359, 81.68348, 
    81.68291, 81.68356, 81.68208, 81.6831, 81.68118, 81.68223, 81.68112, 
    81.68131, 81.68098, 81.6807, 81.68033, 81.67966, 81.67982, 81.67925, 
    81.68501, 81.68468, 81.6847, 81.68434, 81.68407, 81.68349, 81.68256, 
    81.68291, 81.68227, 81.68214, 81.68311, 81.68253, 81.68445, 81.68414, 
    81.68432, 81.68499, 81.68285, 81.68395, 81.6819, 81.6825, 81.68074, 
    81.68163, 81.6799, 81.67919, 81.67847, 81.67769, 81.68449, 81.68472, 
    81.6843, 81.68373, 81.68318, 81.68246, 81.68238, 81.68225, 81.6819, 
    81.6816, 81.68222, 81.68153, 81.6841, 81.68275, 81.68481, 81.6842, 
    81.68376, 81.68394, 81.68295, 81.68272, 81.68179, 81.68226, 81.67937, 
    81.68066, 81.67706, 81.67807, 81.6848, 81.68448, 81.6834, 81.68391, 
    81.68241, 81.68204, 81.68174, 81.68137, 81.68131, 81.68109, 81.68146, 
    81.6811, 81.68246, 81.68185, 81.6835, 81.68311, 81.68329, 81.68349, 
    81.68286, 81.68221, 81.68218, 81.68198, 81.68142, 81.6824, 81.67924, 
    81.68122, 81.68414, 81.68355, 81.68345, 81.68368, 81.68208, 81.68266, 
    81.68109, 81.68152, 81.68082, 81.68117, 81.68122, 81.68166, 81.68194, 
    81.68264, 81.6832, 81.68364, 81.68354, 81.68305, 81.68217, 81.68132, 
    81.6815, 81.68088, 81.68252, 81.68184, 81.68211, 81.6814, 81.68292, 
    81.68168, 81.68325, 81.68311, 81.68267, 81.6818, 81.68159, 81.68138, 
    81.6815, 81.68214, 81.68224, 81.68268, 81.68281, 81.68314, 81.68342, 
    81.68317, 81.68291, 81.68214, 81.68145, 81.6807, 81.68051, 81.67967, 
    81.68037, 81.67923, 81.68024, 81.67848, 81.68158, 81.68024, 81.68265, 
    81.68238, 81.68192, 81.68083, 81.6814, 81.68073, 81.68224, 81.68304, 
    81.68324, 81.68362, 81.68323, 81.68326, 81.68288, 81.683, 81.68211, 
    81.68259, 81.68123, 81.68073, 81.67931, 81.67846, 81.67755, 81.67716, 
    81.67704, 81.67699 ;

 RH2M_R =
  81.68652, 81.68572, 81.68587, 81.68524, 81.68559, 81.68517, 81.68635, 
    81.6857, 81.68611, 81.68644, 81.68403, 81.68521, 81.68273, 81.6835, 
    81.68156, 81.68286, 81.68129, 81.68158, 81.68067, 81.68093, 81.6798, 
    81.68055, 81.67919, 81.67997, 81.67986, 81.68058, 81.68496, 81.68418, 
    81.68501, 81.68489, 81.68494, 81.68559, 81.68591, 81.68657, 81.68645, 
    81.68596, 81.68484, 81.68521, 81.68425, 81.68427, 81.68321, 81.68369, 
    81.68189, 81.6824, 81.68092, 81.6813, 81.68094, 81.68105, 81.68094, 
    81.68149, 81.68125, 81.68173, 81.6836, 81.68306, 81.68469, 81.68569, 
    81.68633, 81.68678, 81.68671, 81.68659, 81.68596, 81.68535, 81.68488, 
    81.68458, 81.68427, 81.6834, 81.68289, 81.6818, 81.68198, 81.68166, 
    81.68133, 81.6808, 81.68089, 81.68065, 81.68166, 81.68099, 81.68209, 
    81.68179, 81.68425, 81.68511, 81.68552, 81.68584, 81.68667, 81.6861, 
    81.68633, 81.68578, 81.68545, 81.68561, 81.68457, 81.68497, 81.68286, 
    81.68378, 81.68137, 81.68195, 81.68123, 81.68159, 81.68098, 81.68153, 
    81.68056, 81.68036, 81.6805, 81.67994, 81.68156, 81.68095, 81.68562, 
    81.68559, 81.68546, 81.68604, 81.68607, 81.68657, 81.68612, 81.68593, 
    81.68542, 81.68513, 81.68485, 81.68424, 81.68356, 81.68261, 81.68191, 
    81.68144, 81.68172, 81.68147, 81.68176, 81.68188, 81.68044, 81.68125, 
    81.68002, 81.68008, 81.68065, 81.68008, 81.68557, 81.68572, 81.68628, 
    81.68584, 81.68663, 81.6862, 81.68595, 81.68498, 81.68475, 81.68456, 
    81.68417, 81.68367, 81.68279, 81.68202, 81.68131, 81.68136, 81.68134, 
    81.68119, 81.68158, 81.68113, 81.68105, 81.68125, 81.68009, 81.68042, 
    81.68008, 81.6803, 81.68568, 81.68541, 81.68555, 81.68529, 81.68548, 
    81.68465, 81.68439, 81.6832, 81.68368, 81.68291, 81.68359, 81.68348, 
    81.68291, 81.68356, 81.68208, 81.6831, 81.68118, 81.68223, 81.68112, 
    81.68131, 81.68098, 81.6807, 81.68033, 81.67966, 81.67982, 81.67925, 
    81.68501, 81.68468, 81.6847, 81.68434, 81.68407, 81.68349, 81.68256, 
    81.68291, 81.68227, 81.68214, 81.68311, 81.68253, 81.68445, 81.68414, 
    81.68432, 81.68499, 81.68285, 81.68395, 81.6819, 81.6825, 81.68074, 
    81.68163, 81.6799, 81.67919, 81.67847, 81.67769, 81.68449, 81.68472, 
    81.6843, 81.68373, 81.68318, 81.68246, 81.68238, 81.68225, 81.6819, 
    81.6816, 81.68222, 81.68153, 81.6841, 81.68275, 81.68481, 81.6842, 
    81.68376, 81.68394, 81.68295, 81.68272, 81.68179, 81.68226, 81.67937, 
    81.68066, 81.67706, 81.67807, 81.6848, 81.68448, 81.6834, 81.68391, 
    81.68241, 81.68204, 81.68174, 81.68137, 81.68131, 81.68109, 81.68146, 
    81.6811, 81.68246, 81.68185, 81.6835, 81.68311, 81.68329, 81.68349, 
    81.68286, 81.68221, 81.68218, 81.68198, 81.68142, 81.6824, 81.67924, 
    81.68122, 81.68414, 81.68355, 81.68345, 81.68368, 81.68208, 81.68266, 
    81.68109, 81.68152, 81.68082, 81.68117, 81.68122, 81.68166, 81.68194, 
    81.68264, 81.6832, 81.68364, 81.68354, 81.68305, 81.68217, 81.68132, 
    81.6815, 81.68088, 81.68252, 81.68184, 81.68211, 81.6814, 81.68292, 
    81.68168, 81.68325, 81.68311, 81.68267, 81.6818, 81.68159, 81.68138, 
    81.6815, 81.68214, 81.68224, 81.68268, 81.68281, 81.68314, 81.68342, 
    81.68317, 81.68291, 81.68214, 81.68145, 81.6807, 81.68051, 81.67967, 
    81.68037, 81.67923, 81.68024, 81.67848, 81.68158, 81.68024, 81.68265, 
    81.68238, 81.68192, 81.68083, 81.6814, 81.68073, 81.68224, 81.68304, 
    81.68324, 81.68362, 81.68323, 81.68326, 81.68288, 81.683, 81.68211, 
    81.68259, 81.68123, 81.68073, 81.67931, 81.67846, 81.67755, 81.67716, 
    81.67704, 81.67699 ;

 RH2M_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 RR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABG =
  0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 0.05229128, 
    0.05229128, 0.05229128 ;

 SABG_PEN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SABV =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SEEDN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN =
  0.0004362622, 0.0004381055, 0.0004377471, 0.0004392338, 0.000438409, 
    0.0004393824, 0.0004366357, 0.0004381783, 0.0004371935, 0.0004364277, 
    0.0004421185, 0.0004392997, 0.0004450469, 0.0004432489, 0.0004477654, 
    0.0004447669, 0.0004483699, 0.0004476788, 0.0004497589, 0.0004491629, 
    0.0004518233, 0.0004500338, 0.0004532024, 0.0004513958, 0.0004516784, 
    0.0004499745, 0.0004398674, 0.0004417679, 0.0004397547, 0.0004400257, 
    0.000439904, 0.0004384258, 0.0004376808, 0.0004361209, 0.000436404, 
    0.0004375498, 0.0004401472, 0.0004392654, 0.0004414876, 0.0004414374, 
    0.0004439113, 0.0004427959, 0.0004469542, 0.0004457723, 0.0004491877, 
    0.0004483286, 0.0004491473, 0.0004488989, 0.0004491503, 0.0004478905, 
    0.0004484302, 0.0004473217, 0.0004430054, 0.0004442741, 0.0004404899, 
    0.0004382143, 0.0004367031, 0.0004356307, 0.0004357822, 0.0004360712, 
    0.0004375563, 0.0004389527, 0.0004400169, 0.0004407287, 0.00044143, 
    0.000443553, 0.0004446768, 0.0004471931, 0.000446739, 0.0004475082, 
    0.0004482431, 0.0004494769, 0.0004492739, 0.0004498174, 0.0004474876, 
    0.0004490359, 0.0004464799, 0.0004471789, 0.000441621, 0.0004395035, 
    0.0004386033, 0.0004378155, 0.0004358987, 0.0004372223, 0.0004367005, 
    0.0004379418, 0.0004387306, 0.0004383404, 0.0004407481, 0.0004398119, 
    0.0004447433, 0.0004426192, 0.0004481575, 0.0004468321, 0.000448475, 
    0.0004476366, 0.000449073, 0.0004477802, 0.0004500196, 0.0004505072, 
    0.0004501739, 0.0004514541, 0.0004477082, 0.0004491467, 0.0004383297, 
    0.0004383934, 0.0004386897, 0.0004373866, 0.0004373069, 0.0004361128, 
    0.0004371752, 0.0004376276, 0.0004387762, 0.0004394554, 0.0004401012, 
    0.0004415212, 0.000443107, 0.0004453246, 0.0004469179, 0.0004479859, 
    0.000447331, 0.0004479091, 0.0004472627, 0.0004469597, 0.0004503244, 
    0.000448435, 0.0004512698, 0.000451113, 0.0004498299, 0.0004511305, 
    0.0004384379, 0.0004380717, 0.0004368005, 0.0004377952, 0.0004359827, 
    0.0004369972, 0.0004375805, 0.0004398313, 0.0004403259, 0.0004407845, 
    0.0004416902, 0.0004428525, 0.0004448917, 0.0004466659, 0.0004482857, 
    0.0004481669, 0.0004482087, 0.0004485704, 0.0004476741, 0.0004487174, 
    0.0004488925, 0.0004484346, 0.0004510918, 0.0004503326, 0.0004511094, 
    0.000450615, 0.0004381907, 0.0004388067, 0.0004384737, 0.0004390997, 
    0.0004386585, 0.0004406196, 0.0004412075, 0.0004439588, 0.0004428296, 
    0.0004446267, 0.0004430121, 0.0004432982, 0.000444685, 0.0004430992, 
    0.0004465678, 0.000444216, 0.0004485844, 0.0004462357, 0.0004487315, 
    0.0004482782, 0.0004490285, 0.0004497005, 0.0004505458, 0.0004521057, 
    0.0004517444, 0.000453049, 0.0004397251, 0.000440524, 0.0004404537, 
    0.0004412899, 0.0004419083, 0.0004432489, 0.0004453989, 0.0004445903, 
    0.0004460746, 0.0004463725, 0.0004441174, 0.0004455019, 0.0004410583, 
    0.0004417761, 0.0004413487, 0.0004397873, 0.0004447761, 0.0004422156, 
    0.0004469436, 0.0004455564, 0.0004496045, 0.0004475912, 0.0004515455, 
    0.0004532359, 0.000454827, 0.0004566862, 0.0004409602, 0.0004404171, 
    0.0004413893, 0.0004427343, 0.0004439824, 0.0004456417, 0.0004458114, 
    0.0004461222, 0.0004469274, 0.0004476044, 0.0004462203, 0.000447774, 
    0.0004419424, 0.0004449983, 0.0004402111, 0.0004416525, 0.0004426543, 
    0.0004422149, 0.0004444972, 0.000445035, 0.0004472209, 0.0004460909, 
    0.0004528185, 0.000449842, 0.0004581019, 0.0004557935, 0.0004402273, 
    0.0004409581, 0.0004435015, 0.0004422913, 0.0004457523, 0.0004466043, 
    0.0004472968, 0.0004481821, 0.0004482776, 0.0004488022, 0.0004479425, 
    0.0004487681, 0.0004456446, 0.0004470404, 0.0004432102, 0.0004441423, 
    0.0004437135, 0.000443243, 0.0004446947, 0.0004462414, 0.0004462745, 
    0.0004467704, 0.0004481677, 0.0004457654, 0.0004532023, 0.0004486091, 
    0.0004417549, 0.0004431625, 0.0004433636, 0.0004428183, 0.0004465187, 
    0.0004451779, 0.0004487894, 0.0004478132, 0.0004494125, 0.0004486178, 
    0.0004485007, 0.00044748, 0.0004468444, 0.0004452389, 0.0004439325, 
    0.0004428967, 0.0004431375, 0.0004442753, 0.0004463359, 0.0004482855, 
    0.0004478584, 0.0004492902, 0.0004455002, 0.0004470894, 0.0004464751, 
    0.0004480767, 0.0004445686, 0.0004475566, 0.0004438047, 0.0004441336, 
    0.0004451511, 0.0004471979, 0.0004476508, 0.0004481343, 0.0004478359, 
    0.0004463887, 0.0004461515, 0.000445126, 0.0004448428, 0.0004440615, 
    0.0004434145, 0.0004440055, 0.000444626, 0.0004463889, 0.0004479774, 
    0.0004497094, 0.0004501333, 0.0004521567, 0.0004505093, 0.0004532276, 
    0.0004509163, 0.0004549173, 0.0004477297, 0.0004508496, 0.0004451974, 
    0.0004458063, 0.0004469075, 0.0004494335, 0.0004480698, 0.0004496647, 
    0.0004461422, 0.0004443146, 0.0004438418, 0.0004429596, 0.0004438618, 
    0.0004437884, 0.0004446518, 0.0004443743, 0.0004464472, 0.0004453337, 
    0.000448497, 0.0004496514, 0.0004529117, 0.0004549102, 0.0004569448, 
    0.000457843, 0.0004581164, 0.0004582306 ;

 SMINN_TO_NPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_PLANT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMINN_TO_SOIL1N_L1 =
  3.476285e-14, 3.485807e-14, 3.483957e-14, 3.491631e-14, 3.487376e-14, 
    3.492399e-14, 3.478217e-14, 3.486183e-14, 3.4811e-14, 3.477145e-14, 
    3.506505e-14, 3.491974e-14, 3.521595e-14, 3.512339e-14, 3.535582e-14, 
    3.520153e-14, 3.538691e-14, 3.53514e-14, 3.545831e-14, 3.54277e-14, 
    3.556425e-14, 3.547244e-14, 3.563502e-14, 3.554235e-14, 3.555683e-14, 
    3.54694e-14, 3.494903e-14, 3.504696e-14, 3.494321e-14, 3.495719e-14, 
    3.495092e-14, 3.487463e-14, 3.483614e-14, 3.475559e-14, 3.477023e-14, 
    3.48294e-14, 3.496347e-14, 3.491799e-14, 3.503263e-14, 3.503005e-14, 
    3.515753e-14, 3.510007e-14, 3.531415e-14, 3.525335e-14, 3.542898e-14, 
    3.538483e-14, 3.54269e-14, 3.541415e-14, 3.542706e-14, 3.536231e-14, 
    3.539006e-14, 3.533307e-14, 3.511082e-14, 3.517617e-14, 3.498114e-14, 
    3.486367e-14, 3.478566e-14, 3.473026e-14, 3.473809e-14, 3.475302e-14, 
    3.482974e-14, 3.490186e-14, 3.495678e-14, 3.49935e-14, 3.502967e-14, 
    3.513902e-14, 3.519692e-14, 3.532642e-14, 3.530309e-14, 3.534263e-14, 
    3.538044e-14, 3.544384e-14, 3.543341e-14, 3.546133e-14, 3.534161e-14, 
    3.542118e-14, 3.528979e-14, 3.532574e-14, 3.503939e-14, 3.493027e-14, 
    3.488376e-14, 3.484312e-14, 3.474411e-14, 3.481249e-14, 3.478554e-14, 
    3.484967e-14, 3.489039e-14, 3.487026e-14, 3.499451e-14, 3.494621e-14, 
    3.520035e-14, 3.509095e-14, 3.537603e-14, 3.530788e-14, 3.539236e-14, 
    3.534927e-14, 3.542308e-14, 3.535665e-14, 3.547172e-14, 3.549675e-14, 
    3.547965e-14, 3.554538e-14, 3.535296e-14, 3.542688e-14, 3.486969e-14, 
    3.487297e-14, 3.488828e-14, 3.482098e-14, 3.481686e-14, 3.475519e-14, 
    3.481008e-14, 3.483344e-14, 3.489276e-14, 3.492782e-14, 3.496114e-14, 
    3.503437e-14, 3.511609e-14, 3.52303e-14, 3.53123e-14, 3.536722e-14, 
    3.533356e-14, 3.536328e-14, 3.533005e-14, 3.531447e-14, 3.548737e-14, 
    3.539031e-14, 3.553593e-14, 3.552788e-14, 3.546199e-14, 3.552878e-14, 
    3.487528e-14, 3.485638e-14, 3.479071e-14, 3.484211e-14, 3.474847e-14, 
    3.480088e-14, 3.483099e-14, 3.49472e-14, 3.497274e-14, 3.499639e-14, 
    3.50431e-14, 3.510301e-14, 3.520802e-14, 3.529933e-14, 3.538264e-14, 
    3.537654e-14, 3.537869e-14, 3.539728e-14, 3.53512e-14, 3.540484e-14, 
    3.541383e-14, 3.539031e-14, 3.55268e-14, 3.548782e-14, 3.552771e-14, 
    3.550233e-14, 3.486253e-14, 3.489433e-14, 3.487714e-14, 3.490945e-14, 
    3.488668e-14, 3.498785e-14, 3.501817e-14, 3.515996e-14, 3.510182e-14, 
    3.519437e-14, 3.511123e-14, 3.512596e-14, 3.519734e-14, 3.511574e-14, 
    3.529427e-14, 3.517322e-14, 3.5398e-14, 3.527717e-14, 3.540556e-14, 
    3.538228e-14, 3.542084e-14, 3.545535e-14, 3.549877e-14, 3.557882e-14, 
    3.556029e-14, 3.562722e-14, 3.494173e-14, 3.498294e-14, 3.497933e-14, 
    3.502246e-14, 3.505433e-14, 3.512343e-14, 3.523413e-14, 3.519252e-14, 
    3.526893e-14, 3.528425e-14, 3.516818e-14, 3.523944e-14, 3.501052e-14, 
    3.504752e-14, 3.502551e-14, 3.494497e-14, 3.520208e-14, 3.507019e-14, 
    3.531365e-14, 3.524229e-14, 3.545043e-14, 3.534694e-14, 3.555009e-14, 
    3.563676e-14, 3.571837e-14, 3.581353e-14, 3.500544e-14, 3.497745e-14, 
    3.502759e-14, 3.509689e-14, 3.516121e-14, 3.524664e-14, 3.525538e-14, 
    3.527137e-14, 3.531281e-14, 3.534762e-14, 3.527641e-14, 3.535635e-14, 
    3.505605e-14, 3.521353e-14, 3.496684e-14, 3.504115e-14, 3.509281e-14, 
    3.507018e-14, 3.518777e-14, 3.521547e-14, 3.532791e-14, 3.526981e-14, 
    3.561535e-14, 3.546261e-14, 3.5886e-14, 3.576784e-14, 3.496766e-14, 
    3.500536e-14, 3.513643e-14, 3.507409e-14, 3.525235e-14, 3.529617e-14, 
    3.533181e-14, 3.537731e-14, 3.538224e-14, 3.540919e-14, 3.536502e-14, 
    3.540745e-14, 3.524682e-14, 3.531863e-14, 3.512148e-14, 3.516949e-14, 
    3.514742e-14, 3.512318e-14, 3.519795e-14, 3.527753e-14, 3.527926e-14, 
    3.530476e-14, 3.537651e-14, 3.525307e-14, 3.563499e-14, 3.539922e-14, 
    3.504645e-14, 3.511895e-14, 3.512935e-14, 3.510126e-14, 3.529178e-14, 
    3.522278e-14, 3.540854e-14, 3.535837e-14, 3.544056e-14, 3.539973e-14, 
    3.539372e-14, 3.534125e-14, 3.530856e-14, 3.522594e-14, 3.515868e-14, 
    3.510534e-14, 3.511775e-14, 3.517634e-14, 3.52824e-14, 3.538267e-14, 
    3.53607e-14, 3.543432e-14, 3.523943e-14, 3.532118e-14, 3.528958e-14, 
    3.537196e-14, 3.519141e-14, 3.534507e-14, 3.515209e-14, 3.516903e-14, 
    3.522141e-14, 3.532669e-14, 3.535003e-14, 3.537487e-14, 3.535955e-14, 
    3.52851e-14, 3.527291e-14, 3.522015e-14, 3.520556e-14, 3.516535e-14, 
    3.513202e-14, 3.516246e-14, 3.519441e-14, 3.528514e-14, 3.536683e-14, 
    3.545584e-14, 3.547762e-14, 3.558141e-14, 3.549688e-14, 3.563629e-14, 
    3.551771e-14, 3.572294e-14, 3.535402e-14, 3.551429e-14, 3.522381e-14, 
    3.525514e-14, 3.531177e-14, 3.544161e-14, 3.537157e-14, 3.545349e-14, 
    3.527243e-14, 3.517834e-14, 3.515403e-14, 3.510858e-14, 3.515507e-14, 
    3.515129e-14, 3.519575e-14, 3.518147e-14, 3.528815e-14, 3.523086e-14, 
    3.539355e-14, 3.545286e-14, 3.562019e-14, 3.572262e-14, 3.582684e-14, 
    3.587279e-14, 3.588678e-14, 3.589262e-14 ;

 SMINN_TO_SOIL1N_L2 =
  1.15589e-14, 1.159059e-14, 1.158443e-14, 1.160997e-14, 1.159581e-14, 
    1.161253e-14, 1.156533e-14, 1.159184e-14, 1.157492e-14, 1.156176e-14, 
    1.165948e-14, 1.161111e-14, 1.170971e-14, 1.16789e-14, 1.175627e-14, 
    1.170491e-14, 1.176661e-14, 1.17548e-14, 1.179038e-14, 1.178019e-14, 
    1.182564e-14, 1.179508e-14, 1.18492e-14, 1.181835e-14, 1.182317e-14, 
    1.179407e-14, 1.162086e-14, 1.165346e-14, 1.161893e-14, 1.162358e-14, 
    1.16215e-14, 1.15961e-14, 1.158329e-14, 1.155648e-14, 1.156135e-14, 
    1.158105e-14, 1.162567e-14, 1.161054e-14, 1.164869e-14, 1.164783e-14, 
    1.169026e-14, 1.167114e-14, 1.174239e-14, 1.172216e-14, 1.178062e-14, 
    1.176592e-14, 1.177992e-14, 1.177568e-14, 1.177998e-14, 1.175843e-14, 
    1.176766e-14, 1.174869e-14, 1.167472e-14, 1.169647e-14, 1.163155e-14, 
    1.159245e-14, 1.156649e-14, 1.154805e-14, 1.155066e-14, 1.155562e-14, 
    1.158116e-14, 1.160517e-14, 1.162345e-14, 1.163567e-14, 1.164771e-14, 
    1.16841e-14, 1.170338e-14, 1.174648e-14, 1.173871e-14, 1.175188e-14, 
    1.176446e-14, 1.178556e-14, 1.178209e-14, 1.179138e-14, 1.175154e-14, 
    1.177802e-14, 1.173429e-14, 1.174625e-14, 1.165094e-14, 1.161462e-14, 
    1.159914e-14, 1.158562e-14, 1.155266e-14, 1.157542e-14, 1.156645e-14, 
    1.15878e-14, 1.160135e-14, 1.159465e-14, 1.1636e-14, 1.161993e-14, 
    1.170452e-14, 1.166811e-14, 1.176299e-14, 1.174031e-14, 1.176843e-14, 
    1.175408e-14, 1.177866e-14, 1.175654e-14, 1.179484e-14, 1.180318e-14, 
    1.179748e-14, 1.181936e-14, 1.175532e-14, 1.177992e-14, 1.159446e-14, 
    1.159555e-14, 1.160065e-14, 1.157824e-14, 1.157688e-14, 1.155635e-14, 
    1.157462e-14, 1.158239e-14, 1.160214e-14, 1.161381e-14, 1.16249e-14, 
    1.164927e-14, 1.167647e-14, 1.171449e-14, 1.174178e-14, 1.176006e-14, 
    1.174886e-14, 1.175875e-14, 1.174769e-14, 1.17425e-14, 1.180005e-14, 
    1.176774e-14, 1.181621e-14, 1.181354e-14, 1.17916e-14, 1.181384e-14, 
    1.159632e-14, 1.159003e-14, 1.156817e-14, 1.158528e-14, 1.155411e-14, 
    1.157155e-14, 1.158158e-14, 1.162026e-14, 1.162876e-14, 1.163663e-14, 
    1.165218e-14, 1.167212e-14, 1.170707e-14, 1.173746e-14, 1.176519e-14, 
    1.176316e-14, 1.176388e-14, 1.177006e-14, 1.175473e-14, 1.177258e-14, 
    1.177557e-14, 1.176775e-14, 1.181318e-14, 1.18002e-14, 1.181348e-14, 
    1.180503e-14, 1.159207e-14, 1.160266e-14, 1.159694e-14, 1.160769e-14, 
    1.160011e-14, 1.163379e-14, 1.164388e-14, 1.169107e-14, 1.167172e-14, 
    1.170253e-14, 1.167486e-14, 1.167976e-14, 1.170352e-14, 1.167635e-14, 
    1.173578e-14, 1.169549e-14, 1.177031e-14, 1.173009e-14, 1.177282e-14, 
    1.176507e-14, 1.177791e-14, 1.17894e-14, 1.180385e-14, 1.183049e-14, 
    1.182433e-14, 1.18466e-14, 1.161844e-14, 1.163215e-14, 1.163095e-14, 
    1.164531e-14, 1.165592e-14, 1.167891e-14, 1.171576e-14, 1.170191e-14, 
    1.172734e-14, 1.173244e-14, 1.169381e-14, 1.171753e-14, 1.164133e-14, 
    1.165365e-14, 1.164632e-14, 1.161951e-14, 1.170509e-14, 1.166119e-14, 
    1.174223e-14, 1.171848e-14, 1.178776e-14, 1.175331e-14, 1.182093e-14, 
    1.184978e-14, 1.187694e-14, 1.190862e-14, 1.163964e-14, 1.163032e-14, 
    1.164701e-14, 1.167008e-14, 1.169149e-14, 1.171992e-14, 1.172284e-14, 
    1.172816e-14, 1.174195e-14, 1.175354e-14, 1.172983e-14, 1.175644e-14, 
    1.165649e-14, 1.170891e-14, 1.16268e-14, 1.165153e-14, 1.166872e-14, 
    1.166119e-14, 1.170033e-14, 1.170955e-14, 1.174698e-14, 1.172764e-14, 
    1.184265e-14, 1.179181e-14, 1.193274e-14, 1.189341e-14, 1.162707e-14, 
    1.163961e-14, 1.168324e-14, 1.166249e-14, 1.172183e-14, 1.173641e-14, 
    1.174827e-14, 1.176342e-14, 1.176506e-14, 1.177403e-14, 1.175933e-14, 
    1.177345e-14, 1.171998e-14, 1.174389e-14, 1.167827e-14, 1.169424e-14, 
    1.16869e-14, 1.167883e-14, 1.170372e-14, 1.173021e-14, 1.173078e-14, 
    1.173927e-14, 1.176315e-14, 1.172207e-14, 1.184919e-14, 1.177071e-14, 
    1.165329e-14, 1.167742e-14, 1.168088e-14, 1.167154e-14, 1.173495e-14, 
    1.171198e-14, 1.177381e-14, 1.175712e-14, 1.178447e-14, 1.177088e-14, 
    1.176888e-14, 1.175141e-14, 1.174053e-14, 1.171304e-14, 1.169065e-14, 
    1.167289e-14, 1.167702e-14, 1.169652e-14, 1.173183e-14, 1.17652e-14, 
    1.175789e-14, 1.17824e-14, 1.171753e-14, 1.174473e-14, 1.173422e-14, 
    1.176164e-14, 1.170154e-14, 1.175269e-14, 1.168845e-14, 1.169409e-14, 
    1.171153e-14, 1.174657e-14, 1.175434e-14, 1.176261e-14, 1.175751e-14, 
    1.173273e-14, 1.172867e-14, 1.171111e-14, 1.170625e-14, 1.169287e-14, 
    1.168178e-14, 1.16919e-14, 1.170254e-14, 1.173274e-14, 1.175993e-14, 
    1.178956e-14, 1.179681e-14, 1.183136e-14, 1.180322e-14, 1.184962e-14, 
    1.181015e-14, 1.187846e-14, 1.175567e-14, 1.180901e-14, 1.171233e-14, 
    1.172276e-14, 1.17416e-14, 1.178482e-14, 1.176151e-14, 1.178878e-14, 
    1.172851e-14, 1.169719e-14, 1.16891e-14, 1.167397e-14, 1.168944e-14, 
    1.168819e-14, 1.170299e-14, 1.169823e-14, 1.173374e-14, 1.171467e-14, 
    1.176883e-14, 1.178856e-14, 1.184426e-14, 1.187836e-14, 1.191305e-14, 
    1.192835e-14, 1.1933e-14, 1.193495e-14 ;

 SMINN_TO_SOIL1N_S2 =
  -8.146111e-11, -8.18206e-11, -8.175072e-11, -8.204067e-11, -8.187984e-11, 
    -8.206969e-11, -8.1534e-11, -8.183487e-11, -8.16428e-11, -8.149349e-11, 
    -8.260338e-11, -8.205361e-11, -8.317459e-11, -8.282391e-11, 
    -8.370489e-11, -8.312001e-11, -8.382284e-11, -8.368804e-11, 
    -8.409381e-11, -8.397756e-11, -8.449655e-11, -8.414747e-11, 
    -8.476563e-11, -8.44132e-11, -8.446832e-11, -8.413595e-11, -8.216426e-11, 
    -8.253492e-11, -8.21423e-11, -8.219515e-11, -8.217144e-11, -8.188315e-11, 
    -8.173786e-11, -8.143364e-11, -8.148888e-11, -8.171232e-11, 
    -8.221892e-11, -8.204696e-11, -8.248039e-11, -8.247061e-11, 
    -8.295316e-11, -8.273558e-11, -8.354671e-11, -8.331617e-11, 
    -8.398242e-11, -8.381485e-11, -8.397454e-11, -8.392612e-11, 
    -8.397517e-11, -8.372943e-11, -8.383471e-11, -8.361848e-11, 
    -8.277632e-11, -8.302381e-11, -8.228571e-11, -8.18419e-11, -8.154719e-11, 
    -8.133805e-11, -8.136762e-11, -8.142398e-11, -8.171363e-11, 
    -8.198599e-11, -8.219354e-11, -8.233238e-11, -8.24692e-11, -8.288327e-11, 
    -8.310248e-11, -8.359332e-11, -8.350476e-11, -8.365481e-11, 
    -8.379818e-11, -8.403889e-11, -8.399927e-11, -8.410531e-11, 
    -8.365086e-11, -8.395288e-11, -8.345431e-11, -8.359066e-11, 
    -8.250632e-11, -8.209336e-11, -8.191778e-11, -8.176415e-11, 
    -8.139035e-11, -8.164848e-11, -8.154672e-11, -8.178883e-11, 
    -8.194267e-11, -8.186658e-11, -8.233619e-11, -8.215361e-11, 
    -8.311547e-11, -8.270115e-11, -8.378146e-11, -8.352294e-11, 
    -8.384343e-11, -8.367989e-11, -8.39601e-11, -8.370792e-11, -8.414479e-11, 
    -8.423991e-11, -8.41749e-11, -8.442464e-11, -8.369393e-11, -8.397454e-11, 
    -8.186445e-11, -8.187686e-11, -8.193467e-11, -8.168054e-11, 
    -8.166499e-11, -8.143213e-11, -8.163933e-11, -8.172757e-11, 
    -8.195159e-11, -8.208409e-11, -8.221005e-11, -8.2487e-11, -8.279632e-11, 
    -8.322889e-11, -8.35397e-11, -8.374804e-11, -8.362028e-11, -8.373307e-11, 
    -8.360699e-11, -8.35479e-11, -8.420426e-11, -8.38357e-11, -8.438873e-11, 
    -8.435812e-11, -8.410783e-11, -8.436157e-11, -8.188557e-11, 
    -8.181417e-11, -8.156624e-11, -8.176027e-11, -8.140677e-11, 
    -8.160463e-11, -8.17184e-11, -8.215741e-11, -8.225389e-11, -8.234333e-11, 
    -8.251999e-11, -8.274671e-11, -8.314446e-11, -8.349055e-11, 
    -8.380653e-11, -8.378338e-11, -8.379153e-11, -8.386211e-11, 
    -8.368727e-11, -8.389081e-11, -8.392497e-11, -8.383565e-11, 
    -8.435402e-11, -8.420593e-11, -8.435747e-11, -8.426105e-11, 
    -8.183738e-11, -8.195753e-11, -8.18926e-11, -8.201469e-11, -8.192868e-11, 
    -8.231115e-11, -8.242583e-11, -8.296248e-11, -8.274225e-11, 
    -8.309277e-11, -8.277786e-11, -8.283366e-11, -8.310418e-11, 
    -8.279488e-11, -8.347146e-11, -8.301273e-11, -8.386485e-11, 
    -8.340671e-11, -8.389356e-11, -8.380516e-11, -8.395153e-11, 
    -8.408262e-11, -8.424755e-11, -8.455185e-11, -8.448139e-11, -8.47359e-11, 
    -8.213667e-11, -8.229251e-11, -8.22788e-11, -8.244191e-11, -8.256253e-11, 
    -8.282401e-11, -8.324338e-11, -8.308568e-11, -8.337522e-11, 
    -8.343334e-11, -8.299347e-11, -8.326353e-11, -8.239683e-11, 
    -8.253683e-11, -8.245348e-11, -8.214895e-11, -8.312201e-11, 
    -8.262261e-11, -8.354483e-11, -8.327427e-11, -8.406392e-11, 
    -8.367119e-11, -8.44426e-11, -8.477236e-11, -8.508279e-11, -8.544553e-11, 
    -8.237758e-11, -8.227168e-11, -8.246131e-11, -8.272365e-11, 
    -8.296711e-11, -8.329076e-11, -8.332389e-11, -8.338452e-11, -8.35416e-11, 
    -8.367366e-11, -8.340368e-11, -8.370676e-11, -8.256928e-11, 
    -8.316536e-11, -8.223164e-11, -8.251277e-11, -8.270819e-11, 
    -8.262248e-11, -8.306766e-11, -8.317259e-11, -8.359898e-11, 
    -8.337857e-11, -8.469096e-11, -8.411029e-11, -8.572177e-11, 
    -8.527139e-11, -8.223468e-11, -8.237722e-11, -8.287332e-11, 
    -8.263727e-11, -8.331238e-11, -8.347856e-11, -8.361367e-11, 
    -8.378636e-11, -8.380502e-11, -8.390734e-11, -8.373966e-11, 
    -8.390072e-11, -8.329146e-11, -8.356372e-11, -8.281663e-11, 
    -8.299845e-11, -8.291481e-11, -8.282305e-11, -8.310624e-11, 
    -8.340793e-11, -8.341439e-11, -8.351114e-11, -8.37837e-11, -8.331512e-11, 
    -8.476587e-11, -8.386986e-11, -8.253266e-11, -8.28072e-11, -8.284644e-11, 
    -8.274009e-11, -8.34619e-11, -8.320035e-11, -8.390485e-11, -8.371445e-11, 
    -8.402642e-11, -8.387139e-11, -8.384858e-11, -8.364948e-11, 
    -8.352551e-11, -8.321234e-11, -8.295754e-11, -8.275551e-11, 
    -8.280249e-11, -8.302441e-11, -8.342639e-11, -8.38067e-11, -8.372338e-11, 
    -8.400271e-11, -8.326343e-11, -8.357341e-11, -8.345359e-11, 
    -8.376601e-11, -8.308149e-11, -8.366433e-11, -8.293252e-11, 
    -8.299668e-11, -8.319516e-11, -8.359442e-11, -8.368278e-11, -8.37771e-11, 
    -8.37189e-11, -8.34366e-11, -8.339036e-11, -8.319034e-11, -8.31351e-11, 
    -8.298271e-11, -8.285653e-11, -8.297181e-11, -8.309287e-11, 
    -8.343672e-11, -8.374661e-11, -8.408448e-11, -8.416717e-11, 
    -8.456193e-11, -8.424055e-11, -8.477086e-11, -8.431996e-11, 
    -8.510054e-11, -8.369814e-11, -8.430674e-11, -8.320419e-11, 
    -8.332297e-11, -8.353779e-11, -8.403055e-11, -8.376454e-11, 
    -8.407565e-11, -8.338855e-11, -8.303207e-11, -8.293986e-11, 
    -8.276779e-11, -8.294379e-11, -8.292948e-11, -8.30979e-11, -8.304377e-11, 
    -8.344814e-11, -8.323094e-11, -8.3848e-11, -8.40732e-11, -8.470922e-11, 
    -8.509914e-11, -8.54961e-11, -8.567135e-11, -8.57247e-11, -8.5747e-11 ;

 SMINN_TO_SOIL1N_S3 =
  -1.963369e-12, -1.972031e-12, -1.970347e-12, -1.977334e-12, -1.973459e-12, 
    -1.978034e-12, -1.965125e-12, -1.972375e-12, -1.967747e-12, 
    -1.964149e-12, -1.990894e-12, -1.977646e-12, -2.004658e-12, 
    -1.996208e-12, -2.017436e-12, -2.003343e-12, -2.020278e-12, -2.01703e-12, 
    -2.026808e-12, -2.024007e-12, -2.036513e-12, -2.028101e-12, 
    -2.042996e-12, -2.034504e-12, -2.035832e-12, -2.027823e-12, 
    -1.980313e-12, -1.989244e-12, -1.979783e-12, -1.981057e-12, 
    -1.980485e-12, -1.973539e-12, -1.970037e-12, -1.962707e-12, 
    -1.964038e-12, -1.969422e-12, -1.981629e-12, -1.977486e-12, -1.98793e-12, 
    -1.987694e-12, -1.999322e-12, -1.994079e-12, -2.013625e-12, 
    -2.008069e-12, -2.024124e-12, -2.020086e-12, -2.023934e-12, 
    -2.022767e-12, -2.023949e-12, -2.018028e-12, -2.020565e-12, 
    -2.015354e-12, -1.995061e-12, -2.001025e-12, -1.983239e-12, 
    -1.972545e-12, -1.965443e-12, -1.960403e-12, -1.961116e-12, 
    -1.962474e-12, -1.969454e-12, -1.976017e-12, -1.981018e-12, 
    -1.984364e-12, -1.98766e-12, -1.997638e-12, -2.00292e-12, -2.014748e-12, 
    -2.012614e-12, -2.01623e-12, -2.019685e-12, -2.025484e-12, -2.02453e-12, 
    -2.027085e-12, -2.016134e-12, -2.023412e-12, -2.011398e-12, 
    -2.014684e-12, -1.988555e-12, -1.978604e-12, -1.974373e-12, 
    -1.970671e-12, -1.961664e-12, -1.967884e-12, -1.965432e-12, 
    -1.971266e-12, -1.974973e-12, -1.973139e-12, -1.984455e-12, 
    -1.980056e-12, -2.003234e-12, -1.99325e-12, -2.019281e-12, -2.013052e-12, 
    -2.020775e-12, -2.016834e-12, -2.023586e-12, -2.017509e-12, 
    -2.028036e-12, -2.030329e-12, -2.028762e-12, -2.03478e-12, -2.017172e-12, 
    -2.023934e-12, -1.973088e-12, -1.973387e-12, -1.97478e-12, -1.968656e-12, 
    -1.968282e-12, -1.96267e-12, -1.967663e-12, -1.96979e-12, -1.975188e-12, 
    -1.978381e-12, -1.981416e-12, -1.98809e-12, -1.995543e-12, -2.005966e-12, 
    -2.013456e-12, -2.018476e-12, -2.015398e-12, -2.018115e-12, 
    -2.015077e-12, -2.013653e-12, -2.029469e-12, -2.020588e-12, 
    -2.033914e-12, -2.033177e-12, -2.027146e-12, -2.03326e-12, -1.973597e-12, 
    -1.971876e-12, -1.965902e-12, -1.970577e-12, -1.962059e-12, 
    -1.966827e-12, -1.969568e-12, -1.980147e-12, -1.982472e-12, 
    -1.984627e-12, -1.988884e-12, -1.994348e-12, -2.003932e-12, 
    -2.012272e-12, -2.019886e-12, -2.019328e-12, -2.019524e-12, 
    -2.021225e-12, -2.017012e-12, -2.021916e-12, -2.02274e-12, -2.020587e-12, 
    -2.033078e-12, -2.02951e-12, -2.033161e-12, -2.030838e-12, -1.972436e-12, 
    -1.975331e-12, -1.973766e-12, -1.976708e-12, -1.974636e-12, 
    -1.983852e-12, -1.986615e-12, -1.999547e-12, -1.99424e-12, -2.002686e-12, 
    -1.995098e-12, -1.996443e-12, -2.002961e-12, -1.995508e-12, 
    -2.011812e-12, -2.000758e-12, -2.021291e-12, -2.010251e-12, 
    -2.021983e-12, -2.019853e-12, -2.02338e-12, -2.026538e-12, -2.030512e-12, 
    -2.037845e-12, -2.036147e-12, -2.04228e-12, -1.979647e-12, -1.983403e-12, 
    -1.983073e-12, -1.987003e-12, -1.98991e-12, -1.99621e-12, -2.006316e-12, 
    -2.002516e-12, -2.009492e-12, -2.010893e-12, -2.000294e-12, 
    -2.006801e-12, -1.985916e-12, -1.98929e-12, -1.987282e-12, -1.979944e-12, 
    -2.003391e-12, -1.991357e-12, -2.013579e-12, -2.00706e-12, -2.026088e-12, 
    -2.016624e-12, -2.035212e-12, -2.043159e-12, -2.050639e-12, -2.05938e-12, 
    -1.985453e-12, -1.982901e-12, -1.98747e-12, -1.993792e-12, -1.999658e-12, 
    -2.007457e-12, -2.008256e-12, -2.009717e-12, -2.013502e-12, 
    -2.016684e-12, -2.010178e-12, -2.017481e-12, -1.990072e-12, 
    -2.004436e-12, -1.981936e-12, -1.98871e-12, -1.993419e-12, -1.991354e-12, 
    -2.002081e-12, -2.00461e-12, -2.014884e-12, -2.009573e-12, -2.041197e-12, 
    -2.027205e-12, -2.066036e-12, -2.055183e-12, -1.982009e-12, 
    -1.985444e-12, -1.997398e-12, -1.99171e-12, -2.007978e-12, -2.011983e-12, 
    -2.015238e-12, -2.0194e-12, -2.019849e-12, -2.022315e-12, -2.018274e-12, 
    -2.022155e-12, -2.007474e-12, -2.014035e-12, -1.996032e-12, 
    -2.000414e-12, -1.998398e-12, -1.996187e-12, -2.003011e-12, 
    -2.010281e-12, -2.010437e-12, -2.012768e-12, -2.019335e-12, 
    -2.008044e-12, -2.043002e-12, -2.021411e-12, -1.98919e-12, -1.995805e-12, 
    -1.996751e-12, -1.994188e-12, -2.011581e-12, -2.005279e-12, 
    -2.022255e-12, -2.017667e-12, -2.025184e-12, -2.021449e-12, 
    -2.020899e-12, -2.016101e-12, -2.013114e-12, -2.005568e-12, 
    -1.999428e-12, -1.99456e-12, -1.995692e-12, -2.001039e-12, -2.010726e-12, 
    -2.019889e-12, -2.017882e-12, -2.024613e-12, -2.006799e-12, 
    -2.014268e-12, -2.011381e-12, -2.018909e-12, -2.002415e-12, 
    -2.016459e-12, -1.998825e-12, -2.000371e-12, -2.005154e-12, 
    -2.014774e-12, -2.016904e-12, -2.019176e-12, -2.017774e-12, 
    -2.010971e-12, -2.009857e-12, -2.005037e-12, -2.003706e-12, 
    -2.000034e-12, -1.996994e-12, -1.999772e-12, -2.002689e-12, 
    -2.010975e-12, -2.018442e-12, -2.026583e-12, -2.028576e-12, 
    -2.038088e-12, -2.030344e-12, -2.043122e-12, -2.032257e-12, 
    -2.051066e-12, -2.017274e-12, -2.031939e-12, -2.005371e-12, 
    -2.008233e-12, -2.01341e-12, -2.025284e-12, -2.018874e-12, -2.02637e-12, 
    -2.009814e-12, -2.001224e-12, -1.999002e-12, -1.994855e-12, 
    -1.999097e-12, -1.998752e-12, -2.00281e-12, -2.001506e-12, -2.01125e-12, 
    -2.006016e-12, -2.020885e-12, -2.026311e-12, -2.041637e-12, 
    -2.051033e-12, -2.060598e-12, -2.064821e-12, -2.066106e-12, -2.066644e-12 ;

 SMINN_TO_SOIL2N_L3 =
  3.754954e-15, 3.765249e-15, 3.763249e-15, 3.771547e-15, 3.766946e-15, 
    3.772377e-15, 3.757043e-15, 3.765656e-15, 3.76016e-15, 3.755883e-15, 
    3.787629e-15, 3.771917e-15, 3.803946e-15, 3.793938e-15, 3.81907e-15, 
    3.802387e-15, 3.822431e-15, 3.818592e-15, 3.830152e-15, 3.826842e-15, 
    3.841607e-15, 3.831679e-15, 3.849259e-15, 3.839239e-15, 3.840806e-15, 
    3.831351e-15, 3.775084e-15, 3.785673e-15, 3.774455e-15, 3.775967e-15, 
    3.775289e-15, 3.76704e-15, 3.762878e-15, 3.754169e-15, 3.755751e-15, 
    3.762149e-15, 3.776646e-15, 3.771729e-15, 3.784124e-15, 3.783845e-15, 
    3.797629e-15, 3.791416e-15, 3.814564e-15, 3.80799e-15, 3.82698e-15, 
    3.822207e-15, 3.826755e-15, 3.825377e-15, 3.826773e-15, 3.819772e-15, 
    3.822771e-15, 3.81661e-15, 3.792579e-15, 3.799645e-15, 3.778557e-15, 
    3.765855e-15, 3.757421e-15, 3.75143e-15, 3.752277e-15, 3.753891e-15, 
    3.762186e-15, 3.769984e-15, 3.775923e-15, 3.779893e-15, 3.783805e-15, 
    3.795627e-15, 3.801889e-15, 3.815891e-15, 3.813368e-15, 3.817644e-15, 
    3.821732e-15, 3.828587e-15, 3.827459e-15, 3.830478e-15, 3.817533e-15, 
    3.826137e-15, 3.81193e-15, 3.815817e-15, 3.784855e-15, 3.773056e-15, 
    3.768027e-15, 3.763633e-15, 3.752928e-15, 3.760321e-15, 3.757407e-15, 
    3.764341e-15, 3.768744e-15, 3.766567e-15, 3.780002e-15, 3.77478e-15, 
    3.802259e-15, 3.790431e-15, 3.821255e-15, 3.813886e-15, 3.823021e-15, 
    3.818361e-15, 3.826343e-15, 3.81916e-15, 3.831603e-15, 3.834309e-15, 
    3.832459e-15, 3.839566e-15, 3.818761e-15, 3.826754e-15, 3.766506e-15, 
    3.766861e-15, 3.768516e-15, 3.761239e-15, 3.760794e-15, 3.754125e-15, 
    3.760061e-15, 3.762586e-15, 3.769001e-15, 3.772791e-15, 3.776394e-15, 
    3.784312e-15, 3.793148e-15, 3.805498e-15, 3.814364e-15, 3.820303e-15, 
    3.816662e-15, 3.819877e-15, 3.816283e-15, 3.814599e-15, 3.833294e-15, 
    3.822799e-15, 3.838545e-15, 3.837674e-15, 3.830549e-15, 3.837772e-15, 
    3.76711e-15, 3.765067e-15, 3.757967e-15, 3.763524e-15, 3.753399e-15, 
    3.759066e-15, 3.762322e-15, 3.774886e-15, 3.777648e-15, 3.780205e-15, 
    3.785256e-15, 3.791734e-15, 3.803089e-15, 3.812962e-15, 3.82197e-15, 
    3.82131e-15, 3.821542e-15, 3.823552e-15, 3.818571e-15, 3.82437e-15, 
    3.825342e-15, 3.822799e-15, 3.837558e-15, 3.833343e-15, 3.837656e-15, 
    3.834912e-15, 3.765731e-15, 3.76917e-15, 3.767312e-15, 3.770805e-15, 
    3.768343e-15, 3.779283e-15, 3.782561e-15, 3.797892e-15, 3.791605e-15, 
    3.801613e-15, 3.792623e-15, 3.794216e-15, 3.801934e-15, 3.79311e-15, 
    3.812415e-15, 3.799325e-15, 3.823631e-15, 3.810566e-15, 3.824449e-15, 
    3.821931e-15, 3.8261e-15, 3.829832e-15, 3.834527e-15, 3.843183e-15, 
    3.84118e-15, 3.848416e-15, 3.774295e-15, 3.778751e-15, 3.778361e-15, 
    3.783024e-15, 3.786471e-15, 3.793942e-15, 3.805912e-15, 3.801413e-15, 
    3.809674e-15, 3.811331e-15, 3.798781e-15, 3.806486e-15, 3.781734e-15, 
    3.785734e-15, 3.783354e-15, 3.774646e-15, 3.802447e-15, 3.788185e-15, 
    3.81451e-15, 3.806794e-15, 3.8293e-15, 3.81811e-15, 3.840076e-15, 
    3.849448e-15, 3.858272e-15, 3.868562e-15, 3.781184e-15, 3.778157e-15, 
    3.783579e-15, 3.791072e-15, 3.798027e-15, 3.807264e-15, 3.80821e-15, 
    3.809939e-15, 3.814419e-15, 3.818184e-15, 3.810483e-15, 3.819127e-15, 
    3.786656e-15, 3.803685e-15, 3.777011e-15, 3.785045e-15, 3.790632e-15, 
    3.788184e-15, 3.800899e-15, 3.803893e-15, 3.816052e-15, 3.80977e-15, 
    3.847133e-15, 3.830617e-15, 3.876398e-15, 3.863622e-15, 3.777099e-15, 
    3.781175e-15, 3.795348e-15, 3.788607e-15, 3.807882e-15, 3.812621e-15, 
    3.816474e-15, 3.821394e-15, 3.821927e-15, 3.82484e-15, 3.820064e-15, 
    3.824653e-15, 3.807284e-15, 3.815049e-15, 3.793731e-15, 3.798922e-15, 
    3.796536e-15, 3.793915e-15, 3.802e-15, 3.810604e-15, 3.810791e-15, 
    3.813549e-15, 3.821307e-15, 3.80796e-15, 3.849256e-15, 3.823763e-15, 
    3.785618e-15, 3.793458e-15, 3.794582e-15, 3.791545e-15, 3.812145e-15, 
    3.804685e-15, 3.82477e-15, 3.819346e-15, 3.828233e-15, 3.823817e-15, 
    3.823167e-15, 3.817494e-15, 3.81396e-15, 3.805026e-15, 3.797754e-15, 
    3.791986e-15, 3.793328e-15, 3.799663e-15, 3.811131e-15, 3.821973e-15, 
    3.819598e-15, 3.827558e-15, 3.806485e-15, 3.815324e-15, 3.811907e-15, 
    3.820815e-15, 3.801292e-15, 3.817907e-15, 3.797041e-15, 3.798872e-15, 
    3.804537e-15, 3.81592e-15, 3.818443e-15, 3.82113e-15, 3.819473e-15, 
    3.811423e-15, 3.810105e-15, 3.8044e-15, 3.802822e-15, 3.798474e-15, 
    3.794871e-15, 3.798162e-15, 3.801616e-15, 3.811428e-15, 3.82026e-15, 
    3.829885e-15, 3.83224e-15, 3.843463e-15, 3.834323e-15, 3.849397e-15, 
    3.836575e-15, 3.858766e-15, 3.818875e-15, 3.836205e-15, 3.804795e-15, 
    3.808184e-15, 3.814307e-15, 3.828346e-15, 3.820773e-15, 3.829631e-15, 
    3.810054e-15, 3.799879e-15, 3.79725e-15, 3.792336e-15, 3.797363e-15, 
    3.796954e-15, 3.801762e-15, 3.800218e-15, 3.811753e-15, 3.805558e-15, 
    3.82315e-15, 3.829562e-15, 3.847656e-15, 3.858732e-15, 3.870001e-15, 
    3.874971e-15, 3.876483e-15, 3.877115e-15 ;

 SMINN_TO_SOIL2N_S1 =
  -8.528931e-09, -8.566539e-09, -8.559229e-09, -8.589563e-09, -8.572736e-09, 
    -8.592599e-09, -8.536556e-09, -8.568032e-09, -8.547939e-09, 
    -8.532318e-09, -8.64843e-09, -8.590916e-09, -8.708187e-09, -8.671502e-09, 
    -8.763664e-09, -8.702478e-09, -8.776003e-09, -8.761901e-09, -8.80435e-09, 
    -8.792189e-09, -8.846483e-09, -8.809963e-09, -8.874632e-09, 
    -8.837763e-09, -8.843529e-09, -8.808758e-09, -8.602492e-09, 
    -8.641269e-09, -8.600194e-09, -8.605724e-09, -8.603243e-09, 
    -8.573084e-09, -8.557883e-09, -8.526058e-09, -8.531837e-09, 
    -8.555212e-09, -8.60821e-09, -8.590221e-09, -8.635564e-09, -8.63454e-09, 
    -8.685022e-09, -8.66226e-09, -8.747117e-09, -8.722998e-09, -8.792697e-09, 
    -8.775168e-09, -8.791874e-09, -8.786809e-09, -8.79194e-09, -8.766231e-09, 
    -8.777246e-09, -8.754625e-09, -8.666523e-09, -8.692413e-09, 
    -8.615197e-09, -8.568768e-09, -8.537937e-09, -8.516057e-09, 
    -8.519151e-09, -8.525046e-09, -8.555348e-09, -8.583842e-09, 
    -8.605555e-09, -8.620081e-09, -8.634393e-09, -8.677711e-09, 
    -8.700645e-09, -8.751993e-09, -8.742727e-09, -8.758425e-09, 
    -8.773424e-09, -8.798605e-09, -8.79446e-09, -8.805554e-09, -8.758012e-09, 
    -8.789607e-09, -8.73745e-09, -8.751715e-09, -8.638277e-09, -8.595074e-09, 
    -8.576706e-09, -8.560634e-09, -8.521528e-09, -8.548533e-09, 
    -8.537888e-09, -8.563216e-09, -8.57931e-09, -8.571351e-09, -8.620478e-09, 
    -8.601377e-09, -8.702004e-09, -8.658659e-09, -8.771675e-09, 
    -8.744629e-09, -8.778158e-09, -8.761049e-09, -8.790363e-09, 
    -8.763981e-09, -8.809684e-09, -8.819635e-09, -8.812834e-09, -8.83896e-09, 
    -8.762518e-09, -8.791873e-09, -8.571127e-09, -8.572425e-09, 
    -8.578473e-09, -8.551886e-09, -8.550261e-09, -8.525899e-09, 
    -8.547577e-09, -8.556808e-09, -8.580243e-09, -8.594105e-09, 
    -8.607282e-09, -8.636256e-09, -8.668615e-09, -8.713868e-09, 
    -8.746382e-09, -8.768177e-09, -8.754814e-09, -8.766612e-09, 
    -8.753423e-09, -8.747241e-09, -8.815905e-09, -8.777348e-09, 
    -8.835202e-09, -8.832001e-09, -8.805817e-09, -8.832362e-09, 
    -8.573337e-09, -8.565866e-09, -8.539929e-09, -8.560227e-09, 
    -8.523246e-09, -8.543945e-09, -8.555848e-09, -8.601775e-09, 
    -8.611869e-09, -8.621226e-09, -8.639707e-09, -8.663426e-09, 
    -8.705035e-09, -8.741242e-09, -8.774297e-09, -8.771875e-09, 
    -8.772727e-09, -8.780112e-09, -8.761821e-09, -8.783115e-09, 
    -8.786688e-09, -8.777344e-09, -8.831572e-09, -8.816079e-09, 
    -8.831933e-09, -8.821845e-09, -8.568295e-09, -8.580865e-09, 
    -8.574072e-09, -8.586845e-09, -8.577846e-09, -8.617859e-09, 
    -8.629856e-09, -8.685998e-09, -8.662958e-09, -8.699628e-09, 
    -8.666683e-09, -8.67252e-09, -8.700821e-09, -8.668464e-09, -8.739244e-09, 
    -8.691255e-09, -8.780399e-09, -8.73247e-09, -8.783402e-09, -8.774154e-09, 
    -8.789466e-09, -8.80318e-09, -8.820433e-09, -8.852267e-09, -8.844896e-09, 
    -8.871521e-09, -8.599605e-09, -8.615909e-09, -8.614474e-09, 
    -8.631538e-09, -8.644157e-09, -8.671512e-09, -8.715385e-09, 
    -8.698887e-09, -8.729176e-09, -8.735257e-09, -8.68924e-09, -8.717492e-09, 
    -8.626822e-09, -8.641469e-09, -8.632749e-09, -8.600891e-09, 
    -8.702687e-09, -8.650442e-09, -8.74692e-09, -8.718615e-09, -8.801224e-09, 
    -8.760138e-09, -8.840838e-09, -8.875336e-09, -8.90781e-09, -8.945757e-09, 
    -8.624808e-09, -8.61373e-09, -8.633568e-09, -8.661012e-09, -8.686482e-09, 
    -8.720341e-09, -8.723807e-09, -8.730149e-09, -8.746581e-09, 
    -8.760397e-09, -8.732154e-09, -8.763861e-09, -8.644863e-09, 
    -8.707222e-09, -8.609541e-09, -8.638952e-09, -8.659396e-09, 
    -8.650429e-09, -8.697001e-09, -8.707978e-09, -8.752584e-09, 
    -8.729526e-09, -8.86682e-09, -8.806074e-09, -8.974655e-09, -8.92754e-09, 
    -8.609859e-09, -8.624771e-09, -8.67667e-09, -8.651977e-09, -8.722602e-09, 
    -8.739987e-09, -8.754121e-09, -8.772187e-09, -8.774139e-09, 
    -8.784843e-09, -8.767302e-09, -8.78415e-09, -8.720414e-09, -8.748896e-09, 
    -8.67074e-09, -8.689761e-09, -8.681011e-09, -8.671412e-09, -8.701037e-09, 
    -8.732598e-09, -8.733275e-09, -8.743394e-09, -8.771909e-09, 
    -8.722889e-09, -8.874657e-09, -8.780922e-09, -8.641032e-09, 
    -8.669754e-09, -8.673858e-09, -8.662732e-09, -8.738244e-09, 
    -8.710883e-09, -8.784583e-09, -8.764664e-09, -8.797301e-09, 
    -8.781083e-09, -8.778696e-09, -8.757867e-09, -8.744899e-09, 
    -8.712137e-09, -8.685481e-09, -8.664346e-09, -8.669261e-09, 
    -8.692477e-09, -8.73453e-09, -8.774315e-09, -8.765599e-09, -8.794821e-09, 
    -8.717481e-09, -8.749909e-09, -8.737375e-09, -8.770058e-09, 
    -8.698448e-09, -8.759422e-09, -8.682862e-09, -8.689575e-09, 
    -8.710339e-09, -8.752107e-09, -8.761352e-09, -8.771218e-09, -8.76513e-09, 
    -8.735597e-09, -8.730759e-09, -8.709835e-09, -8.704057e-09, 
    -8.688114e-09, -8.674914e-09, -8.686974e-09, -8.699638e-09, -8.73561e-09, 
    -8.768028e-09, -8.803374e-09, -8.812026e-09, -8.853321e-09, 
    -8.819701e-09, -8.875178e-09, -8.828009e-09, -8.909667e-09, 
    -8.762958e-09, -8.826625e-09, -8.711285e-09, -8.723711e-09, 
    -8.746183e-09, -8.797732e-09, -8.769905e-09, -8.80245e-09, -8.73057e-09, 
    -8.693277e-09, -8.683632e-09, -8.665631e-09, -8.684043e-09, 
    -8.682545e-09, -8.700164e-09, -8.694503e-09, -8.736805e-09, 
    -8.714082e-09, -8.778636e-09, -8.802194e-09, -8.86873e-09, -8.90952e-09, 
    -8.951047e-09, -8.969381e-09, -8.974961e-09, -8.977294e-09 ;

 SMINN_TO_SOIL3N_S1 =
  -1.012121e-10, -1.016586e-10, -1.015718e-10, -1.019319e-10, -1.017321e-10, 
    -1.019679e-10, -1.013026e-10, -1.016763e-10, -1.014377e-10, 
    -1.012523e-10, -1.026307e-10, -1.01948e-10, -1.033402e-10, -1.029046e-10, 
    -1.039988e-10, -1.032724e-10, -1.041453e-10, -1.039779e-10, 
    -1.044818e-10, -1.043374e-10, -1.04982e-10, -1.045485e-10, -1.053162e-10, 
    -1.048785e-10, -1.04947e-10, -1.045341e-10, -1.020854e-10, -1.025457e-10, 
    -1.020581e-10, -1.021237e-10, -1.020943e-10, -1.017362e-10, 
    -1.015558e-10, -1.01178e-10, -1.012466e-10, -1.015241e-10, -1.021533e-10, 
    -1.019397e-10, -1.02478e-10, -1.024658e-10, -1.030651e-10, -1.027949e-10, 
    -1.038023e-10, -1.03516e-10, -1.043435e-10, -1.041354e-10, -1.043337e-10, 
    -1.042735e-10, -1.043345e-10, -1.040293e-10, -1.0416e-10, -1.038915e-10, 
    -1.028455e-10, -1.031529e-10, -1.022362e-10, -1.01685e-10, -1.01319e-10, 
    -1.010593e-10, -1.01096e-10, -1.01166e-10, -1.015257e-10, -1.01864e-10, 
    -1.021217e-10, -1.022942e-10, -1.024641e-10, -1.029783e-10, 
    -1.032506e-10, -1.038602e-10, -1.037502e-10, -1.039366e-10, 
    -1.041146e-10, -1.044136e-10, -1.043644e-10, -1.044961e-10, 
    -1.039317e-10, -1.043068e-10, -1.036876e-10, -1.038569e-10, 
    -1.025102e-10, -1.019973e-10, -1.017793e-10, -1.015885e-10, 
    -1.011242e-10, -1.014448e-10, -1.013184e-10, -1.016191e-10, 
    -1.018102e-10, -1.017157e-10, -1.022989e-10, -1.020721e-10, 
    -1.032667e-10, -1.027522e-10, -1.040939e-10, -1.037728e-10, 
    -1.041708e-10, -1.039677e-10, -1.043158e-10, -1.040025e-10, 
    -1.045451e-10, -1.046633e-10, -1.045825e-10, -1.048927e-10, 
    -1.039852e-10, -1.043337e-10, -1.01713e-10, -1.017284e-10, -1.018002e-10, 
    -1.014846e-10, -1.014653e-10, -1.011761e-10, -1.014334e-10, -1.01543e-10, 
    -1.018212e-10, -1.019858e-10, -1.021422e-10, -1.024862e-10, 
    -1.028704e-10, -1.034076e-10, -1.037936e-10, -1.040524e-10, 
    -1.038937e-10, -1.040338e-10, -1.038772e-10, -1.038038e-10, -1.04619e-10, 
    -1.041612e-10, -1.048481e-10, -1.048101e-10, -1.044992e-10, 
    -1.048144e-10, -1.017392e-10, -1.016506e-10, -1.013427e-10, 
    -1.015836e-10, -1.011446e-10, -1.013903e-10, -1.015316e-10, 
    -1.020769e-10, -1.021967e-10, -1.023078e-10, -1.025272e-10, 
    -1.028087e-10, -1.033027e-10, -1.037326e-10, -1.04125e-10, -1.040963e-10, 
    -1.041064e-10, -1.04194e-10, -1.039769e-10, -1.042297e-10, -1.042721e-10, 
    -1.041612e-10, -1.04805e-10, -1.046211e-10, -1.048093e-10, -1.046895e-10, 
    -1.016794e-10, -1.018286e-10, -1.01748e-10, -1.018996e-10, -1.017928e-10, 
    -1.022678e-10, -1.024102e-10, -1.030767e-10, -1.028032e-10, 
    -1.032385e-10, -1.028474e-10, -1.029167e-10, -1.032527e-10, 
    -1.028686e-10, -1.037089e-10, -1.031391e-10, -1.041974e-10, 
    -1.036284e-10, -1.042331e-10, -1.041233e-10, -1.043051e-10, 
    -1.044679e-10, -1.046727e-10, -1.050507e-10, -1.049632e-10, 
    -1.052793e-10, -1.020511e-10, -1.022447e-10, -1.022276e-10, 
    -1.024302e-10, -1.0258e-10, -1.029047e-10, -1.034256e-10, -1.032297e-10, 
    -1.035893e-10, -1.036615e-10, -1.031152e-10, -1.034506e-10, 
    -1.023742e-10, -1.025481e-10, -1.024446e-10, -1.020664e-10, 
    -1.032748e-10, -1.026546e-10, -1.038e-10, -1.03464e-10, -1.044447e-10, 
    -1.039569e-10, -1.04915e-10, -1.053246e-10, -1.057101e-10, -1.061607e-10, 
    -1.023503e-10, -1.022188e-10, -1.024543e-10, -1.027801e-10, 
    -1.030825e-10, -1.034844e-10, -1.035256e-10, -1.036009e-10, -1.03796e-10, 
    -1.0396e-10, -1.036247e-10, -1.040011e-10, -1.025884e-10, -1.033287e-10, 
    -1.02169e-10, -1.025182e-10, -1.027609e-10, -1.026545e-10, -1.032074e-10, 
    -1.033377e-10, -1.038672e-10, -1.035935e-10, -1.052235e-10, 
    -1.045023e-10, -1.065038e-10, -1.059444e-10, -1.021728e-10, 
    -1.023499e-10, -1.02966e-10, -1.026728e-10, -1.035113e-10, -1.037177e-10, 
    -1.038855e-10, -1.041e-10, -1.041231e-10, -1.042502e-10, -1.04042e-10, 
    -1.04242e-10, -1.034853e-10, -1.038234e-10, -1.028956e-10, -1.031214e-10, 
    -1.030175e-10, -1.029036e-10, -1.032553e-10, -1.0363e-10, -1.03638e-10, 
    -1.037581e-10, -1.040967e-10, -1.035147e-10, -1.053165e-10, 
    -1.042037e-10, -1.025429e-10, -1.028839e-10, -1.029326e-10, 
    -1.028005e-10, -1.03697e-10, -1.033722e-10, -1.042471e-10, -1.040106e-10, 
    -1.043981e-10, -1.042056e-10, -1.041772e-10, -1.0393e-10, -1.03776e-10, 
    -1.03387e-10, -1.030706e-10, -1.028197e-10, -1.02878e-10, -1.031536e-10, 
    -1.036529e-10, -1.041252e-10, -1.040217e-10, -1.043687e-10, 
    -1.034505e-10, -1.038355e-10, -1.036867e-10, -1.040747e-10, 
    -1.032245e-10, -1.039484e-10, -1.030395e-10, -1.031192e-10, 
    -1.033657e-10, -1.038616e-10, -1.039713e-10, -1.040885e-10, 
    -1.040162e-10, -1.036656e-10, -1.036081e-10, -1.033597e-10, 
    -1.032911e-10, -1.031018e-10, -1.029451e-10, -1.030883e-10, 
    -1.032387e-10, -1.036657e-10, -1.040506e-10, -1.044702e-10, 
    -1.045729e-10, -1.050632e-10, -1.046641e-10, -1.053227e-10, 
    -1.047627e-10, -1.057322e-10, -1.039904e-10, -1.047463e-10, 
    -1.033769e-10, -1.035244e-10, -1.037912e-10, -1.044032e-10, 
    -1.040729e-10, -1.044593e-10, -1.036059e-10, -1.031631e-10, 
    -1.030486e-10, -1.028349e-10, -1.030535e-10, -1.030357e-10, 
    -1.032449e-10, -1.031777e-10, -1.036799e-10, -1.034101e-10, 
    -1.041765e-10, -1.044562e-10, -1.052462e-10, -1.057304e-10, 
    -1.062235e-10, -1.064411e-10, -1.065074e-10, -1.065351e-10 ;

 SMINN_TO_SOIL3N_S2 =
  -8.394119e-12, -8.431162e-12, -8.423961e-12, -8.453839e-12, -8.437267e-12, 
    -8.45683e-12, -8.40163e-12, -8.432632e-12, -8.412842e-12, -8.397455e-12, 
    -8.511824e-12, -8.455173e-12, -8.570683e-12, -8.534548e-12, 
    -8.625329e-12, -8.565059e-12, -8.637482e-12, -8.623592e-12, 
    -8.665404e-12, -8.653426e-12, -8.706905e-12, -8.670933e-12, 
    -8.734632e-12, -8.698316e-12, -8.703995e-12, -8.669746e-12, 
    -8.466576e-12, -8.50477e-12, -8.464312e-12, -8.469758e-12, -8.467315e-12, 
    -8.437608e-12, -8.422637e-12, -8.391289e-12, -8.39698e-12, -8.420005e-12, 
    -8.472207e-12, -8.454488e-12, -8.49915e-12, -8.498141e-12, -8.547866e-12, 
    -8.525446e-12, -8.609029e-12, -8.585273e-12, -8.653926e-12, 
    -8.636659e-12, -8.653115e-12, -8.648125e-12, -8.65318e-12, -8.627856e-12, 
    -8.638706e-12, -8.616424e-12, -8.529645e-12, -8.555146e-12, 
    -8.479089e-12, -8.433357e-12, -8.402989e-12, -8.381439e-12, 
    -8.384485e-12, -8.390293e-12, -8.42014e-12, -8.448205e-12, -8.469592e-12, 
    -8.483899e-12, -8.497997e-12, -8.540665e-12, -8.563253e-12, 
    -8.613832e-12, -8.604705e-12, -8.620168e-12, -8.634942e-12, 
    -8.659745e-12, -8.655662e-12, -8.66659e-12, -8.619761e-12, -8.650882e-12, 
    -8.599507e-12, -8.613558e-12, -8.501823e-12, -8.459269e-12, 
    -8.441177e-12, -8.425345e-12, -8.386828e-12, -8.413426e-12, 
    -8.402941e-12, -8.427889e-12, -8.44374e-12, -8.435901e-12, -8.484291e-12, 
    -8.465477e-12, -8.564593e-12, -8.521898e-12, -8.633218e-12, 
    -8.606579e-12, -8.639604e-12, -8.622753e-12, -8.651626e-12, -8.62564e-12, 
    -8.670657e-12, -8.680459e-12, -8.67376e-12, -8.699495e-12, -8.624199e-12, 
    -8.653114e-12, -8.435681e-12, -8.436959e-12, -8.442917e-12, -8.41673e-12, 
    -8.415128e-12, -8.391132e-12, -8.412484e-12, -8.421577e-12, -8.44466e-12, 
    -8.458314e-12, -8.471293e-12, -8.499832e-12, -8.531705e-12, 
    -8.576279e-12, -8.608306e-12, -8.629774e-12, -8.61661e-12, -8.628232e-12, 
    -8.61524e-12, -8.609151e-12, -8.676786e-12, -8.638807e-12, -8.695793e-12, 
    -8.69264e-12, -8.666849e-12, -8.692995e-12, -8.437857e-12, -8.430499e-12, 
    -8.404952e-12, -8.424945e-12, -8.38852e-12, -8.408908e-12, -8.420631e-12, 
    -8.465869e-12, -8.47581e-12, -8.485027e-12, -8.503231e-12, -8.526593e-12, 
    -8.567579e-12, -8.603242e-12, -8.635801e-12, -8.633416e-12, 
    -8.634256e-12, -8.641528e-12, -8.623512e-12, -8.644486e-12, 
    -8.648006e-12, -8.638803e-12, -8.692218e-12, -8.676958e-12, 
    -8.692574e-12, -8.682637e-12, -8.432892e-12, -8.445272e-12, 
    -8.438582e-12, -8.451163e-12, -8.442299e-12, -8.481711e-12, 
    -8.493528e-12, -8.548827e-12, -8.526133e-12, -8.562252e-12, 
    -8.529803e-12, -8.535552e-12, -8.563428e-12, -8.531557e-12, 
    -8.601274e-12, -8.554005e-12, -8.641811e-12, -8.594602e-12, -8.64477e-12, 
    -8.635661e-12, -8.650743e-12, -8.664251e-12, -8.681246e-12, 
    -8.712604e-12, -8.705342e-12, -8.731568e-12, -8.463731e-12, 
    -8.479791e-12, -8.478378e-12, -8.495185e-12, -8.507615e-12, 
    -8.534558e-12, -8.577773e-12, -8.561522e-12, -8.591358e-12, 
    -8.597347e-12, -8.552021e-12, -8.579849e-12, -8.490539e-12, 
    -8.504966e-12, -8.496377e-12, -8.464998e-12, -8.565266e-12, 
    -8.513805e-12, -8.608835e-12, -8.580955e-12, -8.662324e-12, 
    -8.621856e-12, -8.701345e-12, -8.735325e-12, -8.767314e-12, 
    -8.804691e-12, -8.488556e-12, -8.477644e-12, -8.497184e-12, 
    -8.524217e-12, -8.549304e-12, -8.582655e-12, -8.586068e-12, 
    -8.592316e-12, -8.608502e-12, -8.62211e-12, -8.59429e-12, -8.625521e-12, 
    -8.50831e-12, -8.569733e-12, -8.473518e-12, -8.502487e-12, -8.522624e-12, 
    -8.513791e-12, -8.559665e-12, -8.570478e-12, -8.614415e-12, 
    -8.591702e-12, -8.726938e-12, -8.667103e-12, -8.833156e-12, 
    -8.786747e-12, -8.473831e-12, -8.48852e-12, -8.539639e-12, -8.515316e-12, 
    -8.584882e-12, -8.602006e-12, -8.615928e-12, -8.633723e-12, 
    -8.635646e-12, -8.64619e-12, -8.628912e-12, -8.645507e-12, -8.582727e-12, 
    -8.610781e-12, -8.533798e-12, -8.552534e-12, -8.543915e-12, -8.53446e-12, 
    -8.56364e-12, -8.594728e-12, -8.595394e-12, -8.605363e-12, -8.63345e-12, 
    -8.585165e-12, -8.734656e-12, -8.642326e-12, -8.504536e-12, 
    -8.532826e-12, -8.53687e-12, -8.52591e-12, -8.60029e-12, -8.573338e-12, 
    -8.645933e-12, -8.626312e-12, -8.65846e-12, -8.642485e-12, -8.640135e-12, 
    -8.619618e-12, -8.606844e-12, -8.574573e-12, -8.548318e-12, -8.5275e-12, 
    -8.532341e-12, -8.555209e-12, -8.59663e-12, -8.635819e-12, -8.627234e-12, 
    -8.656017e-12, -8.579838e-12, -8.61178e-12, -8.599433e-12, -8.631627e-12, 
    -8.56109e-12, -8.621149e-12, -8.545739e-12, -8.552351e-12, -8.572803e-12, 
    -8.613945e-12, -8.62305e-12, -8.632769e-12, -8.626772e-12, -8.597682e-12, 
    -8.592917e-12, -8.572306e-12, -8.566614e-12, -8.550912e-12, -8.53791e-12, 
    -8.549788e-12, -8.562263e-12, -8.597695e-12, -8.629627e-12, 
    -8.664442e-12, -8.672964e-12, -8.713641e-12, -8.680525e-12, 
    -8.735171e-12, -8.688708e-12, -8.769142e-12, -8.624633e-12, 
    -8.687345e-12, -8.573735e-12, -8.585974e-12, -8.608109e-12, 
    -8.658885e-12, -8.631475e-12, -8.663533e-12, -8.592731e-12, 
    -8.555997e-12, -8.546496e-12, -8.528765e-12, -8.546901e-12, 
    -8.545427e-12, -8.562781e-12, -8.557204e-12, -8.598872e-12, 
    -8.576489e-12, -8.640076e-12, -8.66328e-12, -8.728819e-12, -8.768998e-12, 
    -8.809903e-12, -8.827962e-12, -8.833458e-12, -8.835756e-12 ;

 SMIN_NH4 =
  0.0004350498, 0.0004368826, 0.0004365262, 0.0004380044, 0.0004371844, 
    0.0004381522, 0.0004354211, 0.0004369549, 0.0004359757, 0.0004352143, 
    0.0004408726, 0.00043807, 0.0004437841, 0.0004419966, 0.0004464868, 
    0.0004435058, 0.0004470879, 0.0004464008, 0.0004484687, 0.0004478762, 
    0.000450521, 0.000448742, 0.000451892, 0.0004500961, 0.0004503769, 
    0.000448683, 0.0004386345, 0.000440524, 0.0004385223, 0.0004387918, 
    0.0004386709, 0.0004372011, 0.0004364603, 0.0004349092, 0.0004351908, 
    0.00043633, 0.0004389126, 0.0004380359, 0.0004402453, 0.0004401955, 
    0.0004426551, 0.0004415461, 0.0004456804, 0.0004445053, 0.0004479008, 
    0.0004470468, 0.0004478606, 0.0004476138, 0.0004478637, 0.0004466113, 
    0.0004471477, 0.0004460457, 0.0004417544, 0.0004430158, 0.0004392533, 
    0.0004369908, 0.0004354881, 0.0004344218, 0.0004345725, 0.0004348598, 
    0.0004363365, 0.000437725, 0.0004387831, 0.0004394908, 0.0004401881, 
    0.0004422989, 0.0004434162, 0.0004459178, 0.0004454664, 0.0004462311, 
    0.0004469618, 0.0004481884, 0.0004479865, 0.0004485268, 0.0004462107, 
    0.0004477499, 0.0004452088, 0.0004459038, 0.000440378, 0.0004382726, 
    0.0004373775, 0.0004365942, 0.0004346884, 0.0004360044, 0.0004354855, 
    0.0004367198, 0.0004375041, 0.0004371161, 0.0004395101, 0.0004385793, 
    0.0004434823, 0.0004413704, 0.0004468766, 0.000445559, 0.0004471923, 
    0.0004463588, 0.0004477868, 0.0004465015, 0.0004487279, 0.0004492127, 
    0.0004488813, 0.000450154, 0.0004464299, 0.00044786, 0.0004371055, 
    0.0004371688, 0.0004374635, 0.0004361678, 0.0004360885, 0.0004349012, 
    0.0004359575, 0.0004364074, 0.0004375494, 0.0004382248, 0.0004388669, 
    0.0004402787, 0.0004418554, 0.0004440602, 0.0004456443, 0.000446706, 
    0.0004460549, 0.0004466297, 0.0004459871, 0.0004456858, 0.0004490309, 
    0.0004471525, 0.0004499707, 0.0004498148, 0.0004485393, 0.0004498322, 
    0.0004372131, 0.000436849, 0.000435585, 0.0004365741, 0.0004347718, 
    0.0004357806, 0.0004363605, 0.0004385986, 0.0004390903, 0.0004395463, 
    0.0004404468, 0.0004416024, 0.0004436298, 0.0004453937, 0.0004470041, 
    0.000446886, 0.0004469275, 0.0004472872, 0.0004463961, 0.0004474334, 
    0.0004476074, 0.0004471522, 0.0004497938, 0.0004490391, 0.0004498113, 
    0.0004493198, 0.0004369673, 0.0004375798, 0.0004372487, 0.0004378711, 
    0.0004374325, 0.0004393823, 0.0004399669, 0.0004427023, 0.0004415796, 
    0.0004433664, 0.000441761, 0.0004420455, 0.0004434244, 0.0004418477, 
    0.0004452962, 0.000442958, 0.0004473011, 0.000444966, 0.0004474473, 
    0.0004469967, 0.0004477426, 0.0004484106, 0.000449251, 0.0004508018, 
    0.0004504426, 0.0004517395, 0.0004384929, 0.0004392873, 0.0004392174, 
    0.0004400488, 0.0004406636, 0.0004419965, 0.0004441341, 0.0004433302, 
    0.0004448058, 0.0004451021, 0.00044286, 0.0004442365, 0.0004398185, 
    0.0004405321, 0.0004401072, 0.0004385547, 0.0004435148, 0.0004409692, 
    0.0004456698, 0.0004442907, 0.0004483152, 0.0004463137, 0.0004502448, 
    0.0004519253, 0.000453507, 0.0004553551, 0.0004397209, 0.000439181, 
    0.0004401476, 0.0004414849, 0.0004427258, 0.0004443755, 0.0004445442, 
    0.0004448532, 0.0004456537, 0.0004463268, 0.0004449507, 0.0004464953, 
    0.0004406975, 0.0004437358, 0.0004389761, 0.0004404093, 0.0004414053, 
    0.0004409684, 0.0004432376, 0.0004437723, 0.0004459455, 0.0004448221, 
    0.0004515103, 0.0004485513, 0.0004567624, 0.0004544677, 0.0004389923, 
    0.0004397189, 0.0004422477, 0.0004410445, 0.0004444855, 0.0004453325, 
    0.000446021, 0.0004469011, 0.0004469961, 0.0004475176, 0.0004466629, 
    0.0004474837, 0.0004443784, 0.0004457661, 0.0004419581, 0.0004428848, 
    0.0004424584, 0.0004419906, 0.000443434, 0.0004449718, 0.0004450046, 
    0.0004454976, 0.0004468868, 0.0004444984, 0.0004518919, 0.0004473257, 
    0.0004405112, 0.0004419106, 0.0004421105, 0.0004415684, 0.0004452474, 
    0.0004439143, 0.0004475049, 0.0004465344, 0.0004481243, 0.0004473342, 
    0.0004472179, 0.0004462031, 0.0004455712, 0.000443975, 0.0004426762, 
    0.0004416464, 0.0004418857, 0.0004430169, 0.0004450657, 0.000447004, 
    0.0004465793, 0.0004480028, 0.0004442348, 0.0004458148, 0.000445204, 
    0.0004467963, 0.0004433086, 0.0004462793, 0.0004425491, 0.0004428761, 
    0.0004438877, 0.0004459227, 0.0004463729, 0.0004468536, 0.0004465569, 
    0.0004451181, 0.0004448823, 0.0004438628, 0.0004435812, 0.0004428044, 
    0.0004421611, 0.0004427487, 0.0004433657, 0.0004451183, 0.0004466976, 
    0.0004484195, 0.0004488409, 0.0004508524, 0.0004492147, 0.000451917, 
    0.0004496193, 0.0004535968, 0.0004464514, 0.000449553, 0.0004439338, 
    0.0004445391, 0.000445634, 0.0004481452, 0.0004467895, 0.000448375, 
    0.0004448731, 0.000443056, 0.0004425859, 0.0004417089, 0.0004426059, 
    0.0004425329, 0.0004433913, 0.0004431154, 0.0004451764, 0.0004440693, 
    0.0004472142, 0.0004483619, 0.0004516029, 0.0004535897, 0.0004556122, 
    0.000456505, 0.0004567768, 0.0004568903 ;

 SMIN_NH4_vr =
  0.002842416, 0.00284735, 0.002846385, 0.002850361, 0.002848153, 0.00285075, 
    0.002843402, 0.002847523, 0.002844889, 0.002842835, 0.00285804, 
    0.002850514, 0.002865857, 0.002861057, 0.002873096, 0.002865101, 
    0.002874704, 0.00287286, 0.002878399, 0.002876807, 0.002883879, 
    0.002879123, 0.002887541, 0.002882739, 0.002883486, 0.00287895, 
    0.002852054, 0.002857126, 0.002851746, 0.002852471, 0.002852143, 
    0.002848184, 0.002846188, 0.002842012, 0.002842766, 0.002845831, 
    0.002852774, 0.002850413, 0.002856349, 0.002856215, 0.002862813, 
    0.002859837, 0.002870926, 0.002867771, 0.00287687, 0.002874577, 
    0.002876756, 0.002876091, 0.002876756, 0.002873401, 0.002874832, 
    0.00287188, 0.002860431, 0.002863812, 0.002853706, 0.002847614, 
    0.002843569, 0.0028407, 0.002841099, 0.002841873, 0.002845843, 
    0.002849575, 0.002852419, 0.002854317, 0.002856187, 0.002861851, 
    0.002864848, 0.002871554, 0.002870345, 0.002872388, 0.002874346, 
    0.002877627, 0.002877085, 0.002878527, 0.002872319, 0.002876443, 
    0.002869628, 0.002871491, 0.002856719, 0.002851063, 0.002848651, 
    0.002846542, 0.002841409, 0.002844951, 0.002843551, 0.002846869, 
    0.002848977, 0.00284793, 0.002854365, 0.002851859, 0.002865021, 
    0.002859354, 0.002874122, 0.002870586, 0.002874959, 0.002872727, 
    0.002876545, 0.002873104, 0.00287906, 0.002880357, 0.002879464, 
    0.002882872, 0.002872893, 0.002876724, 0.002847919, 0.002848089, 
    0.002848878, 0.002845386, 0.002845172, 0.002841972, 0.002844812, 
    0.002846022, 0.002849092, 0.002850903, 0.002852625, 0.002856421, 
    0.00286065, 0.002866563, 0.002870811, 0.002873653, 0.002871907, 
    0.002873442, 0.002871718, 0.002870907, 0.002879862, 0.002874833, 
    0.002882373, 0.002881956, 0.002878537, 0.002881994, 0.002848202, 
    0.002847219, 0.002843815, 0.002846473, 0.002841618, 0.002844333, 
    0.002845889, 0.002851905, 0.002853225, 0.00285445, 0.002856866, 
    0.002859965, 0.002865405, 0.002870132, 0.002874448, 0.002874127, 
    0.002874237, 0.002875195, 0.002872807, 0.002875581, 0.002876043, 
    0.002874825, 0.002881891, 0.002879872, 0.002881935, 0.002880615, 
    0.002847534, 0.002849176, 0.002848282, 0.002849956, 0.00284877, 
    0.002854011, 0.002855578, 0.00286292, 0.002859904, 0.0028647, 
    0.002860385, 0.002861149, 0.002864842, 0.002860611, 0.00286986, 
    0.002863582, 0.002875229, 0.002868962, 0.002875615, 0.002874404, 
    0.002876398, 0.002878187, 0.002880431, 0.002884579, 0.002883612, 
    0.002887082, 0.002851628, 0.002853758, 0.002853571, 0.0028558, 
    0.002857447, 0.002861028, 0.00286676, 0.002864599, 0.002868555, 
    0.002869349, 0.002863328, 0.002867021, 0.002855155, 0.002857067, 
    0.002855926, 0.002851748, 0.002865068, 0.002858229, 0.002870844, 
    0.002867141, 0.002877923, 0.00287256, 0.002883082, 0.002887573, 
    0.0028918, 0.002896726, 0.002854921, 0.002853466, 0.00285606, 0.00285965, 
    0.002862977, 0.002867404, 0.002867854, 0.002868677, 0.00287082, 
    0.002872625, 0.00286893, 0.002873068, 0.002857504, 0.002865661, 
    0.002852875, 0.002856725, 0.002859395, 0.002858224, 0.002864313, 
    0.002865743, 0.002871565, 0.002868556, 0.002886454, 0.002878539, 
    0.002900477, 0.002894353, 0.002852955, 0.002854904, 0.00286169, 
    0.002858461, 0.002867691, 0.002869963, 0.002871803, 0.002874161, 
    0.00287441, 0.002875807, 0.002873511, 0.002875711, 0.00286738, 
    0.002871102, 0.002860882, 0.002863364, 0.00286222, 0.002860959, 
    0.002864829, 0.002868952, 0.002869039, 0.002870355, 0.002874069, 
    0.002867671, 0.002887459, 0.002875236, 0.002857029, 0.00286078, 
    0.002861315, 0.002859861, 0.002869726, 0.002866151, 0.002875773, 
    0.002873169, 0.002877424, 0.002875308, 0.00287499, 0.002872271, 
    0.002870571, 0.00286629, 0.002862798, 0.002860036, 0.002860671, 
    0.002863707, 0.002869196, 0.002874393, 0.002873251, 0.002877061, 
    0.002866958, 0.002871194, 0.00286955, 0.00287382, 0.002864529, 
    0.002872489, 0.002862488, 0.002863361, 0.002866071, 0.002871526, 
    0.00287273, 0.002874017, 0.002873217, 0.002869359, 0.002868724, 
    0.002865985, 0.002865225, 0.002863142, 0.002861409, 0.002862986, 
    0.002864635, 0.002869337, 0.002873566, 0.002878174, 0.002879302, 
    0.002884674, 0.002880292, 0.002887511, 0.002881363, 0.002891996, 
    0.002872945, 0.002881251, 0.002866196, 0.002867815, 0.002870747, 
    0.00287747, 0.002873838, 0.002878083, 0.002868697, 0.002863816, 
    0.002862553, 0.002860199, 0.002862601, 0.002862405, 0.002864706, 
    0.002863961, 0.002869484, 0.002866516, 0.00287494, 0.002878013, 
    0.002886682, 0.002891985, 0.002897387, 0.002899764, 0.002900488, 
    0.002900787,
  0.001592185, 0.001598216, 0.001597044, 0.001601904, 0.001599209, 
    0.001602391, 0.001593409, 0.001598454, 0.001595234, 0.001592729, 
    0.001611324, 0.001602121, 0.001620875, 0.001615015, 0.001629726, 
    0.001619962, 0.001631693, 0.001629446, 0.00163621, 0.001634273, 
    0.001642913, 0.001637104, 0.001647389, 0.001641527, 0.001642444, 
    0.001636912, 0.001603976, 0.001610178, 0.001603608, 0.001604493, 
    0.001604096, 0.001599264, 0.001596827, 0.001591725, 0.001592652, 
    0.0015964, 0.001604891, 0.001602011, 0.001609269, 0.001609105, 
    0.001617176, 0.001613538, 0.001627088, 0.00162324, 0.001634354, 
    0.001631561, 0.001634222, 0.001633416, 0.001634233, 0.001630136, 
    0.001631891, 0.001628286, 0.001614219, 0.001618356, 0.001606009, 
    0.001598571, 0.00159363, 0.00159012, 0.001590616, 0.001591562, 
    0.001596422, 0.001600989, 0.001604466, 0.001606792, 0.001609082, 
    0.001616005, 0.00161967, 0.001627865, 0.001626388, 0.001628891, 
    0.001631283, 0.001635294, 0.001634634, 0.001636401, 0.001628826, 
    0.001633861, 0.001625546, 0.001627822, 0.001609699, 0.001602788, 
    0.001599844, 0.001597269, 0.001590998, 0.001595329, 0.001593622, 
    0.001597684, 0.001600263, 0.001598987, 0.001606855, 0.001603797, 
    0.001619887, 0.001612962, 0.001631004, 0.001626692, 0.001632037, 
    0.00162931, 0.001633981, 0.001629778, 0.001637059, 0.001638642, 
    0.00163756, 0.001641718, 0.001629544, 0.001634222, 0.001598952, 
    0.001599159, 0.001600129, 0.001595867, 0.001595606, 0.001591699, 
    0.001595176, 0.001596656, 0.001600413, 0.001602633, 0.001604743, 
    0.00160938, 0.001614553, 0.001621782, 0.001626971, 0.001630447, 
    0.001628316, 0.001630197, 0.001628094, 0.001627108, 0.001638049, 
    0.001631908, 0.00164112, 0.001640611, 0.001636443, 0.001640668, 
    0.001599306, 0.001598109, 0.00159395, 0.001597205, 0.001591274, 
    0.001594594, 0.001596501, 0.00160386, 0.001605477, 0.001606974, 
    0.001609932, 0.001613725, 0.001620372, 0.001626151, 0.001631422, 
    0.001631036, 0.001631172, 0.001632348, 0.001629433, 0.001632827, 
    0.001633396, 0.001631907, 0.001640543, 0.001638077, 0.0016406, 
    0.001638995, 0.001598498, 0.001600512, 0.001599424, 0.00160147, 
    0.001600028, 0.001606435, 0.001608354, 0.001617331, 0.00161365, 
    0.001619508, 0.001614245, 0.001615178, 0.001619697, 0.00161453, 
    0.001625831, 0.00161817, 0.001632394, 0.00162475, 0.001632873, 
    0.001631399, 0.001633839, 0.001636023, 0.00163877, 0.001643834, 
    0.001642662, 0.001646895, 0.001603513, 0.001606123, 0.001605894, 
    0.001608625, 0.001610643, 0.001615017, 0.001622025, 0.001619391, 
    0.001624226, 0.001625196, 0.00161785, 0.001622361, 0.00160787, 
    0.001610212, 0.001608818, 0.001603719, 0.001619997, 0.001611648, 
    0.001627057, 0.001622541, 0.001635711, 0.001629164, 0.001642016, 
    0.0016475, 0.00165266, 0.00165868, 0.001607548, 0.001605775, 0.00160895, 
    0.001613338, 0.001617409, 0.001622816, 0.001623369, 0.001624381, 
    0.001627003, 0.001629206, 0.0016247, 0.001629758, 0.001610753, 
    0.001620721, 0.001605104, 0.001609809, 0.00161308, 0.001611646, 
    0.00161909, 0.001620843, 0.00162796, 0.001624282, 0.001646146, 
    0.001636483, 0.001663262, 0.00165579, 0.001605155, 0.001607542, 
    0.001615841, 0.001611894, 0.001623177, 0.001625951, 0.001628206, 
    0.001631085, 0.001631397, 0.001633102, 0.001630307, 0.001632992, 
    0.001622827, 0.001627372, 0.001614894, 0.001617933, 0.001616535, 
    0.001615001, 0.001619734, 0.001624771, 0.00162488, 0.001626494, 
    0.001631037, 0.001623223, 0.001647389, 0.001632474, 0.001610144, 
    0.001614735, 0.001615392, 0.001613614, 0.001625673, 0.001621306, 
    0.001633061, 0.001629886, 0.001635087, 0.001632503, 0.001632123, 
    0.001628803, 0.001626735, 0.001621506, 0.001617249, 0.001613872, 
    0.001614658, 0.001618367, 0.001625079, 0.001631424, 0.001630035, 
    0.001634692, 0.00162236, 0.001627533, 0.001625534, 0.001630746, 
    0.00161932, 0.001629047, 0.001616831, 0.001617904, 0.001621219, 
    0.001627883, 0.001629358, 0.001630931, 0.001629961, 0.00162525, 
    0.001624479, 0.001621139, 0.001620216, 0.00161767, 0.001615561, 
    0.001617488, 0.00161951, 0.001625253, 0.001630422, 0.001636054, 
    0.001637432, 0.001643999, 0.001638651, 0.001647472, 0.001639971, 
    0.001652951, 0.001629612, 0.001639753, 0.001621371, 0.001623354, 
    0.001626938, 0.001635154, 0.001630722, 0.001635906, 0.001624448, 
    0.001618494, 0.001616954, 0.001614077, 0.00161702, 0.001616781, 
    0.001619595, 0.001618691, 0.001625443, 0.001621817, 0.001632113, 
    0.001635865, 0.001646451, 0.00165293, 0.001659521, 0.001662427, 
    0.001663311, 0.001663681,
  0.001500654, 0.00150729, 0.001506001, 0.00151135, 0.001508383, 0.001511885, 
    0.001502, 0.001507553, 0.001504009, 0.001501253, 0.001521721, 
    0.001511588, 0.001532239, 0.001525784, 0.001541993, 0.001531235, 
    0.001544161, 0.001541683, 0.001549139, 0.001547004, 0.001556532, 
    0.001550125, 0.001561469, 0.001555003, 0.001556014, 0.001549913, 
    0.001513629, 0.00152046, 0.001513224, 0.001514198, 0.001513761, 
    0.001508444, 0.001505763, 0.001500148, 0.001501168, 0.001505292, 
    0.001514637, 0.001511466, 0.001519457, 0.001519276, 0.001528164, 
    0.001524158, 0.001539085, 0.001534845, 0.001547093, 0.001544014, 
    0.001546948, 0.001546059, 0.00154696, 0.001542444, 0.001544379, 
    0.001540405, 0.001524908, 0.001529465, 0.001515868, 0.001507682, 
    0.001502244, 0.001498382, 0.001498928, 0.001499969, 0.001505316, 
    0.001510341, 0.001514169, 0.001516729, 0.00151925, 0.001526877, 
    0.001530912, 0.001539942, 0.001538313, 0.001541072, 0.001543708, 
    0.00154813, 0.001547403, 0.00154935, 0.001541, 0.00154655, 0.001537386, 
    0.001539893, 0.001519933, 0.001512322, 0.001509083, 0.001506248, 
    0.001499348, 0.001504114, 0.001502235, 0.001506704, 0.001509542, 
    0.001508139, 0.001516799, 0.001513433, 0.001531152, 0.001523523, 
    0.0015434, 0.001538648, 0.001544539, 0.001541534, 0.001546683, 
    0.001542049, 0.001550075, 0.001551822, 0.001550628, 0.001555213, 
    0.001541792, 0.001546948, 0.001508099, 0.001508328, 0.001509395, 
    0.001504705, 0.001504418, 0.00150012, 0.001503945, 0.001505573, 
    0.001509707, 0.001512151, 0.001514473, 0.001519578, 0.001525276, 
    0.001533239, 0.001538956, 0.001542786, 0.001540438, 0.001542511, 
    0.001540193, 0.001539107, 0.001551167, 0.001544397, 0.001554554, 
    0.001553992, 0.001549397, 0.001554056, 0.001508489, 0.001507172, 
    0.001502596, 0.001506177, 0.001499651, 0.001503304, 0.001505404, 
    0.001513502, 0.001515282, 0.00151693, 0.001520186, 0.001524363, 
    0.001531685, 0.001538052, 0.001543861, 0.001543436, 0.001543586, 
    0.001544883, 0.001541669, 0.00154541, 0.001546037, 0.001544396, 
    0.001553917, 0.001551198, 0.00155398, 0.00155221, 0.0015076, 0.001509816, 
    0.001508619, 0.001510871, 0.001509284, 0.001516337, 0.00151845, 
    0.001528335, 0.00152428, 0.001530734, 0.001524936, 0.001525964, 
    0.001530943, 0.00152525, 0.001537701, 0.00152926, 0.001544933, 
    0.001536509, 0.00154546, 0.001543836, 0.001546526, 0.001548933, 
    0.001551962, 0.001557547, 0.001556255, 0.001560924, 0.00151312, 
    0.001515993, 0.001515741, 0.001518747, 0.00152097, 0.001525786, 
    0.001533506, 0.001530604, 0.001535931, 0.001537, 0.001528907, 
    0.001533876, 0.001517916, 0.001520496, 0.00151896, 0.001513347, 
    0.001531272, 0.001522076, 0.00153905, 0.001534074, 0.00154859, 
    0.001541373, 0.001555543, 0.001561592, 0.001567284, 0.001573929, 
    0.001517562, 0.00151561, 0.001519105, 0.001523938, 0.001528421, 
    0.001534377, 0.001534987, 0.001536102, 0.001538991, 0.001541419, 
    0.001536454, 0.001542028, 0.001521093, 0.00153207, 0.001514871, 
    0.001520053, 0.001523653, 0.001522074, 0.001530272, 0.001532203, 
    0.001540046, 0.001535993, 0.001560099, 0.001549441, 0.001578987, 
    0.001570739, 0.001514928, 0.001517555, 0.001526694, 0.001522347, 
    0.001534775, 0.001537832, 0.001540316, 0.00154349, 0.001543833, 
    0.001545714, 0.001542632, 0.001545592, 0.00153439, 0.001539398, 
    0.00152565, 0.001528998, 0.001527458, 0.001525769, 0.001530982, 
    0.001536532, 0.001536652, 0.001538431, 0.00154344, 0.001534826, 
    0.001561472, 0.001545024, 0.00152042, 0.001525476, 0.001526199, 
    0.001524241, 0.001537525, 0.001532714, 0.001545668, 0.001542169, 
    0.001547901, 0.001545053, 0.001544634, 0.001540974, 0.001538695, 
    0.001532934, 0.001528245, 0.001524525, 0.00152539, 0.001529476, 
    0.001536872, 0.001543864, 0.001542333, 0.001547466, 0.001533875, 
    0.001539576, 0.001537372, 0.001543116, 0.001530526, 0.001541246, 
    0.001527784, 0.001528965, 0.001532618, 0.001539962, 0.001541587, 
    0.00154332, 0.001542251, 0.00153706, 0.001536209, 0.00153253, 
    0.001531513, 0.001528708, 0.001526385, 0.001528508, 0.001530736, 
    0.001537062, 0.00154276, 0.001548968, 0.001550487, 0.001557732, 
    0.001551833, 0.001561564, 0.00155329, 0.001567608, 0.001541868, 
    0.001553048, 0.001532785, 0.00153497, 0.001538921, 0.001547977, 
    0.001543089, 0.001548805, 0.001536176, 0.001529616, 0.001527919, 
    0.001524751, 0.001527992, 0.001527728, 0.001530829, 0.001529832, 
    0.001537272, 0.001533277, 0.001544623, 0.00154876, 0.001560434, 
    0.001567583, 0.001574856, 0.001578064, 0.00157904, 0.001579448,
  0.001428956, 0.001435721, 0.001434406, 0.001439862, 0.001436835, 
    0.001440408, 0.001430328, 0.00143599, 0.001432375, 0.001429565, 
    0.001450447, 0.001440105, 0.001461186, 0.001454593, 0.001471153, 
    0.00146016, 0.001473369, 0.001470836, 0.00147846, 0.001476276, 
    0.001486025, 0.001479468, 0.001491078, 0.00148446, 0.001485495, 
    0.001479252, 0.001442187, 0.001449159, 0.001441773, 0.001442768, 
    0.001442322, 0.001436898, 0.001434164, 0.001428439, 0.001429478, 
    0.001433684, 0.001443215, 0.00143998, 0.001448133, 0.001447949, 
    0.001457023, 0.001452932, 0.00146818, 0.001463847, 0.001476367, 
    0.001473219, 0.00147622, 0.00147531, 0.001476231, 0.001471614, 
    0.001473592, 0.001469529, 0.001453698, 0.001458352, 0.001444471, 
    0.001436122, 0.001430576, 0.00142664, 0.001427196, 0.001428257, 
    0.001433708, 0.001438833, 0.001442737, 0.001445349, 0.001447922, 
    0.00145571, 0.001459831, 0.001469056, 0.001467392, 0.001470212, 
    0.001472906, 0.001477428, 0.001476684, 0.001478676, 0.001470138, 
    0.001475813, 0.001466444, 0.001469006, 0.001448621, 0.001440853, 
    0.00143755, 0.001434659, 0.001427624, 0.001432482, 0.001430567, 
    0.001435123, 0.001438018, 0.001436586, 0.001445421, 0.001441986, 
    0.001460075, 0.001452285, 0.001472592, 0.001467734, 0.001473756, 
    0.001470683, 0.001475948, 0.00147121, 0.001479418, 0.001481205, 
    0.001479984, 0.001484674, 0.001470947, 0.00147622, 0.001436546, 
    0.001436779, 0.001437867, 0.001433085, 0.001432793, 0.00142841, 
    0.00143231, 0.001433971, 0.001438185, 0.001440678, 0.001443048, 
    0.001448257, 0.001454074, 0.001462207, 0.001468049, 0.001471964, 
    0.001469563, 0.001471682, 0.001469313, 0.001468203, 0.001480535, 
    0.001473611, 0.001484, 0.001483425, 0.001478724, 0.00148349, 0.001436943, 
    0.0014356, 0.001430934, 0.001434586, 0.001427933, 0.001431657, 
    0.001433798, 0.001442058, 0.001443872, 0.001445555, 0.001448878, 
    0.001453141, 0.00146062, 0.001467125, 0.001473063, 0.001472628, 
    0.001472781, 0.001474107, 0.001470822, 0.001474646, 0.001475288, 
    0.00147361, 0.001483348, 0.001480566, 0.001483413, 0.001481602, 
    0.001436037, 0.001438297, 0.001437076, 0.001439373, 0.001437754, 
    0.00144495, 0.001447107, 0.001457199, 0.001453057, 0.001459648, 
    0.001453727, 0.001454776, 0.001459863, 0.001454047, 0.001466766, 
    0.001458143, 0.001474159, 0.001465549, 0.001474698, 0.001473037, 
    0.001475787, 0.00147825, 0.001481348, 0.001487064, 0.00148574, 
    0.00149052, 0.001441667, 0.001444599, 0.001444341, 0.001447409, 
    0.001449678, 0.001454595, 0.001462479, 0.001459515, 0.001464957, 
    0.00146605, 0.001457781, 0.001462858, 0.001446561, 0.001449195, 
    0.001447627, 0.001441899, 0.001460198, 0.001450808, 0.001468145, 
    0.00146306, 0.001477899, 0.00147052, 0.001485012, 0.001491205, 
    0.001497032, 0.001503841, 0.001446199, 0.001444207, 0.001447774, 
    0.001452708, 0.001457285, 0.00146337, 0.001463992, 0.001465132, 
    0.001468084, 0.001470566, 0.001465492, 0.001471188, 0.001449805, 
    0.001461013, 0.001443454, 0.001448742, 0.001452417, 0.001450805, 
    0.001459176, 0.001461148, 0.001469163, 0.00146502, 0.001489676, 
    0.00147877, 0.001509024, 0.001500573, 0.001443511, 0.001446192, 
    0.001455522, 0.001451083, 0.001463776, 0.0014669, 0.001469439, 
    0.001472684, 0.001473034, 0.001474957, 0.001471806, 0.001474833, 
    0.001463383, 0.0014685, 0.001454456, 0.001457875, 0.001456302, 
    0.001454577, 0.001459901, 0.001465572, 0.001465694, 0.001467512, 
    0.001472635, 0.001463828, 0.001491083, 0.001474253, 0.001449116, 
    0.001454279, 0.001455017, 0.001453017, 0.001466586, 0.00146167, 
    0.00147491, 0.001471332, 0.001477194, 0.001474282, 0.001473853, 
    0.001470112, 0.001467782, 0.001461896, 0.001457106, 0.001453307, 
    0.00145419, 0.001458363, 0.001465919, 0.001473066, 0.001471501, 
    0.001476749, 0.001462856, 0.001468682, 0.00146643, 0.001472301, 
    0.001459436, 0.001470392, 0.001456635, 0.001457841, 0.001461573, 
    0.001469077, 0.001470737, 0.00147251, 0.001471416, 0.001466111, 
    0.001465242, 0.001461482, 0.001460444, 0.001457579, 0.001455206, 
    0.001457374, 0.00145965, 0.001466113, 0.001471937, 0.001478285, 
    0.001479838, 0.001487253, 0.001481217, 0.001491177, 0.001482709, 
    0.001497366, 0.001471027, 0.00148246, 0.001461742, 0.001463975, 
    0.001468013, 0.001477272, 0.001472274, 0.001478119, 0.001465208, 
    0.001458507, 0.001456773, 0.001453538, 0.001456847, 0.001456578, 
    0.001459744, 0.001458727, 0.001466328, 0.001462245, 0.001473842, 
    0.001478073, 0.001490019, 0.001497339, 0.00150479, 0.001508078, 
    0.001509079, 0.001509498,
  0.00134304, 0.00134928, 0.001348067, 0.001353102, 0.001350308, 0.001353606, 
    0.001344305, 0.001349528, 0.001346193, 0.001343602, 0.001362882, 
    0.001353327, 0.001372815, 0.001366714, 0.001382048, 0.001371866, 
    0.001384102, 0.001381754, 0.001388824, 0.001386798, 0.001395847, 
    0.001389759, 0.001400541, 0.001394393, 0.001395354, 0.001389558, 
    0.001355248, 0.001361692, 0.001354867, 0.001355785, 0.001355373, 
    0.001350366, 0.001347844, 0.001342563, 0.001343522, 0.0013474, 
    0.001356198, 0.001353211, 0.001360741, 0.001360571, 0.001368962, 
    0.001365178, 0.001379293, 0.001375279, 0.001386882, 0.001383963, 
    0.001386745, 0.001385901, 0.001386756, 0.001382475, 0.001384309, 
    0.001380542, 0.001365887, 0.001370192, 0.001357358, 0.001349651, 
    0.001344534, 0.001340905, 0.001341418, 0.001342396, 0.001347423, 
    0.001352152, 0.001355757, 0.001358169, 0.001360547, 0.001367748, 
    0.001371561, 0.001380105, 0.001378562, 0.001381175, 0.001383672, 
    0.001387866, 0.001387176, 0.001389024, 0.001381106, 0.001386368, 
    0.001377683, 0.001380058, 0.001361194, 0.001354016, 0.001350968, 
    0.0013483, 0.001341812, 0.001346292, 0.001344526, 0.001348728, 
    0.001351399, 0.001350078, 0.001358235, 0.001355063, 0.001371787, 
    0.00136458, 0.001383381, 0.001378878, 0.00138446, 0.001381612, 
    0.001386494, 0.0013821, 0.001389712, 0.001391371, 0.001390237, 
    0.001394592, 0.001381856, 0.001386745, 0.001350041, 0.001350257, 
    0.00135126, 0.001346849, 0.001346579, 0.001342537, 0.001346133, 
    0.001347665, 0.001351554, 0.001353855, 0.001356044, 0.001360857, 
    0.001366235, 0.00137376, 0.00137917, 0.001382799, 0.001380573, 
    0.001382538, 0.001380342, 0.001379313, 0.001390749, 0.001384326, 
    0.001393965, 0.001393432, 0.001389068, 0.001393492, 0.001350408, 
    0.001349168, 0.001344864, 0.001348232, 0.001342097, 0.001345531, 
    0.001347506, 0.00135513, 0.001356805, 0.00135836, 0.00136143, 
    0.001365372, 0.001372291, 0.001378315, 0.001383818, 0.001383414, 
    0.001383556, 0.001384786, 0.00138174, 0.001385286, 0.001385882, 
    0.001384325, 0.00139336, 0.001390778, 0.00139342, 0.001391739, 
    0.001349571, 0.001351657, 0.00135053, 0.00135265, 0.001351157, 
    0.001357801, 0.001359794, 0.001369125, 0.001365294, 0.001371391, 
    0.001365913, 0.001366884, 0.001371591, 0.001366209, 0.001377983, 
    0.001369999, 0.001384834, 0.001376856, 0.001385334, 0.001383794, 
    0.001386344, 0.001388629, 0.001391504, 0.001396811, 0.001395582, 
    0.001400022, 0.001354769, 0.001357477, 0.001357238, 0.001360073, 
    0.00136217, 0.001366716, 0.001374012, 0.001371268, 0.001376307, 
    0.001377319, 0.001369663, 0.001374363, 0.001359289, 0.001361723, 
    0.001360274, 0.001354982, 0.0013719, 0.001363214, 0.00137926, 
    0.001374549, 0.001388303, 0.001381461, 0.001394905, 0.001400659, 
    0.001406077, 0.001412414, 0.001358955, 0.001357114, 0.00136041, 
    0.001364971, 0.001369205, 0.001374837, 0.001375413, 0.001376469, 
    0.001379203, 0.001381503, 0.001376803, 0.00138208, 0.001362288, 
    0.001372655, 0.001356419, 0.001361305, 0.001364702, 0.001363212, 
    0.001370954, 0.00137278, 0.001380203, 0.001376365, 0.001399239, 
    0.001389112, 0.001417242, 0.001409372, 0.001356472, 0.001358948, 
    0.001367574, 0.001363469, 0.001375213, 0.001378106, 0.001380458, 
    0.001383467, 0.001383791, 0.001385574, 0.001382653, 0.001385459, 
    0.001374849, 0.001379589, 0.001366587, 0.00136975, 0.001368295, 
    0.001366699, 0.001371625, 0.001376877, 0.001376989, 0.001378673, 
    0.001383423, 0.00137526, 0.001400548, 0.001384923, 0.00136165, 
    0.001366424, 0.001367106, 0.001365256, 0.001377816, 0.001373263, 
    0.001385531, 0.001382213, 0.001387649, 0.001384948, 0.00138455, 
    0.001381082, 0.001378923, 0.001373472, 0.001369039, 0.001365524, 
    0.001366341, 0.001370202, 0.001377198, 0.001383821, 0.00138237, 
    0.001387236, 0.001374361, 0.001379758, 0.001377671, 0.001383112, 
    0.001371195, 0.001381343, 0.001368603, 0.001369719, 0.001373173, 
    0.001380124, 0.001381662, 0.001383305, 0.001382291, 0.001377376, 
    0.00137657, 0.001373089, 0.001372128, 0.001369476, 0.001367281, 
    0.001369287, 0.001371393, 0.001377377, 0.001382774, 0.001388661, 
    0.001390102, 0.001396988, 0.001391383, 0.001400635, 0.001392769, 
    0.001406389, 0.001381931, 0.001392537, 0.00137333, 0.001375397, 
    0.001379138, 0.001387722, 0.001383086, 0.001388508, 0.001376539, 
    0.001370335, 0.001368731, 0.001365738, 0.001368799, 0.00136855, 
    0.00137148, 0.001370538, 0.001377576, 0.001373795, 0.00138454, 
    0.001388465, 0.001399557, 0.001406363, 0.001413297, 0.00141636, 
    0.001417292, 0.001417682,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3 =
  1.21246e-06, 1.222928e-06, 1.220889e-06, 1.229358e-06, 1.224656e-06, 
    1.230207e-06, 1.214578e-06, 1.223343e-06, 1.217744e-06, 1.213399e-06, 
    1.24588e-06, 1.229736e-06, 1.262769e-06, 1.252386e-06, 1.278553e-06, 
    1.26115e-06, 1.282077e-06, 1.278049e-06, 1.290193e-06, 1.286707e-06, 
    1.302304e-06, 1.291802e-06, 1.310428e-06, 1.299792e-06, 1.301452e-06, 
    1.291456e-06, 1.232978e-06, 1.243865e-06, 1.232334e-06, 1.233883e-06, 
    1.233188e-06, 1.224753e-06, 1.220513e-06, 1.211661e-06, 1.213265e-06, 
    1.219768e-06, 1.234579e-06, 1.229541e-06, 1.242258e-06, 1.241971e-06, 
    1.256207e-06, 1.249778e-06, 1.273834e-06, 1.266972e-06, 1.286853e-06, 
    1.281837e-06, 1.286616e-06, 1.285166e-06, 1.286635e-06, 1.279284e-06, 
    1.28243e-06, 1.275972e-06, 1.250982e-06, 1.2583e-06, 1.236539e-06, 
    1.223548e-06, 1.214961e-06, 1.208886e-06, 1.209744e-06, 1.21138e-06, 
    1.219806e-06, 1.227757e-06, 1.233834e-06, 1.237908e-06, 1.241929e-06, 
    1.25414e-06, 1.260629e-06, 1.275223e-06, 1.272583e-06, 1.277057e-06, 
    1.281339e-06, 1.288544e-06, 1.287357e-06, 1.290536e-06, 1.276938e-06, 
    1.285967e-06, 1.271079e-06, 1.275142e-06, 1.243023e-06, 1.2309e-06, 
    1.225764e-06, 1.221279e-06, 1.210403e-06, 1.217908e-06, 1.214947e-06, 
    1.221999e-06, 1.22649e-06, 1.224268e-06, 1.238019e-06, 1.232663e-06, 
    1.261014e-06, 1.248761e-06, 1.280839e-06, 1.273124e-06, 1.282692e-06, 
    1.277805e-06, 1.286183e-06, 1.278641e-06, 1.291721e-06, 1.294578e-06, 
    1.292625e-06, 1.300135e-06, 1.278223e-06, 1.286615e-06, 1.224206e-06, 
    1.224568e-06, 1.226257e-06, 1.218842e-06, 1.218389e-06, 1.211616e-06, 
    1.217641e-06, 1.220212e-06, 1.226751e-06, 1.230627e-06, 1.234317e-06, 
    1.242452e-06, 1.25157e-06, 1.264379e-06, 1.273623e-06, 1.27984e-06, 
    1.276026e-06, 1.279392e-06, 1.275629e-06, 1.273867e-06, 1.293506e-06, 
    1.282459e-06, 1.299053e-06, 1.298132e-06, 1.290611e-06, 1.298236e-06, 
    1.224823e-06, 1.222738e-06, 1.215514e-06, 1.221165e-06, 1.210879e-06, 
    1.216631e-06, 1.219944e-06, 1.232774e-06, 1.235603e-06, 1.238228e-06, 
    1.243423e-06, 1.250105e-06, 1.261873e-06, 1.272159e-06, 1.281588e-06, 
    1.280895e-06, 1.281139e-06, 1.283249e-06, 1.278024e-06, 1.284108e-06, 
    1.28513e-06, 1.282458e-06, 1.298008e-06, 1.293556e-06, 1.298112e-06, 
    1.295212e-06, 1.223415e-06, 1.226925e-06, 1.225027e-06, 1.228596e-06, 
    1.226081e-06, 1.237284e-06, 1.240653e-06, 1.256482e-06, 1.249973e-06, 
    1.260341e-06, 1.251024e-06, 1.252672e-06, 1.260678e-06, 1.251526e-06, 
    1.27159e-06, 1.257969e-06, 1.283331e-06, 1.269662e-06, 1.28419e-06, 
    1.281546e-06, 1.285925e-06, 1.289854e-06, 1.294806e-06, 1.303969e-06, 
    1.301844e-06, 1.309526e-06, 1.232167e-06, 1.236737e-06, 1.236334e-06, 
    1.241126e-06, 1.244675e-06, 1.252388e-06, 1.264809e-06, 1.26013e-06, 
    1.268726e-06, 1.270456e-06, 1.257399e-06, 1.265407e-06, 1.239799e-06, 
    1.243917e-06, 1.241464e-06, 1.232525e-06, 1.261206e-06, 1.246443e-06, 
    1.273775e-06, 1.265724e-06, 1.289293e-06, 1.277543e-06, 1.300675e-06, 
    1.310628e-06, 1.320034e-06, 1.331069e-06, 1.239235e-06, 1.236125e-06, 
    1.241696e-06, 1.249425e-06, 1.256619e-06, 1.266216e-06, 1.2672e-06, 
    1.269003e-06, 1.273679e-06, 1.277618e-06, 1.269573e-06, 1.278606e-06, 
    1.244873e-06, 1.262492e-06, 1.234948e-06, 1.243208e-06, 1.248966e-06, 
    1.246439e-06, 1.259595e-06, 1.262705e-06, 1.275388e-06, 1.268824e-06, 
    1.308167e-06, 1.290683e-06, 1.339503e-06, 1.325765e-06, 1.235039e-06, 
    1.239224e-06, 1.253845e-06, 1.246877e-06, 1.266858e-06, 1.271802e-06, 
    1.275828e-06, 1.280984e-06, 1.281542e-06, 1.284603e-06, 1.279588e-06, 
    1.284404e-06, 1.266235e-06, 1.274338e-06, 1.252168e-06, 1.257544e-06, 
    1.255069e-06, 1.252357e-06, 1.260737e-06, 1.269697e-06, 1.269889e-06, 
    1.27277e-06, 1.280903e-06, 1.266937e-06, 1.310431e-06, 1.283478e-06, 
    1.243795e-06, 1.251891e-06, 1.25305e-06, 1.249909e-06, 1.271305e-06, 
    1.26353e-06, 1.284528e-06, 1.278835e-06, 1.288169e-06, 1.283526e-06, 
    1.282844e-06, 1.276895e-06, 1.273199e-06, 1.263885e-06, 1.256333e-06, 
    1.250363e-06, 1.251749e-06, 1.258313e-06, 1.270246e-06, 1.28159e-06, 
    1.2791e-06, 1.287457e-06, 1.265401e-06, 1.274625e-06, 1.271055e-06, 
    1.280373e-06, 1.260006e-06, 1.27734e-06, 1.255594e-06, 1.257493e-06, 
    1.263376e-06, 1.275253e-06, 1.27789e-06, 1.280707e-06, 1.278968e-06, 
    1.270551e-06, 1.269175e-06, 1.263232e-06, 1.261593e-06, 1.257078e-06, 
    1.253346e-06, 1.256755e-06, 1.260341e-06, 1.270554e-06, 1.279794e-06, 
    1.289908e-06, 1.29239e-06, 1.304271e-06, 1.294594e-06, 1.310581e-06, 
    1.296981e-06, 1.320571e-06, 1.278349e-06, 1.296586e-06, 1.263644e-06, 
    1.267172e-06, 1.273565e-06, 1.288293e-06, 1.280331e-06, 1.289645e-06, 
    1.269121e-06, 1.25854e-06, 1.25581e-06, 1.250725e-06, 1.255926e-06, 
    1.255503e-06, 1.26049e-06, 1.258886e-06, 1.270893e-06, 1.264436e-06, 
    1.282825e-06, 1.28957e-06, 1.308718e-06, 1.320529e-06, 1.332609e-06, 
    1.33796e-06, 1.339592e-06, 1.340273e-06 ;

 SMIN_NO3_LEACHED =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_RUNOFF =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SMIN_NO3_vr =
  7.531931e-06, 7.565989e-06, 7.559351e-06, 7.586841e-06, 7.571584e-06, 
    7.589571e-06, 7.538798e-06, 7.567281e-06, 7.549087e-06, 7.534936e-06, 
    7.640187e-06, 7.588005e-06, 7.694573e-06, 7.661181e-06, 7.745125e-06, 
    7.689343e-06, 7.756383e-06, 7.743511e-06, 7.782272e-06, 7.771149e-06, 
    7.820747e-06, 7.78738e-06, 7.846511e-06, 7.81277e-06, 7.818027e-06, 
    7.786238e-06, 7.598571e-06, 7.633738e-06, 7.596469e-06, 7.601483e-06, 
    7.599227e-06, 7.571859e-06, 7.558071e-06, 7.529267e-06, 7.534484e-06, 
    7.55564e-06, 7.603679e-06, 7.587356e-06, 7.628506e-06, 7.627578e-06, 
    7.673451e-06, 7.652751e-06, 7.730014e-06, 7.708019e-06, 7.771604e-06, 
    7.755582e-06, 7.770833e-06, 7.766196e-06, 7.770869e-06, 7.747397e-06, 
    7.757433e-06, 7.736794e-06, 7.656719e-06, 7.680261e-06, 7.610067e-06, 
    7.567921e-06, 7.54001e-06, 7.52022e-06, 7.522999e-06, 7.528331e-06, 
    7.555747e-06, 7.581566e-06, 7.601261e-06, 7.614432e-06, 7.62742e-06, 
    7.666767e-06, 7.687643e-06, 7.734434e-06, 7.725993e-06, 7.740287e-06, 
    7.753982e-06, 7.776962e-06, 7.773175e-06, 7.783293e-06, 7.739877e-06, 
    7.768713e-06, 7.721112e-06, 7.734117e-06, 7.630979e-06, 7.591794e-06, 
    7.57511e-06, 7.560551e-06, 7.525143e-06, 7.549581e-06, 7.539933e-06, 
    7.562866e-06, 7.577447e-06, 7.570223e-06, 7.614783e-06, 7.597433e-06, 
    7.688869e-06, 7.649441e-06, 7.752394e-06, 7.727707e-06, 7.75829e-06, 
    7.742679e-06, 7.769414e-06, 7.745338e-06, 7.787053e-06, 7.796144e-06, 
    7.789913e-06, 7.813809e-06, 7.743951e-06, 7.770745e-06, 7.570065e-06, 
    7.571243e-06, 7.576717e-06, 7.552604e-06, 7.55113e-06, 7.529072e-06, 
    7.548681e-06, 7.557039e-06, 7.578275e-06, 7.590828e-06, 7.602773e-06, 
    7.629082e-06, 7.658475e-06, 7.699655e-06, 7.729296e-06, 7.749171e-06, 
    7.736975e-06, 7.747726e-06, 7.735688e-06, 7.730039e-06, 7.79271e-06, 
    7.757491e-06, 7.810347e-06, 7.807423e-06, 7.783467e-06, 7.807728e-06, 
    7.572053e-06, 7.565274e-06, 7.541774e-06, 7.560148e-06, 7.526657e-06, 
    7.545386e-06, 7.556146e-06, 7.597771e-06, 7.606933e-06, 7.615424e-06, 
    7.632203e-06, 7.653747e-06, 7.691602e-06, 7.724585e-06, 7.754747e-06, 
    7.752525e-06, 7.753299e-06, 7.760023e-06, 7.743326e-06, 7.762749e-06, 
    7.765996e-06, 7.757472e-06, 7.807006e-06, 7.792843e-06, 7.807327e-06, 
    7.798092e-06, 7.567466e-06, 7.578844e-06, 7.572677e-06, 7.584254e-06, 
    7.576076e-06, 7.612367e-06, 7.623247e-06, 7.674276e-06, 7.65332e-06, 
    7.686681e-06, 7.656695e-06, 7.662001e-06, 7.687719e-06, 7.658296e-06, 
    7.722728e-06, 7.678989e-06, 7.760276e-06, 7.71651e-06, 7.763003e-06, 
    7.75455e-06, 7.768521e-06, 7.781044e-06, 7.796798e-06, 7.825909e-06, 
    7.81915e-06, 7.843523e-06, 7.595831e-06, 7.610606e-06, 7.609312e-06, 
    7.624791e-06, 7.636241e-06, 7.661116e-06, 7.701038e-06, 7.686005e-06, 
    7.713588e-06, 7.719129e-06, 7.677198e-06, 7.702915e-06, 7.620433e-06, 
    7.633715e-06, 7.625803e-06, 7.596866e-06, 7.689382e-06, 7.641838e-06, 
    7.729686e-06, 7.703874e-06, 7.779233e-06, 7.741713e-06, 7.815432e-06, 
    7.846988e-06, 7.876761e-06, 7.911533e-06, 7.618683e-06, 7.608618e-06, 
    7.626621e-06, 7.651547e-06, 7.674708e-06, 7.705543e-06, 7.708695e-06, 
    7.71446e-06, 7.729435e-06, 7.742038e-06, 7.716257e-06, 7.745176e-06, 
    7.636768e-06, 7.693515e-06, 7.604701e-06, 7.631395e-06, 7.649967e-06, 
    7.641824e-06, 7.684186e-06, 7.694167e-06, 7.734802e-06, 7.71379e-06, 
    7.839163e-06, 7.783614e-06, 7.938068e-06, 7.894807e-06, 7.605094e-06, 
    7.61862e-06, 7.665769e-06, 7.643323e-06, 7.707585e-06, 7.72343e-06, 
    7.736307e-06, 7.752786e-06, 7.754555e-06, 7.764326e-06, 7.7483e-06, 
    7.763681e-06, 7.70552e-06, 7.731491e-06, 7.660298e-06, 7.677585e-06, 
    7.669625e-06, 7.66088e-06, 7.68783e-06, 7.716568e-06, 7.71719e-06, 
    7.726395e-06, 7.752355e-06, 7.707696e-06, 7.846276e-06, 7.76056e-06, 
    7.633381e-06, 7.659458e-06, 7.663197e-06, 7.653084e-06, 7.721816e-06, 
    7.696884e-06, 7.76409e-06, 7.745897e-06, 7.775685e-06, 7.760874e-06, 
    7.758676e-06, 7.739671e-06, 7.727821e-06, 7.697959e-06, 7.673672e-06, 
    7.654457e-06, 7.658907e-06, 7.680024e-06, 7.718307e-06, 7.754607e-06, 
    7.746638e-06, 7.773317e-06, 7.702751e-06, 7.732305e-06, 7.720855e-06, 
    7.750679e-06, 7.685569e-06, 7.741096e-06, 7.67138e-06, 7.677475e-06, 
    7.696365e-06, 7.734422e-06, 7.742858e-06, 7.751857e-06, 7.74629e-06, 
    7.719344e-06, 7.714929e-06, 7.695856e-06, 7.690576e-06, 7.676073e-06, 
    7.664044e-06, 7.675016e-06, 7.686519e-06, 7.719298e-06, 7.748853e-06, 
    7.781118e-06, 7.789027e-06, 7.826745e-06, 7.795998e-06, 7.84671e-06, 
    7.803537e-06, 7.878315e-06, 7.74432e-06, 7.802473e-06, 7.697233e-06, 
    7.708541e-06, 7.729006e-06, 7.776041e-06, 7.750639e-06, 7.780346e-06, 
    7.714752e-06, 7.680758e-06, 7.671984e-06, 7.65561e-06, 7.672344e-06, 
    7.670983e-06, 7.68701e-06, 7.681843e-06, 7.720364e-06, 7.699662e-06, 
    7.758508e-06, 7.780019e-06, 7.840868e-06, 7.878219e-06, 7.916331e-06, 
    7.933151e-06, 7.938275e-06, 7.940408e-06,
  3.965845e-06, 3.995977e-06, 3.990114e-06, 4.014464e-06, 4.000952e-06, 
    4.016904e-06, 3.97195e-06, 3.997172e-06, 3.981066e-06, 3.968558e-06, 
    4.061866e-06, 4.015552e-06, 4.110216e-06, 4.080519e-06, 4.15528e-06, 
    4.105585e-06, 4.165328e-06, 4.153851e-06, 4.188449e-06, 4.178527e-06, 
    4.222878e-06, 4.193031e-06, 4.245948e-06, 4.215747e-06, 4.220464e-06, 
    4.192047e-06, 4.024863e-06, 4.056087e-06, 4.023015e-06, 4.027461e-06, 
    4.025467e-06, 4.001229e-06, 3.98903e-06, 3.96355e-06, 3.968173e-06, 
    3.986892e-06, 4.029461e-06, 4.014997e-06, 4.051503e-06, 4.050677e-06, 
    4.091457e-06, 4.073052e-06, 4.141825e-06, 4.122237e-06, 4.178941e-06, 
    4.164653e-06, 4.178268e-06, 4.174139e-06, 4.178322e-06, 4.157374e-06, 
    4.166344e-06, 4.147931e-06, 4.076495e-06, 4.097439e-06, 4.035087e-06, 
    3.997758e-06, 3.973053e-06, 3.955553e-06, 3.958025e-06, 3.962738e-06, 
    3.987001e-06, 4.009871e-06, 4.02733e-06, 4.039024e-06, 4.050559e-06, 
    4.08553e-06, 4.104102e-06, 4.145787e-06, 4.138259e-06, 4.151019e-06, 
    4.163232e-06, 4.183758e-06, 4.180378e-06, 4.189429e-06, 4.150687e-06, 
    4.176418e-06, 4.133972e-06, 4.145564e-06, 4.053672e-06, 4.018898e-06, 
    4.00413e-06, 3.99124e-06, 3.959926e-06, 3.98154e-06, 3.973013e-06, 
    3.993314e-06, 4.00623e-06, 3.999841e-06, 4.039343e-06, 4.023968e-06, 
    4.105204e-06, 4.070138e-06, 4.161807e-06, 4.139804e-06, 4.167089e-06, 
    4.153159e-06, 4.177035e-06, 4.155545e-06, 4.192801e-06, 4.200927e-06, 
    4.195373e-06, 4.216731e-06, 4.154354e-06, 4.178265e-06, 3.999661e-06, 
    4.000703e-06, 4.00556e-06, 3.984227e-06, 3.982924e-06, 3.963422e-06, 
    3.980776e-06, 3.988172e-06, 4.006982e-06, 4.018118e-06, 4.028718e-06, 
    4.052059e-06, 4.078183e-06, 4.114825e-06, 4.141229e-06, 4.158961e-06, 
    4.148086e-06, 4.157686e-06, 4.146954e-06, 4.141928e-06, 4.19788e-06, 
    4.166426e-06, 4.213657e-06, 4.211039e-06, 4.189643e-06, 4.211334e-06, 
    4.001435e-06, 3.995441e-06, 3.97465e-06, 3.990917e-06, 3.961301e-06, 
    3.977865e-06, 3.9874e-06, 4.024283e-06, 4.03241e-06, 4.039944e-06, 
    4.054843e-06, 4.073992e-06, 4.107664e-06, 4.137049e-06, 4.163945e-06, 
    4.161972e-06, 4.162666e-06, 4.16868e-06, 4.153786e-06, 4.171127e-06, 
    4.174038e-06, 4.166426e-06, 4.210688e-06, 4.198026e-06, 4.210983e-06, 
    4.202738e-06, 3.99739e-06, 4.00748e-06, 4.002026e-06, 4.012282e-06, 
    4.005054e-06, 4.037228e-06, 4.046893e-06, 4.092241e-06, 4.073614e-06, 
    4.103282e-06, 4.076626e-06, 4.081343e-06, 4.10424e-06, 4.078066e-06, 
    4.135421e-06, 4.096495e-06, 4.168914e-06, 4.129914e-06, 4.171362e-06, 
    4.163828e-06, 4.176306e-06, 4.187491e-06, 4.201583e-06, 4.227621e-06, 
    4.221587e-06, 4.2434e-06, 4.022542e-06, 4.03566e-06, 4.034509e-06, 
    4.048256e-06, 4.058433e-06, 4.08053e-06, 4.116057e-06, 4.102686e-06, 
    4.127252e-06, 4.132188e-06, 4.094874e-06, 4.117765e-06, 4.044452e-06, 
    4.056258e-06, 4.049231e-06, 4.023574e-06, 4.105759e-06, 4.0635e-06, 
    4.141665e-06, 4.118679e-06, 4.185895e-06, 4.152412e-06, 4.218266e-06, 
    4.246519e-06, 4.273196e-06, 4.30442e-06, 4.042831e-06, 4.03391e-06, 
    4.049894e-06, 4.072038e-06, 4.092639e-06, 4.120078e-06, 4.122892e-06, 
    4.12804e-06, 4.141392e-06, 4.152628e-06, 4.129664e-06, 4.155447e-06, 
    4.058989e-06, 4.109437e-06, 4.030534e-06, 4.054227e-06, 4.070734e-06, 
    4.063495e-06, 4.101159e-06, 4.110054e-06, 4.146269e-06, 4.127536e-06, 
    4.239535e-06, 4.189848e-06, 4.328265e-06, 4.289418e-06, 4.030793e-06, 
    4.042803e-06, 4.084698e-06, 4.064745e-06, 4.121915e-06, 4.136031e-06, 
    4.147523e-06, 4.162223e-06, 4.163815e-06, 4.172535e-06, 4.158248e-06, 
    4.171972e-06, 4.120137e-06, 4.143272e-06, 4.079906e-06, 4.095293e-06, 
    4.088214e-06, 4.08045e-06, 4.104428e-06, 4.130024e-06, 4.130579e-06, 
    4.138798e-06, 4.161976e-06, 4.122148e-06, 4.245949e-06, 4.169321e-06, 
    4.055913e-06, 4.079101e-06, 4.082426e-06, 4.073434e-06, 4.134615e-06, 
    4.112407e-06, 4.172324e-06, 4.156101e-06, 4.182696e-06, 4.169472e-06, 
    4.167527e-06, 4.15057e-06, 4.140023e-06, 4.113422e-06, 4.091828e-06, 
    4.074739e-06, 4.07871e-06, 4.097491e-06, 4.131593e-06, 4.163956e-06, 
    4.156857e-06, 4.180673e-06, 4.11776e-06, 4.144094e-06, 4.133905e-06, 
    4.160491e-06, 4.102329e-06, 4.151815e-06, 4.089712e-06, 4.095145e-06, 
    4.111966e-06, 4.145877e-06, 4.153404e-06, 4.161434e-06, 4.15648e-06, 
    4.132462e-06, 4.128535e-06, 4.111559e-06, 4.106872e-06, 4.093963e-06, 
    4.083282e-06, 4.093038e-06, 4.103291e-06, 4.132475e-06, 4.158836e-06, 
    4.187649e-06, 4.194715e-06, 4.228473e-06, 4.200974e-06, 4.246376e-06, 
    4.207748e-06, 4.274704e-06, 4.1547e-06, 4.20663e-06, 4.112735e-06, 
    4.122815e-06, 4.141061e-06, 4.18304e-06, 4.160366e-06, 4.186891e-06, 
    4.128382e-06, 4.098136e-06, 4.090334e-06, 4.075775e-06, 4.090667e-06, 
    4.089455e-06, 4.103721e-06, 4.099135e-06, 4.133446e-06, 4.115003e-06, 
    4.167476e-06, 4.186683e-06, 4.241109e-06, 4.274594e-06, 4.30879e-06, 
    4.323913e-06, 4.328521e-06, 4.330447e-06,
  3.780339e-06, 3.813908e-06, 3.807373e-06, 3.834519e-06, 3.819452e-06, 
    3.83724e-06, 3.787136e-06, 3.815241e-06, 3.79729e-06, 3.783358e-06, 
    3.88743e-06, 3.835733e-06, 3.941459e-06, 3.908257e-06, 3.991896e-06, 
    3.936283e-06, 4.00315e-06, 3.990291e-06, 4.029057e-06, 4.017935e-06, 
    4.067682e-06, 4.034194e-06, 4.093577e-06, 4.059676e-06, 4.06497e-06, 
    4.033091e-06, 3.846116e-06, 3.880976e-06, 3.844054e-06, 3.849016e-06, 
    3.84679e-06, 3.819761e-06, 3.806169e-06, 3.777782e-06, 3.782929e-06, 
    3.803784e-06, 3.851248e-06, 3.83511e-06, 3.875845e-06, 3.874923e-06, 
    3.920481e-06, 3.899912e-06, 3.976826e-06, 3.954902e-06, 4.0184e-06, 
    4.00239e-06, 4.017646e-06, 4.013018e-06, 4.017706e-06, 3.994237e-06, 
    4.004286e-06, 3.983661e-06, 3.90376e-06, 3.927169e-06, 3.857524e-06, 
    3.815898e-06, 3.788366e-06, 3.768879e-06, 3.771631e-06, 3.77688e-06, 
    3.803906e-06, 3.829394e-06, 3.848867e-06, 3.861915e-06, 3.874791e-06, 
    3.913865e-06, 3.934623e-06, 3.981263e-06, 3.972832e-06, 3.987122e-06, 
    4.000799e-06, 4.0238e-06, 4.020011e-06, 4.030157e-06, 3.986747e-06, 
    4.015574e-06, 3.968033e-06, 3.981012e-06, 3.87828e-06, 3.839462e-06, 
    3.823001e-06, 3.808628e-06, 3.773748e-06, 3.79782e-06, 3.788322e-06, 
    3.810937e-06, 3.825336e-06, 3.818212e-06, 3.862272e-06, 3.845116e-06, 
    3.935854e-06, 3.89666e-06, 3.999202e-06, 3.974563e-06, 4.005118e-06, 
    3.989515e-06, 4.016265e-06, 3.992187e-06, 4.033937e-06, 4.043051e-06, 
    4.036822e-06, 4.060777e-06, 3.990854e-06, 4.017645e-06, 3.818012e-06, 
    3.819173e-06, 3.824587e-06, 3.800814e-06, 3.799362e-06, 3.77764e-06, 
    3.796967e-06, 3.805209e-06, 3.826172e-06, 3.838592e-06, 3.850416e-06, 
    3.876467e-06, 3.905648e-06, 3.946613e-06, 3.976158e-06, 3.996013e-06, 
    3.983834e-06, 3.994586e-06, 3.982567e-06, 3.97694e-06, 4.039634e-06, 
    4.004378e-06, 4.057328e-06, 4.054391e-06, 4.030398e-06, 4.054722e-06, 
    3.819989e-06, 3.813307e-06, 3.790144e-06, 3.808266e-06, 3.775277e-06, 
    3.793726e-06, 3.80435e-06, 3.845471e-06, 3.854535e-06, 3.862943e-06, 
    3.879575e-06, 3.900963e-06, 3.938603e-06, 3.97148e-06, 4.001596e-06, 
    3.999386e-06, 4.000164e-06, 4.006902e-06, 3.990218e-06, 4.009644e-06, 
    4.012907e-06, 4.004376e-06, 4.053998e-06, 4.039795e-06, 4.054329e-06, 
    4.045079e-06, 3.815479e-06, 3.826728e-06, 3.820648e-06, 3.832085e-06, 
    3.824025e-06, 3.859916e-06, 3.870704e-06, 3.921361e-06, 3.900541e-06, 
    3.933703e-06, 3.903906e-06, 3.909177e-06, 3.934781e-06, 3.905514e-06, 
    3.969662e-06, 3.926118e-06, 4.007164e-06, 3.963502e-06, 4.009906e-06, 
    4.001465e-06, 4.015447e-06, 4.027985e-06, 4.043784e-06, 4.073e-06, 
    4.066228e-06, 4.090713e-06, 3.843526e-06, 3.858164e-06, 3.856876e-06, 
    3.872221e-06, 3.883584e-06, 3.908267e-06, 3.94799e-06, 3.933033e-06, 
    3.960513e-06, 3.966038e-06, 3.924299e-06, 3.949901e-06, 3.867976e-06, 
    3.88116e-06, 3.87331e-06, 3.844678e-06, 3.936474e-06, 3.889247e-06, 
    3.976646e-06, 3.950922e-06, 4.026196e-06, 3.988683e-06, 4.062501e-06, 
    4.094223e-06, 4.124186e-06, 4.1593e-06, 3.866166e-06, 3.856208e-06, 
    3.874048e-06, 3.898784e-06, 3.921802e-06, 3.952488e-06, 3.955635e-06, 
    3.961396e-06, 3.976339e-06, 3.988921e-06, 3.963216e-06, 3.992077e-06, 
    3.884215e-06, 3.940586e-06, 3.852444e-06, 3.878892e-06, 3.897325e-06, 
    3.889237e-06, 3.931326e-06, 3.941273e-06, 3.981802e-06, 3.960831e-06, 
    4.086382e-06, 4.030631e-06, 4.186129e-06, 4.142426e-06, 3.852731e-06, 
    3.866132e-06, 3.912927e-06, 3.890633e-06, 3.954542e-06, 3.97034e-06, 
    3.983204e-06, 3.999669e-06, 4.001451e-06, 4.011222e-06, 3.995215e-06, 
    4.010591e-06, 3.952554e-06, 3.978445e-06, 3.907569e-06, 3.924769e-06, 
    3.916854e-06, 3.908177e-06, 3.934982e-06, 3.96362e-06, 3.964237e-06, 
    3.973438e-06, 3.999408e-06, 3.954802e-06, 4.093592e-06, 4.007634e-06, 
    3.880769e-06, 3.906676e-06, 3.910387e-06, 3.900338e-06, 3.968754e-06, 
    3.943906e-06, 4.010984e-06, 3.99281e-06, 4.022608e-06, 4.007789e-06, 
    4.00561e-06, 3.986615e-06, 3.974808e-06, 3.945043e-06, 3.920896e-06, 
    3.901795e-06, 3.906233e-06, 3.927228e-06, 3.965376e-06, 4.00161e-06, 
    3.99366e-06, 4.02034e-06, 3.949893e-06, 3.979367e-06, 3.967963e-06, 
    3.997728e-06, 3.932635e-06, 3.988024e-06, 3.918528e-06, 3.924602e-06, 
    3.943414e-06, 3.981366e-06, 3.98979e-06, 3.998785e-06, 3.993235e-06, 
    3.966347e-06, 3.961951e-06, 3.942956e-06, 3.937717e-06, 3.92328e-06, 
    3.911342e-06, 3.922247e-06, 3.933713e-06, 3.96636e-06, 3.995876e-06, 
    4.028162e-06, 4.036082e-06, 4.073965e-06, 4.04311e-06, 4.094073e-06, 
    4.050719e-06, 4.125893e-06, 3.99125e-06, 4.049455e-06, 3.944272e-06, 
    3.955548e-06, 3.975974e-06, 4.023e-06, 3.997588e-06, 4.027316e-06, 
    3.961779e-06, 3.927951e-06, 3.919224e-06, 3.902955e-06, 3.919596e-06, 
    3.918241e-06, 3.934191e-06, 3.929063e-06, 3.967446e-06, 3.946809e-06, 
    4.005554e-06, 4.027082e-06, 4.088143e-06, 4.125762e-06, 4.16421e-06, 
    4.181228e-06, 4.186414e-06, 4.188583e-06,
  3.868284e-06, 3.905084e-06, 3.897917e-06, 3.927694e-06, 3.911163e-06, 
    3.93068e-06, 3.875731e-06, 3.906548e-06, 3.886862e-06, 3.87159e-06, 
    3.985792e-06, 3.929025e-06, 4.04518e-06, 4.008669e-06, 4.100689e-06, 
    4.039487e-06, 4.113084e-06, 4.098919e-06, 4.141627e-06, 4.12937e-06, 
    4.184225e-06, 4.147289e-06, 4.212799e-06, 4.175391e-06, 4.181232e-06, 
    4.146073e-06, 3.940419e-06, 3.978703e-06, 3.938156e-06, 3.943603e-06, 
    3.941158e-06, 3.911503e-06, 3.8966e-06, 3.865478e-06, 3.87112e-06, 
    3.893982e-06, 3.946053e-06, 3.92834e-06, 3.973056e-06, 3.972044e-06, 
    4.022106e-06, 3.999497e-06, 4.084093e-06, 4.059963e-06, 4.129881e-06, 
    4.112243e-06, 4.129052e-06, 4.123951e-06, 4.129118e-06, 4.103265e-06, 
    4.114332e-06, 4.091618e-06, 4.003726e-06, 4.029461e-06, 3.952942e-06, 
    3.907271e-06, 3.87708e-06, 3.855725e-06, 3.85874e-06, 3.864492e-06, 
    3.894116e-06, 3.922069e-06, 3.943436e-06, 3.95776e-06, 3.971898e-06, 
    4.014839e-06, 4.03766e-06, 4.08898e-06, 4.079696e-06, 4.095431e-06, 
    4.110491e-06, 4.135833e-06, 4.131657e-06, 4.142841e-06, 4.095016e-06, 
    4.12677e-06, 4.074413e-06, 4.088701e-06, 3.975743e-06, 3.933116e-06, 
    3.915061e-06, 3.899294e-06, 3.86106e-06, 3.887444e-06, 3.877032e-06, 
    3.901824e-06, 3.917617e-06, 3.909802e-06, 3.958152e-06, 3.939321e-06, 
    4.039014e-06, 3.995925e-06, 4.108732e-06, 4.081601e-06, 4.115248e-06, 
    4.098063e-06, 4.127531e-06, 4.101005e-06, 4.147007e-06, 4.157056e-06, 
    4.150188e-06, 4.176603e-06, 4.099537e-06, 4.129051e-06, 3.909583e-06, 
    3.910857e-06, 3.916795e-06, 3.890726e-06, 3.889134e-06, 3.865324e-06, 
    3.886507e-06, 3.895545e-06, 3.918533e-06, 3.932161e-06, 3.945138e-06, 
    3.973741e-06, 4.005803e-06, 4.050847e-06, 4.083357e-06, 4.105219e-06, 
    4.091808e-06, 4.103647e-06, 4.090413e-06, 4.084217e-06, 4.153289e-06, 
    4.114435e-06, 4.172799e-06, 4.169559e-06, 4.143107e-06, 4.169924e-06, 
    3.911752e-06, 3.904423e-06, 3.879028e-06, 3.898895e-06, 3.862735e-06, 
    3.882955e-06, 3.894605e-06, 3.939713e-06, 3.949659e-06, 3.95889e-06, 
    3.977154e-06, 4.000653e-06, 4.042035e-06, 4.078209e-06, 4.111368e-06, 
    4.108934e-06, 4.109791e-06, 4.117214e-06, 4.098838e-06, 4.120235e-06, 
    4.123831e-06, 4.114431e-06, 4.169125e-06, 4.153464e-06, 4.16949e-06, 
    4.159289e-06, 3.906805e-06, 3.919144e-06, 3.912474e-06, 3.925021e-06, 
    3.91618e-06, 3.955569e-06, 3.967416e-06, 4.023078e-06, 4.000189e-06, 
    4.036646e-06, 4.003885e-06, 4.009681e-06, 4.037837e-06, 4.005653e-06, 
    4.07621e-06, 4.028308e-06, 4.117502e-06, 4.069433e-06, 4.120524e-06, 
    4.111224e-06, 4.126627e-06, 4.140446e-06, 4.157862e-06, 4.19009e-06, 
    4.182617e-06, 4.209637e-06, 3.937575e-06, 3.953644e-06, 3.952229e-06, 
    3.969077e-06, 3.981559e-06, 4.008678e-06, 4.05236e-06, 4.035907e-06, 
    4.066137e-06, 4.072218e-06, 4.026302e-06, 4.054464e-06, 3.964417e-06, 
    3.978898e-06, 3.970274e-06, 3.938841e-06, 4.039694e-06, 3.987783e-06, 
    4.083895e-06, 4.055585e-06, 4.138474e-06, 4.09715e-06, 4.178505e-06, 
    4.213517e-06, 4.246598e-06, 4.285412e-06, 3.962428e-06, 3.951494e-06, 
    3.971083e-06, 3.99826e-06, 4.023558e-06, 4.057309e-06, 4.06077e-06, 
    4.06711e-06, 4.083556e-06, 4.097409e-06, 4.069115e-06, 4.100884e-06, 
    3.98226e-06, 4.044216e-06, 3.947364e-06, 3.976408e-06, 3.996656e-06, 
    3.987768e-06, 4.034029e-06, 4.04497e-06, 4.089573e-06, 4.066487e-06, 
    4.204862e-06, 4.143367e-06, 4.315081e-06, 4.266758e-06, 3.947678e-06, 
    3.962391e-06, 4.013803e-06, 3.989302e-06, 4.059567e-06, 4.076953e-06, 
    4.091113e-06, 4.109248e-06, 4.111209e-06, 4.121974e-06, 4.10434e-06, 
    4.121277e-06, 4.05738e-06, 4.085875e-06, 4.007912e-06, 4.026821e-06, 
    4.018116e-06, 4.008579e-06, 4.03805e-06, 4.06956e-06, 4.070235e-06, 
    4.080365e-06, 4.108972e-06, 4.059853e-06, 4.212829e-06, 4.118032e-06, 
    3.978465e-06, 4.006934e-06, 4.011009e-06, 3.999964e-06, 4.075208e-06, 
    4.047866e-06, 4.121712e-06, 4.101691e-06, 4.134519e-06, 4.118191e-06, 
    4.11579e-06, 4.09487e-06, 4.081871e-06, 4.049118e-06, 4.022563e-06, 
    4.001565e-06, 4.006443e-06, 4.029524e-06, 4.071491e-06, 4.111386e-06, 
    4.102631e-06, 4.13202e-06, 4.054452e-06, 4.086891e-06, 4.074338e-06, 
    4.107108e-06, 4.03547e-06, 4.096433e-06, 4.019958e-06, 4.026635e-06, 
    4.047325e-06, 4.089095e-06, 4.098366e-06, 4.108274e-06, 4.102159e-06, 
    4.07256e-06, 4.067721e-06, 4.046821e-06, 4.04106e-06, 4.025181e-06, 
    4.012058e-06, 4.024047e-06, 4.036657e-06, 4.072572e-06, 4.10507e-06, 
    4.140642e-06, 4.149371e-06, 4.19116e-06, 4.157125e-06, 4.213359e-06, 
    4.165525e-06, 4.248496e-06, 4.099981e-06, 4.164124e-06, 4.048268e-06, 
    4.060674e-06, 4.083159e-06, 4.134956e-06, 4.106954e-06, 4.139712e-06, 
    4.067531e-06, 4.030322e-06, 4.020722e-06, 4.00284e-06, 4.021132e-06, 
    4.019642e-06, 4.03718e-06, 4.03154e-06, 4.073768e-06, 4.051059e-06, 
    4.11573e-06, 4.139453e-06, 4.206801e-06, 4.248344e-06, 4.290835e-06, 
    4.309658e-06, 4.315395e-06, 4.317794e-06,
  4.120483e-06, 4.158956e-06, 4.15146e-06, 4.182609e-06, 4.165313e-06, 
    4.185733e-06, 4.128266e-06, 4.160488e-06, 4.139901e-06, 4.123937e-06, 
    4.243442e-06, 4.184002e-06, 4.30569e-06, 4.267406e-06, 4.36395e-06, 
    4.29972e-06, 4.376968e-06, 4.362088e-06, 4.406957e-06, 4.394076e-06, 
    4.451762e-06, 4.412911e-06, 4.481835e-06, 4.442465e-06, 4.448611e-06, 
    4.411633e-06, 4.195923e-06, 4.236016e-06, 4.193555e-06, 4.199257e-06, 
    4.196697e-06, 4.16567e-06, 4.150086e-06, 4.11755e-06, 4.123445e-06, 
    4.147347e-06, 4.201822e-06, 4.183283e-06, 4.230093e-06, 4.229032e-06, 
    4.281491e-06, 4.257793e-06, 4.346521e-06, 4.321195e-06, 4.394613e-06, 
    4.376082e-06, 4.393742e-06, 4.388382e-06, 4.393812e-06, 4.366652e-06, 
    4.378277e-06, 4.354421e-06, 4.262226e-06, 4.289203e-06, 4.209032e-06, 
    4.161247e-06, 4.129676e-06, 4.107358e-06, 4.110509e-06, 4.11652e-06, 
    4.147487e-06, 4.176722e-06, 4.199081e-06, 4.214075e-06, 4.22888e-06, 
    4.273878e-06, 4.297803e-06, 4.351654e-06, 4.341905e-06, 4.358426e-06, 
    4.374241e-06, 4.400869e-06, 4.39648e-06, 4.408235e-06, 4.357989e-06, 
    4.391346e-06, 4.336358e-06, 4.351358e-06, 4.232916e-06, 4.18828e-06, 
    4.169395e-06, 4.152901e-06, 4.112933e-06, 4.140511e-06, 4.129627e-06, 
    4.155545e-06, 4.172064e-06, 4.163889e-06, 4.214486e-06, 4.194774e-06, 
    4.299223e-06, 4.254052e-06, 4.372395e-06, 4.343905e-06, 4.379239e-06, 
    4.361188e-06, 4.392145e-06, 4.364278e-06, 4.412615e-06, 4.423181e-06, 
    4.415959e-06, 4.443738e-06, 4.362736e-06, 4.393743e-06, 4.16366e-06, 
    4.164993e-06, 4.171204e-06, 4.143943e-06, 4.142278e-06, 4.117388e-06, 
    4.13953e-06, 4.14898e-06, 4.173022e-06, 4.187282e-06, 4.200862e-06, 
    4.230811e-06, 4.264404e-06, 4.311633e-06, 4.345748e-06, 4.368704e-06, 
    4.354619e-06, 4.367053e-06, 4.353155e-06, 4.34665e-06, 4.419221e-06, 
    4.378386e-06, 4.439736e-06, 4.436328e-06, 4.408515e-06, 4.436712e-06, 
    4.165929e-06, 4.158263e-06, 4.131712e-06, 4.152482e-06, 4.114683e-06, 
    4.135818e-06, 4.147998e-06, 4.195187e-06, 4.205594e-06, 4.215259e-06, 
    4.234385e-06, 4.259004e-06, 4.30239e-06, 4.340346e-06, 4.375162e-06, 
    4.372605e-06, 4.373505e-06, 4.381304e-06, 4.362002e-06, 4.384478e-06, 
    4.388257e-06, 4.37838e-06, 4.435872e-06, 4.419403e-06, 4.436256e-06, 
    4.425528e-06, 4.160754e-06, 4.173662e-06, 4.166684e-06, 4.179811e-06, 
    4.170561e-06, 4.211784e-06, 4.224189e-06, 4.282512e-06, 4.258518e-06, 
    4.296739e-06, 4.262391e-06, 4.268466e-06, 4.297991e-06, 4.264243e-06, 
    4.338249e-06, 4.287997e-06, 4.381607e-06, 4.331138e-06, 4.384781e-06, 
    4.375011e-06, 4.391194e-06, 4.405717e-06, 4.424028e-06, 4.45793e-06, 
    4.450066e-06, 4.478503e-06, 4.192947e-06, 4.209768e-06, 4.208284e-06, 
    4.225925e-06, 4.238999e-06, 4.267414e-06, 4.313219e-06, 4.295961e-06, 
    4.327673e-06, 4.334056e-06, 4.285889e-06, 4.315427e-06, 4.221047e-06, 
    4.236215e-06, 4.227179e-06, 4.194273e-06, 4.299936e-06, 4.245521e-06, 
    4.346314e-06, 4.316602e-06, 4.403645e-06, 4.360233e-06, 4.445741e-06, 
    4.482592e-06, 4.517432e-06, 4.558353e-06, 4.218964e-06, 4.207515e-06, 
    4.228025e-06, 4.256499e-06, 4.283013e-06, 4.318411e-06, 4.322042e-06, 
    4.328695e-06, 4.345957e-06, 4.360501e-06, 4.330802e-06, 4.364151e-06, 
    4.23974e-06, 4.304678e-06, 4.203193e-06, 4.233607e-06, 4.254817e-06, 
    4.245504e-06, 4.293991e-06, 4.305465e-06, 4.352276e-06, 4.32804e-06, 
    4.473482e-06, 4.408791e-06, 4.589652e-06, 4.538682e-06, 4.20352e-06, 
    4.218924e-06, 4.272788e-06, 4.24711e-06, 4.32078e-06, 4.339026e-06, 
    4.35389e-06, 4.372937e-06, 4.374995e-06, 4.386306e-06, 4.367781e-06, 
    4.385573e-06, 4.318487e-06, 4.348392e-06, 4.26661e-06, 4.286434e-06, 
    4.277307e-06, 4.26731e-06, 4.298207e-06, 4.331268e-06, 4.331975e-06, 
    4.342608e-06, 4.372658e-06, 4.321079e-06, 4.481875e-06, 4.382173e-06, 
    4.235757e-06, 4.26559e-06, 4.269858e-06, 4.258281e-06, 4.337195e-06, 
    4.308505e-06, 4.38603e-06, 4.364998e-06, 4.399488e-06, 4.38233e-06, 
    4.379809e-06, 4.357836e-06, 4.344188e-06, 4.309818e-06, 4.28197e-06, 
    4.259959e-06, 4.265071e-06, 4.289269e-06, 4.333295e-06, 4.375182e-06, 
    4.365987e-06, 4.396861e-06, 4.315414e-06, 4.34946e-06, 4.336283e-06, 
    4.370689e-06, 4.295503e-06, 4.359486e-06, 4.279237e-06, 4.286238e-06, 
    4.307937e-06, 4.351776e-06, 4.361507e-06, 4.371914e-06, 4.36549e-06, 
    4.334416e-06, 4.329336e-06, 4.307408e-06, 4.301366e-06, 4.284713e-06, 
    4.270956e-06, 4.283525e-06, 4.296749e-06, 4.334428e-06, 4.368549e-06, 
    4.405925e-06, 4.415099e-06, 4.459062e-06, 4.423258e-06, 4.482434e-06, 
    4.432099e-06, 4.51944e-06, 4.363208e-06, 4.430619e-06, 4.308925e-06, 
    4.321941e-06, 4.345542e-06, 4.399951e-06, 4.370527e-06, 4.404948e-06, 
    4.329137e-06, 4.290107e-06, 4.280039e-06, 4.261296e-06, 4.280468e-06, 
    4.278907e-06, 4.297295e-06, 4.291381e-06, 4.335683e-06, 4.311853e-06, 
    4.379746e-06, 4.404676e-06, 4.475519e-06, 4.519275e-06, 4.564069e-06, 
    4.583927e-06, 4.589982e-06, 4.592514e-06,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOBCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNODSTMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOINTABS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMCL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOOCMSL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWDP =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWICE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOWLIQ =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_DEPTH =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SINKS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SNOW_SOURCES =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1C =
  5.778243, 5.778224, 5.778227, 5.778212, 5.778221, 5.778211, 5.778239, 
    5.778223, 5.778234, 5.778241, 5.778182, 5.778212, 5.778152, 5.77817, 
    5.778123, 5.778154, 5.778117, 5.778124, 5.778102, 5.778109, 5.778081, 
    5.7781, 5.778067, 5.778086, 5.778082, 5.7781, 5.778205, 5.778186, 
    5.778207, 5.778204, 5.778205, 5.778221, 5.778228, 5.778244, 5.778242, 
    5.77823, 5.778203, 5.778212, 5.778189, 5.778189, 5.778163, 5.778175, 
    5.778132, 5.778144, 5.778109, 5.778118, 5.778109, 5.778111, 5.778109, 
    5.778122, 5.778116, 5.778128, 5.778173, 5.77816, 5.778199, 5.778223, 
    5.778238, 5.77825, 5.778248, 5.778245, 5.77823, 5.778215, 5.778204, 
    5.778196, 5.778189, 5.778167, 5.778155, 5.778129, 5.778134, 5.778126, 
    5.778118, 5.778106, 5.778108, 5.778102, 5.778126, 5.77811, 5.778137, 
    5.77813, 5.778187, 5.778209, 5.778219, 5.778227, 5.778247, 5.778233, 
    5.778238, 5.778225, 5.778217, 5.778222, 5.778196, 5.778206, 5.778155, 
    5.778177, 5.778119, 5.778133, 5.778116, 5.778125, 5.77811, 5.778123, 
    5.7781, 5.778095, 5.778098, 5.778085, 5.778124, 5.778109, 5.778222, 
    5.778221, 5.778218, 5.778231, 5.778232, 5.778244, 5.778234, 5.778229, 
    5.778217, 5.77821, 5.778203, 5.778188, 5.778172, 5.778149, 5.778132, 
    5.778121, 5.778128, 5.778122, 5.778129, 5.778131, 5.778097, 5.778116, 
    5.778087, 5.778089, 5.778102, 5.778088, 5.77822, 5.778224, 5.778237, 
    5.778227, 5.778246, 5.778235, 5.778229, 5.778206, 5.778201, 5.778196, 
    5.778186, 5.778174, 5.778153, 5.778135, 5.778118, 5.778119, 5.778119, 
    5.778115, 5.778124, 5.778113, 5.778111, 5.778116, 5.778089, 5.778097, 
    5.778089, 5.778094, 5.778223, 5.778216, 5.77822, 5.778214, 5.778218, 
    5.778198, 5.778192, 5.778163, 5.778175, 5.778156, 5.778173, 5.77817, 
    5.778155, 5.778172, 5.778136, 5.77816, 5.778115, 5.778139, 5.778113, 
    5.778118, 5.77811, 5.778103, 5.778094, 5.778078, 5.778082, 5.778069, 
    5.778207, 5.778199, 5.778199, 5.778191, 5.778184, 5.77817, 5.778148, 
    5.778156, 5.778141, 5.778138, 5.778161, 5.778147, 5.778193, 5.778186, 
    5.77819, 5.778206, 5.778154, 5.778181, 5.778132, 5.778146, 5.778104, 
    5.778125, 5.778084, 5.778066, 5.77805, 5.77803, 5.778194, 5.7782, 
    5.77819, 5.778176, 5.778162, 5.778145, 5.778143, 5.778141, 5.778132, 
    5.778125, 5.77814, 5.778123, 5.778184, 5.778152, 5.778202, 5.778187, 
    5.778176, 5.778181, 5.778157, 5.778152, 5.778129, 5.778141, 5.778071, 
    5.778102, 5.778016, 5.77804, 5.778202, 5.778194, 5.778168, 5.77818, 
    5.778144, 5.778135, 5.778128, 5.778119, 5.778118, 5.778112, 5.778121, 
    5.778113, 5.778145, 5.778131, 5.778171, 5.778161, 5.778165, 5.778171, 
    5.778155, 5.778139, 5.778139, 5.778134, 5.778119, 5.778144, 5.778067, 
    5.778114, 5.778186, 5.778171, 5.778169, 5.778175, 5.778136, 5.77815, 
    5.778113, 5.778123, 5.778106, 5.778114, 5.778116, 5.778126, 5.778133, 
    5.77815, 5.778163, 5.778174, 5.778172, 5.77816, 5.778138, 5.778118, 
    5.778122, 5.778108, 5.778147, 5.778131, 5.778137, 5.77812, 5.778157, 
    5.778125, 5.778164, 5.778161, 5.778151, 5.778129, 5.778124, 5.77812, 
    5.778122, 5.778138, 5.77814, 5.778151, 5.778154, 5.778162, 5.778169, 
    5.778162, 5.778156, 5.778138, 5.778121, 5.778103, 5.778099, 5.778078, 
    5.778095, 5.778067, 5.77809, 5.778049, 5.778124, 5.778091, 5.77815, 
    5.778144, 5.778132, 5.778106, 5.77812, 5.778103, 5.77814, 5.778159, 
    5.778164, 5.778173, 5.778164, 5.778165, 5.778156, 5.778159, 5.778137, 
    5.778149, 5.778116, 5.778104, 5.77807, 5.778049, 5.778028, 5.778018, 
    5.778016, 5.778014 ;

 SOIL1C_TO_SOIL2C =
  3.096875e-08, 3.110524e-08, 3.107871e-08, 3.11888e-08, 3.112773e-08, 
    3.119982e-08, 3.099642e-08, 3.111066e-08, 3.103774e-08, 3.098104e-08, 
    3.140244e-08, 3.119371e-08, 3.161931e-08, 3.148617e-08, 3.182064e-08, 
    3.159859e-08, 3.186542e-08, 3.181424e-08, 3.196829e-08, 3.192416e-08, 
    3.212118e-08, 3.198866e-08, 3.222333e-08, 3.208954e-08, 3.211046e-08, 
    3.198429e-08, 3.123573e-08, 3.137646e-08, 3.122739e-08, 3.124745e-08, 
    3.123845e-08, 3.112899e-08, 3.107383e-08, 3.095832e-08, 3.097929e-08, 
    3.106413e-08, 3.125648e-08, 3.119119e-08, 3.135575e-08, 3.135203e-08, 
    3.153524e-08, 3.145264e-08, 3.176059e-08, 3.167306e-08, 3.1926e-08, 
    3.186239e-08, 3.192301e-08, 3.190463e-08, 3.192325e-08, 3.182996e-08, 
    3.186993e-08, 3.178783e-08, 3.14681e-08, 3.156207e-08, 3.128183e-08, 
    3.111333e-08, 3.100143e-08, 3.092203e-08, 3.093325e-08, 3.095465e-08, 
    3.106463e-08, 3.116804e-08, 3.124685e-08, 3.129956e-08, 3.13515e-08, 
    3.150871e-08, 3.159194e-08, 3.177828e-08, 3.174466e-08, 3.180163e-08, 
    3.185606e-08, 3.194744e-08, 3.19324e-08, 3.197266e-08, 3.180013e-08, 
    3.191479e-08, 3.172551e-08, 3.177728e-08, 3.136559e-08, 3.12088e-08, 
    3.114214e-08, 3.108381e-08, 3.094188e-08, 3.103989e-08, 3.100126e-08, 
    3.109318e-08, 3.115159e-08, 3.11227e-08, 3.1301e-08, 3.123168e-08, 
    3.159687e-08, 3.143957e-08, 3.184971e-08, 3.175156e-08, 3.187323e-08, 
    3.181115e-08, 3.191753e-08, 3.182179e-08, 3.198764e-08, 3.202375e-08, 
    3.199908e-08, 3.209388e-08, 3.181648e-08, 3.192301e-08, 3.112189e-08, 
    3.11266e-08, 3.114856e-08, 3.105206e-08, 3.104616e-08, 3.095775e-08, 
    3.103642e-08, 3.106992e-08, 3.115498e-08, 3.120529e-08, 3.125311e-08, 
    3.135826e-08, 3.14757e-08, 3.163993e-08, 3.175792e-08, 3.183702e-08, 
    3.178852e-08, 3.183134e-08, 3.178347e-08, 3.176104e-08, 3.201022e-08, 
    3.18703e-08, 3.208025e-08, 3.206863e-08, 3.197361e-08, 3.206994e-08, 
    3.112991e-08, 3.11028e-08, 3.100867e-08, 3.108233e-08, 3.094812e-08, 
    3.102324e-08, 3.106644e-08, 3.123312e-08, 3.126975e-08, 3.130371e-08, 
    3.137079e-08, 3.145686e-08, 3.160787e-08, 3.173927e-08, 3.185923e-08, 
    3.185044e-08, 3.185353e-08, 3.188033e-08, 3.181395e-08, 3.189123e-08, 
    3.190419e-08, 3.187028e-08, 3.206707e-08, 3.201085e-08, 3.206839e-08, 
    3.203178e-08, 3.111161e-08, 3.115724e-08, 3.113258e-08, 3.117894e-08, 
    3.114628e-08, 3.12915e-08, 3.133503e-08, 3.153878e-08, 3.145517e-08, 
    3.158825e-08, 3.146869e-08, 3.148987e-08, 3.159258e-08, 3.147515e-08, 
    3.173202e-08, 3.155786e-08, 3.188137e-08, 3.170744e-08, 3.189227e-08, 
    3.185871e-08, 3.191428e-08, 3.196404e-08, 3.202665e-08, 3.214218e-08, 
    3.211543e-08, 3.221205e-08, 3.122525e-08, 3.128442e-08, 3.127921e-08, 
    3.134114e-08, 3.138694e-08, 3.148621e-08, 3.164543e-08, 3.158556e-08, 
    3.169548e-08, 3.171755e-08, 3.155055e-08, 3.165308e-08, 3.132402e-08, 
    3.137718e-08, 3.134553e-08, 3.122991e-08, 3.159935e-08, 3.140974e-08, 
    3.175987e-08, 3.165716e-08, 3.195694e-08, 3.180785e-08, 3.21007e-08, 
    3.222589e-08, 3.234373e-08, 3.248143e-08, 3.131672e-08, 3.127651e-08, 
    3.134851e-08, 3.144811e-08, 3.154054e-08, 3.166342e-08, 3.1676e-08, 
    3.169901e-08, 3.175865e-08, 3.180878e-08, 3.170629e-08, 3.182135e-08, 
    3.13895e-08, 3.161581e-08, 3.12613e-08, 3.136804e-08, 3.144224e-08, 
    3.140969e-08, 3.157871e-08, 3.161855e-08, 3.178043e-08, 3.169675e-08, 
    3.219499e-08, 3.197454e-08, 3.25863e-08, 3.241533e-08, 3.126246e-08, 
    3.131658e-08, 3.150493e-08, 3.141531e-08, 3.167163e-08, 3.173471e-08, 
    3.178601e-08, 3.185157e-08, 3.185865e-08, 3.18975e-08, 3.183384e-08, 
    3.189498e-08, 3.166368e-08, 3.176704e-08, 3.148341e-08, 3.155244e-08, 
    3.152068e-08, 3.148585e-08, 3.159336e-08, 3.17079e-08, 3.171035e-08, 
    3.174708e-08, 3.185056e-08, 3.167266e-08, 3.222342e-08, 3.188327e-08, 
    3.13756e-08, 3.147983e-08, 3.149473e-08, 3.145435e-08, 3.172839e-08, 
    3.162909e-08, 3.189655e-08, 3.182427e-08, 3.194271e-08, 3.188385e-08, 
    3.187519e-08, 3.17996e-08, 3.175254e-08, 3.163364e-08, 3.153691e-08, 
    3.14602e-08, 3.147804e-08, 3.15623e-08, 3.171491e-08, 3.185929e-08, 
    3.182766e-08, 3.193371e-08, 3.165304e-08, 3.177072e-08, 3.172524e-08, 
    3.184384e-08, 3.158397e-08, 3.180524e-08, 3.15274e-08, 3.155176e-08, 
    3.162712e-08, 3.17787e-08, 3.181225e-08, 3.184805e-08, 3.182596e-08, 
    3.171878e-08, 3.170123e-08, 3.162529e-08, 3.160432e-08, 3.154646e-08, 
    3.149856e-08, 3.154232e-08, 3.158829e-08, 3.171883e-08, 3.183648e-08, 
    3.196475e-08, 3.199614e-08, 3.2146e-08, 3.2024e-08, 3.222532e-08, 
    3.205414e-08, 3.235047e-08, 3.181808e-08, 3.204912e-08, 3.163055e-08, 
    3.167564e-08, 3.17572e-08, 3.194427e-08, 3.184329e-08, 3.19614e-08, 
    3.170054e-08, 3.15652e-08, 3.15302e-08, 3.146487e-08, 3.153169e-08, 
    3.152625e-08, 3.159019e-08, 3.156965e-08, 3.172316e-08, 3.16407e-08, 
    3.187497e-08, 3.196046e-08, 3.220192e-08, 3.234994e-08, 3.250063e-08, 
    3.256716e-08, 3.25874e-08, 3.259587e-08 ;

 SOIL1C_TO_SOIL3C =
  3.673241e-10, 3.689436e-10, 3.686288e-10, 3.699351e-10, 3.692105e-10, 
    3.700658e-10, 3.676524e-10, 3.690079e-10, 3.681426e-10, 3.674699e-10, 
    3.724701e-10, 3.699933e-10, 3.750434e-10, 3.734636e-10, 3.774324e-10, 
    3.747975e-10, 3.779637e-10, 3.773565e-10, 3.791844e-10, 3.786607e-10, 
    3.809987e-10, 3.794261e-10, 3.822108e-10, 3.806231e-10, 3.808715e-10, 
    3.793742e-10, 3.704919e-10, 3.721617e-10, 3.703929e-10, 3.70631e-10, 
    3.705242e-10, 3.692254e-10, 3.685708e-10, 3.672004e-10, 3.674492e-10, 
    3.684558e-10, 3.707381e-10, 3.699634e-10, 3.71916e-10, 3.718719e-10, 
    3.740458e-10, 3.730656e-10, 3.767198e-10, 3.756812e-10, 3.786826e-10, 
    3.779277e-10, 3.786471e-10, 3.78429e-10, 3.786499e-10, 3.775429e-10, 
    3.780172e-10, 3.770431e-10, 3.732492e-10, 3.743641e-10, 3.710389e-10, 
    3.690396e-10, 3.677119e-10, 3.667697e-10, 3.669029e-10, 3.671568e-10, 
    3.684617e-10, 3.696887e-10, 3.706238e-10, 3.712493e-10, 3.718656e-10, 
    3.73731e-10, 3.747185e-10, 3.769297e-10, 3.765308e-10, 3.772067e-10, 
    3.778526e-10, 3.789369e-10, 3.787585e-10, 3.792362e-10, 3.771889e-10, 
    3.785495e-10, 3.763035e-10, 3.769177e-10, 3.720328e-10, 3.701724e-10, 
    3.693814e-10, 3.686893e-10, 3.670053e-10, 3.681682e-10, 3.677098e-10, 
    3.688005e-10, 3.694935e-10, 3.691508e-10, 3.712664e-10, 3.704438e-10, 
    3.747771e-10, 3.729105e-10, 3.777773e-10, 3.766127e-10, 3.780564e-10, 
    3.773197e-10, 3.785821e-10, 3.77446e-10, 3.79414e-10, 3.798425e-10, 
    3.795497e-10, 3.806747e-10, 3.77383e-10, 3.786471e-10, 3.691412e-10, 
    3.691971e-10, 3.694575e-10, 3.683126e-10, 3.682426e-10, 3.671935e-10, 
    3.68127e-10, 3.685245e-10, 3.695337e-10, 3.701306e-10, 3.706981e-10, 
    3.719458e-10, 3.733393e-10, 3.75288e-10, 3.766882e-10, 3.776267e-10, 
    3.770512e-10, 3.775593e-10, 3.769913e-10, 3.767251e-10, 3.79682e-10, 
    3.780216e-10, 3.805129e-10, 3.803751e-10, 3.792476e-10, 3.803906e-10, 
    3.692363e-10, 3.689146e-10, 3.677977e-10, 3.686718e-10, 3.670793e-10, 
    3.679706e-10, 3.684832e-10, 3.70461e-10, 3.708956e-10, 3.712985e-10, 
    3.720944e-10, 3.731158e-10, 3.749076e-10, 3.764668e-10, 3.778902e-10, 
    3.777859e-10, 3.778226e-10, 3.781406e-10, 3.77353e-10, 3.782699e-10, 
    3.784238e-10, 3.780214e-10, 3.803566e-10, 3.796894e-10, 3.803721e-10, 
    3.799377e-10, 3.690192e-10, 3.695605e-10, 3.69268e-10, 3.69818e-10, 
    3.694305e-10, 3.711536e-10, 3.716702e-10, 3.740878e-10, 3.730957e-10, 
    3.746748e-10, 3.732561e-10, 3.735075e-10, 3.747262e-10, 3.733328e-10, 
    3.763807e-10, 3.743142e-10, 3.78153e-10, 3.76089e-10, 3.782823e-10, 
    3.778841e-10, 3.785434e-10, 3.791339e-10, 3.798769e-10, 3.812478e-10, 
    3.809304e-10, 3.820769e-10, 3.703675e-10, 3.710696e-10, 3.710078e-10, 
    3.717426e-10, 3.722861e-10, 3.73464e-10, 3.753533e-10, 3.746428e-10, 
    3.759472e-10, 3.76209e-10, 3.742275e-10, 3.75444e-10, 3.715395e-10, 
    3.721703e-10, 3.717948e-10, 3.704229e-10, 3.748065e-10, 3.725567e-10, 
    3.767113e-10, 3.754924e-10, 3.790497e-10, 3.772805e-10, 3.807556e-10, 
    3.822411e-10, 3.836396e-10, 3.852736e-10, 3.714528e-10, 3.709758e-10, 
    3.7183e-10, 3.730119e-10, 3.741087e-10, 3.755667e-10, 3.75716e-10, 
    3.759891e-10, 3.766967e-10, 3.772916e-10, 3.760754e-10, 3.774408e-10, 
    3.723165e-10, 3.750018e-10, 3.707954e-10, 3.720619e-10, 3.729423e-10, 
    3.725561e-10, 3.745617e-10, 3.750344e-10, 3.769552e-10, 3.759623e-10, 
    3.818744e-10, 3.792586e-10, 3.86518e-10, 3.844891e-10, 3.708091e-10, 
    3.714512e-10, 3.736862e-10, 3.726228e-10, 3.756641e-10, 3.764127e-10, 
    3.770214e-10, 3.777993e-10, 3.778834e-10, 3.783444e-10, 3.77589e-10, 
    3.783145e-10, 3.755699e-10, 3.767964e-10, 3.734308e-10, 3.742499e-10, 
    3.738731e-10, 3.734597e-10, 3.747355e-10, 3.760945e-10, 3.761237e-10, 
    3.765595e-10, 3.777874e-10, 3.756764e-10, 3.822119e-10, 3.781755e-10, 
    3.721515e-10, 3.733883e-10, 3.735651e-10, 3.730859e-10, 3.763377e-10, 
    3.751594e-10, 3.783331e-10, 3.774754e-10, 3.788808e-10, 3.781824e-10, 
    3.780797e-10, 3.771827e-10, 3.766243e-10, 3.752134e-10, 3.740656e-10, 
    3.731555e-10, 3.733671e-10, 3.743668e-10, 3.761777e-10, 3.778909e-10, 
    3.775157e-10, 3.78774e-10, 3.754436e-10, 3.7684e-10, 3.763002e-10, 
    3.777077e-10, 3.74624e-10, 3.772496e-10, 3.739528e-10, 3.742419e-10, 
    3.75136e-10, 3.769347e-10, 3.773327e-10, 3.777576e-10, 3.774955e-10, 
    3.762237e-10, 3.760154e-10, 3.751143e-10, 3.748655e-10, 3.741789e-10, 
    3.736105e-10, 3.741298e-10, 3.746752e-10, 3.762243e-10, 3.776203e-10, 
    3.791423e-10, 3.795149e-10, 3.812932e-10, 3.798454e-10, 3.822344e-10, 
    3.802031e-10, 3.837195e-10, 3.774019e-10, 3.801436e-10, 3.751768e-10, 
    3.757118e-10, 3.766795e-10, 3.788994e-10, 3.777011e-10, 3.791026e-10, 
    3.760072e-10, 3.744013e-10, 3.739859e-10, 3.732108e-10, 3.740036e-10, 
    3.739392e-10, 3.746979e-10, 3.744541e-10, 3.762757e-10, 3.752972e-10, 
    3.78077e-10, 3.790915e-10, 3.819567e-10, 3.837132e-10, 3.855014e-10, 
    3.862909e-10, 3.865312e-10, 3.866316e-10 ;

 SOIL1C_vr =
  19.98124, 19.98119, 19.9812, 19.98116, 19.98118, 19.98115, 19.98123, 
    19.98119, 19.98121, 19.98124, 19.98108, 19.98116, 19.981, 19.98104, 
    19.98092, 19.981, 19.9809, 19.98092, 19.98086, 19.98088, 19.98081, 
    19.98086, 19.98077, 19.98082, 19.98081, 19.98086, 19.98114, 19.98109, 
    19.98114, 19.98114, 19.98114, 19.98118, 19.9812, 19.98125, 19.98124, 
    19.9812, 19.98113, 19.98116, 19.98109, 19.9811, 19.98103, 19.98106, 
    19.98094, 19.98098, 19.98088, 19.9809, 19.98088, 19.98089, 19.98088, 
    19.98092, 19.9809, 19.98093, 19.98105, 19.98102, 19.98112, 19.98119, 
    19.98123, 19.98126, 19.98125, 19.98125, 19.9812, 19.98116, 19.98114, 
    19.98112, 19.9811, 19.98104, 19.98101, 19.98094, 19.98095, 19.98093, 
    19.98091, 19.98087, 19.98088, 19.98086, 19.98093, 19.98088, 19.98096, 
    19.98094, 19.98109, 19.98115, 19.98118, 19.9812, 19.98125, 19.98121, 
    19.98123, 19.98119, 19.98117, 19.98118, 19.98112, 19.98114, 19.981, 
    19.98106, 19.98091, 19.98095, 19.9809, 19.98092, 19.98088, 19.98092, 
    19.98086, 19.98084, 19.98085, 19.98082, 19.98092, 19.98088, 19.98118, 
    19.98118, 19.98117, 19.98121, 19.98121, 19.98125, 19.98122, 19.9812, 
    19.98117, 19.98115, 19.98113, 19.98109, 19.98105, 19.98099, 19.98094, 
    19.98091, 19.98093, 19.98092, 19.98093, 19.98094, 19.98085, 19.9809, 
    19.98082, 19.98083, 19.98086, 19.98083, 19.98118, 19.98119, 19.98123, 
    19.9812, 19.98125, 19.98122, 19.9812, 19.98114, 19.98113, 19.98112, 
    19.98109, 19.98106, 19.981, 19.98095, 19.98091, 19.98091, 19.98091, 
    19.9809, 19.98092, 19.98089, 19.98089, 19.9809, 19.98083, 19.98085, 
    19.98083, 19.98084, 19.98119, 19.98117, 19.98118, 19.98116, 19.98117, 
    19.98112, 19.9811, 19.98103, 19.98106, 19.98101, 19.98105, 19.98104, 
    19.981, 19.98105, 19.98095, 19.98102, 19.9809, 19.98096, 19.98089, 
    19.98091, 19.98088, 19.98087, 19.98084, 19.9808, 19.98081, 19.98077, 
    19.98114, 19.98112, 19.98112, 19.9811, 19.98108, 19.98104, 19.98099, 
    19.98101, 19.98097, 19.98096, 19.98102, 19.98098, 19.98111, 19.98109, 
    19.9811, 19.98114, 19.981, 19.98108, 19.98094, 19.98098, 19.98087, 
    19.98092, 19.98081, 19.98077, 19.98072, 19.98067, 19.98111, 19.98112, 
    19.9811, 19.98106, 19.98103, 19.98098, 19.98097, 19.98096, 19.98094, 
    19.98092, 19.98096, 19.98092, 19.98108, 19.981, 19.98113, 19.98109, 
    19.98106, 19.98108, 19.98101, 19.981, 19.98093, 19.98097, 19.98078, 
    19.98086, 19.98063, 19.9807, 19.98113, 19.98111, 19.98104, 19.98107, 
    19.98098, 19.98095, 19.98093, 19.98091, 19.98091, 19.98089, 19.98092, 
    19.98089, 19.98098, 19.98094, 19.98105, 19.98102, 19.98103, 19.98105, 
    19.981, 19.98096, 19.98096, 19.98095, 19.98091, 19.98098, 19.98077, 
    19.9809, 19.98109, 19.98105, 19.98104, 19.98106, 19.98096, 19.98099, 
    19.98089, 19.98092, 19.98087, 19.9809, 19.9809, 19.98093, 19.98095, 
    19.98099, 19.98103, 19.98106, 19.98105, 19.98102, 19.98096, 19.98091, 
    19.98092, 19.98088, 19.98098, 19.98094, 19.98096, 19.98091, 19.98101, 
    19.98092, 19.98103, 19.98102, 19.98099, 19.98094, 19.98092, 19.98091, 
    19.98092, 19.98096, 19.98096, 19.98099, 19.981, 19.98102, 19.98104, 
    19.98102, 19.98101, 19.98096, 19.98091, 19.98087, 19.98085, 19.9808, 
    19.98084, 19.98077, 19.98083, 19.98072, 19.98092, 19.98083, 19.98099, 
    19.98097, 19.98094, 19.98087, 19.98091, 19.98087, 19.98096, 19.98102, 
    19.98103, 19.98105, 19.98103, 19.98103, 19.98101, 19.98101, 19.98096, 
    19.98099, 19.9809, 19.98087, 19.98078, 19.98072, 19.98066, 19.98064, 
    19.98063, 19.98063,
  19.9833, 19.98323, 19.98325, 19.98319, 19.98322, 19.98319, 19.98328, 
    19.98323, 19.98326, 19.98329, 19.9831, 19.98319, 19.983, 19.98306, 
    19.9829, 19.98301, 19.98288, 19.98291, 19.98283, 19.98285, 19.98276, 
    19.98282, 19.98272, 19.98278, 19.98277, 19.98283, 19.98317, 19.98311, 
    19.98318, 19.98317, 19.98317, 19.98322, 19.98325, 19.9833, 19.98329, 
    19.98325, 19.98316, 19.98319, 19.98312, 19.98312, 19.98303, 19.98307, 
    19.98293, 19.98297, 19.98285, 19.98288, 19.98285, 19.98286, 19.98285, 
    19.9829, 19.98288, 19.98292, 19.98307, 19.98302, 19.98315, 19.98323, 
    19.98328, 19.98332, 19.98331, 19.9833, 19.98325, 19.9832, 19.98317, 
    19.98314, 19.98312, 19.98305, 19.98301, 19.98292, 19.98294, 19.98291, 
    19.98289, 19.98284, 19.98285, 19.98283, 19.98291, 19.98286, 19.98295, 
    19.98292, 19.98311, 19.98319, 19.98322, 19.98324, 19.98331, 19.98326, 
    19.98328, 19.98324, 19.98321, 19.98322, 19.98314, 19.98318, 19.98301, 
    19.98308, 19.98289, 19.98293, 19.98288, 19.98291, 19.98286, 19.9829, 
    19.98283, 19.98281, 19.98282, 19.98278, 19.9829, 19.98285, 19.98323, 
    19.98322, 19.98321, 19.98326, 19.98326, 19.9833, 19.98327, 19.98325, 
    19.98321, 19.98319, 19.98317, 19.98312, 19.98306, 19.98299, 19.98293, 
    19.98289, 19.98292, 19.9829, 19.98292, 19.98293, 19.98281, 19.98288, 
    19.98278, 19.98279, 19.98283, 19.98279, 19.98322, 19.98323, 19.98328, 
    19.98324, 19.98331, 19.98327, 19.98325, 19.98318, 19.98316, 19.98314, 
    19.98311, 19.98307, 19.983, 19.98294, 19.98289, 19.98289, 19.98289, 
    19.98288, 19.98291, 19.98287, 19.98286, 19.98288, 19.98279, 19.98281, 
    19.98279, 19.98281, 19.98323, 19.98321, 19.98322, 19.9832, 19.98322, 
    19.98315, 19.98313, 19.98303, 19.98307, 19.98301, 19.98306, 19.98306, 
    19.98301, 19.98306, 19.98294, 19.98302, 19.98287, 19.98295, 19.98287, 
    19.98289, 19.98286, 19.98284, 19.98281, 19.98275, 19.98277, 19.98272, 
    19.98318, 19.98315, 19.98315, 19.98312, 19.9831, 19.98306, 19.98298, 
    19.98301, 19.98296, 19.98295, 19.98303, 19.98298, 19.98313, 19.98311, 
    19.98312, 19.98318, 19.98301, 19.98309, 19.98293, 19.98298, 19.98284, 
    19.98291, 19.98277, 19.98272, 19.98266, 19.9826, 19.98314, 19.98315, 
    19.98312, 19.98307, 19.98303, 19.98298, 19.98297, 19.98296, 19.98293, 
    19.98291, 19.98296, 19.9829, 19.9831, 19.983, 19.98316, 19.98311, 
    19.98308, 19.98309, 19.98302, 19.983, 19.98292, 19.98296, 19.98273, 
    19.98283, 19.98255, 19.98263, 19.98316, 19.98314, 19.98305, 19.98309, 
    19.98297, 19.98294, 19.98292, 19.98289, 19.98289, 19.98287, 19.9829, 
    19.98287, 19.98298, 19.98293, 19.98306, 19.98303, 19.98304, 19.98306, 
    19.98301, 19.98295, 19.98295, 19.98294, 19.98289, 19.98297, 19.98272, 
    19.98287, 19.98311, 19.98306, 19.98305, 19.98307, 19.98294, 19.98299, 
    19.98287, 19.9829, 19.98285, 19.98287, 19.98288, 19.98291, 19.98293, 
    19.98299, 19.98303, 19.98307, 19.98306, 19.98302, 19.98295, 19.98289, 
    19.9829, 19.98285, 19.98298, 19.98293, 19.98295, 19.98289, 19.98301, 
    19.98291, 19.98304, 19.98303, 19.98299, 19.98292, 19.98291, 19.98289, 
    19.9829, 19.98295, 19.98296, 19.98299, 19.983, 19.98303, 19.98305, 
    19.98303, 19.98301, 19.98295, 19.98289, 19.98284, 19.98282, 19.98275, 
    19.98281, 19.98272, 19.9828, 19.98266, 19.9829, 19.9828, 19.98299, 
    19.98297, 19.98293, 19.98285, 19.98289, 19.98284, 19.98296, 19.98302, 
    19.98304, 19.98307, 19.98304, 19.98304, 19.98301, 19.98302, 19.98295, 
    19.98299, 19.98288, 19.98284, 19.98273, 19.98266, 19.98259, 19.98256, 
    19.98255, 19.98255,
  19.98426, 19.98419, 19.9842, 19.98414, 19.98418, 19.98414, 19.98424, 
    19.98418, 19.98422, 19.98425, 19.98404, 19.98414, 19.98392, 19.98399, 
    19.98382, 19.98394, 19.9838, 19.98383, 19.98375, 19.98377, 19.98367, 
    19.98374, 19.98362, 19.98368, 19.98368, 19.98374, 19.98412, 19.98405, 
    19.98413, 19.98411, 19.98412, 19.98417, 19.9842, 19.98426, 19.98425, 
    19.98421, 19.98411, 19.98414, 19.98406, 19.98406, 19.98397, 19.98401, 
    19.98385, 19.9839, 19.98377, 19.9838, 19.98377, 19.98378, 19.98377, 
    19.98382, 19.9838, 19.98384, 19.984, 19.98395, 19.9841, 19.98418, 
    19.98424, 19.98428, 19.98428, 19.98426, 19.98421, 19.98416, 19.98412, 
    19.98409, 19.98406, 19.98398, 19.98394, 19.98384, 19.98386, 19.98383, 
    19.9838, 19.98376, 19.98376, 19.98375, 19.98383, 19.98377, 19.98387, 
    19.98384, 19.98405, 19.98413, 19.98417, 19.9842, 19.98427, 19.98422, 
    19.98424, 19.98419, 19.98416, 19.98418, 19.98409, 19.98412, 19.98394, 
    19.98402, 19.98381, 19.98386, 19.9838, 19.98383, 19.98377, 19.98382, 
    19.98374, 19.98372, 19.98373, 19.98368, 19.98382, 19.98377, 19.98418, 
    19.98418, 19.98417, 19.98421, 19.98422, 19.98426, 19.98422, 19.98421, 
    19.98416, 19.98414, 19.98411, 19.98406, 19.984, 19.98391, 19.98385, 
    19.98381, 19.98384, 19.98382, 19.98384, 19.98385, 19.98373, 19.9838, 
    19.98369, 19.9837, 19.98374, 19.9837, 19.98417, 19.98419, 19.98424, 
    19.9842, 19.98427, 19.98423, 19.98421, 19.98412, 19.9841, 19.98409, 
    19.98405, 19.98401, 19.98393, 19.98386, 19.9838, 19.98381, 19.9838, 
    19.98379, 19.98383, 19.98379, 19.98378, 19.9838, 19.9837, 19.98372, 
    19.9837, 19.98372, 19.98418, 19.98416, 19.98417, 19.98415, 19.98417, 
    19.98409, 19.98407, 19.98397, 19.98401, 19.98394, 19.984, 19.98399, 
    19.98394, 19.984, 19.98387, 19.98396, 19.98379, 19.98388, 19.98379, 
    19.9838, 19.98377, 19.98375, 19.98372, 19.98366, 19.98367, 19.98362, 
    19.98413, 19.9841, 19.9841, 19.98407, 19.98404, 19.98399, 19.98391, 
    19.98394, 19.98389, 19.98388, 19.98396, 19.98391, 19.98408, 19.98405, 
    19.98406, 19.98412, 19.98393, 19.98403, 19.98385, 19.98391, 19.98375, 
    19.98383, 19.98368, 19.98362, 19.98356, 19.98349, 19.98408, 19.9841, 
    19.98406, 19.98401, 19.98396, 19.9839, 19.9839, 19.98388, 19.98385, 
    19.98383, 19.98388, 19.98382, 19.98404, 19.98393, 19.98411, 19.98405, 
    19.98401, 19.98403, 19.98395, 19.98392, 19.98384, 19.98388, 19.98363, 
    19.98374, 19.98343, 19.98352, 19.98411, 19.98408, 19.98398, 19.98403, 
    19.9839, 19.98387, 19.98384, 19.98381, 19.9838, 19.98378, 19.98382, 
    19.98378, 19.9839, 19.98385, 19.98399, 19.98396, 19.98397, 19.98399, 
    19.98394, 19.98388, 19.98388, 19.98386, 19.98381, 19.9839, 19.98362, 
    19.98379, 19.98405, 19.984, 19.98399, 19.98401, 19.98387, 19.98392, 
    19.98378, 19.98382, 19.98376, 19.98379, 19.9838, 19.98383, 19.98386, 
    19.98392, 19.98397, 19.98401, 19.984, 19.98395, 19.98388, 19.9838, 
    19.98382, 19.98376, 19.98391, 19.98385, 19.98387, 19.98381, 19.98394, 
    19.98383, 19.98397, 19.98396, 19.98392, 19.98384, 19.98383, 19.98381, 
    19.98382, 19.98387, 19.98388, 19.98392, 19.98393, 19.98396, 19.98399, 
    19.98396, 19.98394, 19.98387, 19.98381, 19.98375, 19.98373, 19.98366, 
    19.98372, 19.98362, 19.9837, 19.98355, 19.98382, 19.98371, 19.98392, 
    19.9839, 19.98385, 19.98376, 19.98381, 19.98375, 19.98388, 19.98395, 
    19.98397, 19.984, 19.98397, 19.98397, 19.98394, 19.98395, 19.98387, 
    19.98391, 19.9838, 19.98375, 19.98363, 19.98355, 19.98348, 19.98344, 
    19.98343, 19.98343,
  19.98501, 19.98494, 19.98495, 19.98489, 19.98492, 19.98489, 19.98499, 
    19.98493, 19.98497, 19.985, 19.98478, 19.98489, 19.98467, 19.98474, 
    19.98456, 19.98468, 19.98454, 19.98457, 19.98449, 19.98451, 19.98441, 
    19.98447, 19.98435, 19.98442, 19.98441, 19.98448, 19.98487, 19.98479, 
    19.98487, 19.98486, 19.98487, 19.98492, 19.98495, 19.98501, 19.985, 
    19.98496, 19.98486, 19.98489, 19.9848, 19.98481, 19.98471, 19.98475, 
    19.98459, 19.98464, 19.98451, 19.98454, 19.98451, 19.98452, 19.98451, 
    19.98456, 19.98454, 19.98458, 19.98475, 19.9847, 19.98484, 19.98493, 
    19.98499, 19.98503, 19.98503, 19.98501, 19.98496, 19.9849, 19.98486, 
    19.98483, 19.98481, 19.98472, 19.98468, 19.98458, 19.9846, 19.98457, 
    19.98454, 19.9845, 19.9845, 19.98448, 19.98457, 19.98451, 19.98461, 
    19.98458, 19.9848, 19.98488, 19.98492, 19.98495, 19.98502, 19.98497, 
    19.98499, 19.98494, 19.98491, 19.98493, 19.98483, 19.98487, 19.98468, 
    19.98476, 19.98455, 19.9846, 19.98454, 19.98457, 19.98451, 19.98456, 
    19.98448, 19.98446, 19.98447, 19.98442, 19.98456, 19.98451, 19.98493, 
    19.98492, 19.98491, 19.98496, 19.98497, 19.98501, 19.98497, 19.98495, 
    19.98491, 19.98488, 19.98486, 19.9848, 19.98474, 19.98466, 19.98459, 
    19.98455, 19.98458, 19.98456, 19.98458, 19.98459, 19.98446, 19.98454, 
    19.98443, 19.98443, 19.98448, 19.98443, 19.98492, 19.98494, 19.98499, 
    19.98495, 19.98502, 19.98498, 19.98495, 19.98487, 19.98485, 19.98483, 
    19.9848, 19.98475, 19.98467, 19.9846, 19.98454, 19.98455, 19.98454, 
    19.98453, 19.98457, 19.98453, 19.98452, 19.98454, 19.98443, 19.98446, 
    19.98443, 19.98445, 19.98493, 19.98491, 19.98492, 19.9849, 19.98491, 
    19.98484, 19.98482, 19.98471, 19.98475, 19.98468, 19.98475, 19.98474, 
    19.98468, 19.98474, 19.98461, 19.9847, 19.98453, 19.98462, 19.98453, 
    19.98454, 19.98451, 19.98449, 19.98446, 19.98439, 19.98441, 19.98436, 
    19.98487, 19.98484, 19.98484, 19.98481, 19.98479, 19.98474, 19.98465, 
    19.98468, 19.98463, 19.98462, 19.9847, 19.98465, 19.98482, 19.98479, 
    19.98481, 19.98487, 19.98468, 19.98478, 19.98459, 19.98465, 19.98449, 
    19.98457, 19.98442, 19.98435, 19.98429, 19.98422, 19.98483, 19.98485, 
    19.98481, 19.98476, 19.98471, 19.98464, 19.98464, 19.98462, 19.98459, 
    19.98457, 19.98462, 19.98456, 19.98479, 19.98467, 19.98485, 19.9848, 
    19.98476, 19.98478, 19.98469, 19.98467, 19.98458, 19.98463, 19.98437, 
    19.98448, 19.98416, 19.98425, 19.98485, 19.98483, 19.98473, 19.98477, 
    19.98464, 19.98461, 19.98458, 19.98455, 19.98454, 19.98452, 19.98456, 
    19.98452, 19.98464, 19.98459, 19.98474, 19.9847, 19.98472, 19.98474, 
    19.98468, 19.98462, 19.98462, 19.9846, 19.98455, 19.98464, 19.98435, 
    19.98453, 19.98479, 19.98474, 19.98473, 19.98475, 19.98461, 19.98466, 
    19.98452, 19.98456, 19.9845, 19.98453, 19.98453, 19.98457, 19.9846, 
    19.98466, 19.98471, 19.98475, 19.98474, 19.9847, 19.98462, 19.98454, 
    19.98456, 19.9845, 19.98465, 19.98459, 19.98461, 19.98455, 19.98469, 
    19.98457, 19.98471, 19.9847, 19.98466, 19.98458, 19.98457, 19.98455, 
    19.98456, 19.98462, 19.98462, 19.98466, 19.98467, 19.9847, 19.98473, 
    19.98471, 19.98468, 19.98462, 19.98455, 19.98449, 19.98447, 19.98439, 
    19.98446, 19.98435, 19.98444, 19.98429, 19.98456, 19.98444, 19.98466, 
    19.98464, 19.9846, 19.9845, 19.98455, 19.98449, 19.98462, 19.9847, 
    19.98471, 19.98475, 19.98471, 19.98472, 19.98468, 19.98469, 19.98461, 
    19.98466, 19.98453, 19.98449, 19.98436, 19.98429, 19.98421, 19.98417, 
    19.98416, 19.98416,
  19.98609, 19.98602, 19.98603, 19.98598, 19.98601, 19.98598, 19.98607, 
    19.98602, 19.98605, 19.98608, 19.98588, 19.98598, 19.98577, 19.98584, 
    19.98568, 19.98578, 19.98566, 19.98568, 19.98561, 19.98563, 19.98554, 
    19.9856, 19.98549, 19.98555, 19.98554, 19.9856, 19.98596, 19.98589, 
    19.98596, 19.98595, 19.98596, 19.98601, 19.98603, 19.98609, 19.98608, 
    19.98604, 19.98595, 19.98598, 19.9859, 19.9859, 19.98582, 19.98586, 
    19.98571, 19.98575, 19.98563, 19.98566, 19.98563, 19.98564, 19.98563, 
    19.98568, 19.98566, 19.98569, 19.98585, 19.9858, 19.98594, 19.98602, 
    19.98607, 19.98611, 19.9861, 19.98609, 19.98604, 19.98599, 19.98595, 
    19.98593, 19.9859, 19.98583, 19.98579, 19.9857, 19.98572, 19.98569, 
    19.98566, 19.98562, 19.98563, 19.98561, 19.98569, 19.98563, 19.98573, 
    19.9857, 19.9859, 19.98597, 19.986, 19.98603, 19.9861, 19.98605, 
    19.98607, 19.98603, 19.986, 19.98601, 19.98593, 19.98596, 19.98579, 
    19.98586, 19.98567, 19.98571, 19.98565, 19.98568, 19.98563, 19.98568, 
    19.9856, 19.98558, 19.98559, 19.98555, 19.98568, 19.98563, 19.98601, 
    19.98601, 19.986, 19.98605, 19.98605, 19.98609, 19.98605, 19.98604, 
    19.986, 19.98597, 19.98595, 19.9859, 19.98584, 19.98577, 19.98571, 
    19.98567, 19.98569, 19.98567, 19.9857, 19.98571, 19.98559, 19.98566, 
    19.98556, 19.98556, 19.98561, 19.98556, 19.98601, 19.98602, 19.98607, 
    19.98603, 19.9861, 19.98606, 19.98604, 19.98596, 19.98594, 19.98593, 
    19.98589, 19.98585, 19.98578, 19.98572, 19.98566, 19.98567, 19.98566, 
    19.98565, 19.98568, 19.98565, 19.98564, 19.98566, 19.98556, 19.98559, 
    19.98556, 19.98558, 19.98602, 19.986, 19.98601, 19.98598, 19.986, 
    19.98593, 19.98591, 19.98581, 19.98585, 19.98579, 19.98585, 19.98584, 
    19.98579, 19.98584, 19.98572, 19.98581, 19.98565, 19.98573, 19.98565, 
    19.98566, 19.98564, 19.98561, 19.98558, 19.98553, 19.98554, 19.98549, 
    19.98596, 19.98594, 19.98594, 19.98591, 19.98589, 19.98584, 19.98576, 
    19.98579, 19.98574, 19.98573, 19.98581, 19.98576, 19.98592, 19.98589, 
    19.98591, 19.98596, 19.98578, 19.98588, 19.98571, 19.98576, 19.98561, 
    19.98569, 19.98555, 19.98549, 19.98543, 19.98536, 19.98592, 19.98594, 
    19.9859, 19.98586, 19.98581, 19.98575, 19.98575, 19.98574, 19.98571, 
    19.98569, 19.98573, 19.98568, 19.98589, 19.98578, 19.98595, 19.9859, 
    19.98586, 19.98588, 19.98579, 19.98577, 19.9857, 19.98574, 19.9855, 
    19.98561, 19.98531, 19.9854, 19.98594, 19.98592, 19.98583, 19.98587, 
    19.98575, 19.98572, 19.9857, 19.98566, 19.98566, 19.98564, 19.98567, 
    19.98564, 19.98575, 19.9857, 19.98584, 19.98581, 19.98582, 19.98584, 
    19.98579, 19.98573, 19.98573, 19.98571, 19.98566, 19.98575, 19.98549, 
    19.98565, 19.98589, 19.98584, 19.98583, 19.98585, 19.98572, 19.98577, 
    19.98564, 19.98568, 19.98562, 19.98565, 19.98565, 19.98569, 19.98571, 
    19.98577, 19.98582, 19.98585, 19.98584, 19.9858, 19.98573, 19.98566, 
    19.98568, 19.98563, 19.98576, 19.9857, 19.98573, 19.98567, 19.98579, 
    19.98569, 19.98582, 19.98581, 19.98577, 19.9857, 19.98568, 19.98567, 
    19.98568, 19.98573, 19.98574, 19.98577, 19.98578, 19.98581, 19.98583, 
    19.98581, 19.98579, 19.98573, 19.98567, 19.98561, 19.9856, 19.98553, 
    19.98558, 19.98549, 19.98557, 19.98543, 19.98568, 19.98557, 19.98577, 
    19.98575, 19.98571, 19.98562, 19.98567, 19.98561, 19.98574, 19.9858, 
    19.98582, 19.98585, 19.98582, 19.98582, 19.98579, 19.9858, 19.98573, 
    19.98577, 19.98565, 19.98561, 19.9855, 19.98543, 19.98536, 19.98532, 
    19.98531, 19.98531,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N =
  0.7222804, 0.722278, 0.7222784, 0.7222765, 0.7222776, 0.7222763, 0.7222799, 
    0.7222779, 0.7222792, 0.7222801, 0.7222728, 0.7222764, 0.7222689, 
    0.7222713, 0.7222654, 0.7222693, 0.7222646, 0.7222655, 0.7222628, 
    0.7222636, 0.7222601, 0.7222624, 0.7222583, 0.7222607, 0.7222603, 
    0.7222626, 0.7222757, 0.7222732, 0.7222759, 0.7222755, 0.7222756, 
    0.7222776, 0.7222785, 0.7222806, 0.7222802, 0.7222787, 0.7222753, 
    0.7222764, 0.7222736, 0.7222736, 0.7222704, 0.7222719, 0.7222665, 
    0.722268, 0.7222636, 0.7222647, 0.7222636, 0.7222639, 0.7222636, 
    0.7222652, 0.7222645, 0.722266, 0.7222716, 0.72227, 0.7222749, 0.7222778, 
    0.7222798, 0.7222812, 0.722281, 0.7222806, 0.7222787, 0.7222769, 
    0.7222755, 0.7222745, 0.7222736, 0.7222709, 0.7222694, 0.7222661, 
    0.7222667, 0.7222657, 0.7222648, 0.7222632, 0.7222635, 0.7222627, 
    0.7222658, 0.7222638, 0.7222671, 0.7222662, 0.7222734, 0.7222762, 
    0.7222773, 0.7222784, 0.7222809, 0.7222791, 0.7222798, 0.7222782, 
    0.7222772, 0.7222777, 0.7222745, 0.7222757, 0.7222694, 0.7222721, 
    0.7222649, 0.7222666, 0.7222645, 0.7222656, 0.7222637, 0.7222654, 
    0.7222625, 0.7222618, 0.7222623, 0.7222606, 0.7222655, 0.7222636, 
    0.7222777, 0.7222776, 0.7222772, 0.7222789, 0.722279, 0.7222806, 
    0.7222792, 0.7222786, 0.7222771, 0.7222762, 0.7222754, 0.7222735, 
    0.7222715, 0.7222686, 0.7222665, 0.7222651, 0.722266, 0.7222652, 
    0.7222661, 0.7222664, 0.7222621, 0.7222645, 0.7222608, 0.7222611, 
    0.7222627, 0.722261, 0.7222775, 0.722278, 0.7222797, 0.7222784, 
    0.7222807, 0.7222794, 0.7222787, 0.7222757, 0.7222751, 0.7222745, 
    0.7222733, 0.7222718, 0.7222692, 0.7222669, 0.7222648, 0.7222649, 
    0.7222648, 0.7222643, 0.7222655, 0.7222642, 0.7222639, 0.7222645, 
    0.7222611, 0.7222621, 0.7222611, 0.7222617, 0.7222779, 0.722277, 
    0.7222775, 0.7222767, 0.7222773, 0.7222747, 0.7222739, 0.7222704, 
    0.7222719, 0.7222695, 0.7222716, 0.7222712, 0.7222694, 0.7222715, 
    0.722267, 0.72227, 0.7222643, 0.7222674, 0.7222642, 0.7222648, 0.7222638, 
    0.7222629, 0.7222618, 0.7222598, 0.7222602, 0.7222586, 0.7222759, 
    0.7222748, 0.7222749, 0.7222738, 0.7222731, 0.7222713, 0.7222685, 
    0.7222695, 0.7222676, 0.7222672, 0.7222701, 0.7222683, 0.7222741, 
    0.7222732, 0.7222738, 0.7222758, 0.7222693, 0.7222726, 0.7222665, 
    0.7222683, 0.722263, 0.7222657, 0.7222605, 0.7222583, 0.7222562, 
    0.7222538, 0.7222742, 0.722275, 0.7222737, 0.722272, 0.7222703, 
    0.7222682, 0.7222679, 0.7222676, 0.7222665, 0.7222656, 0.7222674, 
    0.7222654, 0.722273, 0.722269, 0.7222753, 0.7222733, 0.722272, 0.7222726, 
    0.7222697, 0.7222689, 0.7222661, 0.7222676, 0.7222589, 0.7222627, 
    0.722252, 0.722255, 0.7222752, 0.7222742, 0.722271, 0.7222725, 0.722268, 
    0.7222669, 0.722266, 0.7222649, 0.7222648, 0.7222641, 0.7222652, 
    0.7222641, 0.7222682, 0.7222664, 0.7222713, 0.7222701, 0.7222707, 
    0.7222713, 0.7222694, 0.7222674, 0.7222673, 0.7222667, 0.7222649, 
    0.722268, 0.7222583, 0.7222643, 0.7222732, 0.7222714, 0.7222711, 
    0.7222719, 0.722267, 0.7222688, 0.7222641, 0.7222654, 0.7222633, 
    0.7222643, 0.7222645, 0.7222658, 0.7222666, 0.7222687, 0.7222704, 
    0.7222717, 0.7222714, 0.72227, 0.7222673, 0.7222647, 0.7222653, 
    0.7222635, 0.7222683, 0.7222663, 0.7222671, 0.722265, 0.7222696, 
    0.7222657, 0.7222705, 0.7222701, 0.7222688, 0.7222661, 0.7222655, 
    0.7222649, 0.7222653, 0.7222672, 0.7222675, 0.7222688, 0.7222692, 
    0.7222703, 0.7222711, 0.7222703, 0.7222695, 0.7222672, 0.7222651, 
    0.7222629, 0.7222623, 0.7222597, 0.7222618, 0.7222583, 0.7222613, 
    0.7222561, 0.7222655, 0.7222614, 0.7222688, 0.722268, 0.7222666, 
    0.7222632, 0.722265, 0.7222629, 0.7222675, 0.7222699, 0.7222705, 
    0.7222717, 0.7222705, 0.7222706, 0.7222695, 0.7222698, 0.7222672, 
    0.7222686, 0.7222645, 0.722263, 0.7222587, 0.7222561, 0.7222535, 
    0.7222523, 0.722252, 0.7222518 ;

 SOIL1N_TNDNCY_VERT_TRANS =
  -1.027984e-20, 5.139921e-21, 2.055969e-20, -1.541976e-20, 1.541976e-20, 0, 
    2.055969e-20, 2.569961e-20, 2.006177e-36, 1.027984e-20, 2.055969e-20, 
    -5.139921e-21, 1.027984e-20, 2.569961e-20, -1.541976e-20, 5.139921e-21, 
    5.139921e-21, 5.139921e-21, -1.027984e-20, 2.006177e-36, -1.541976e-20, 
    -1.027984e-20, -1.541976e-20, -3.597945e-20, -5.139921e-21, 2.006177e-36, 
    -1.541976e-20, 0, -5.139921e-21, 5.139921e-21, -5.139921e-21, 
    -1.027984e-20, -1.541976e-20, -5.139921e-21, 1.027984e-20, 1.027984e-20, 
    2.055969e-20, -1.027984e-20, 5.653913e-20, -1.541976e-20, 1.027984e-20, 
    -1.027984e-20, 5.139921e-21, 1.541976e-20, -2.006177e-36, -1.541976e-20, 
    -5.139921e-21, -1.541976e-20, 3.597945e-20, -1.541976e-20, -2.055969e-20, 
    -1.027984e-20, 3.597945e-20, -1.027984e-20, -5.139921e-21, 2.569961e-20, 
    -1.027984e-20, -1.027984e-20, 1.027984e-20, 5.139921e-21, 1.027984e-20, 
    -5.139921e-21, 5.139921e-21, 1.027984e-20, 1.027984e-20, 1.541976e-20, 
    3.083953e-20, 5.139921e-21, -2.569961e-20, 2.006177e-36, -5.139921e-21, 
    5.139921e-21, 2.569961e-20, 0, 2.006177e-36, -5.139921e-21, 2.006177e-36, 
    -1.027984e-20, 2.055969e-20, 5.139921e-21, 3.083953e-20, -2.055969e-20, 
    -5.139921e-21, -5.139921e-21, 1.541976e-20, 1.541976e-20, 5.139921e-21, 
    -2.055969e-20, 5.139921e-21, 1.027984e-20, 2.569961e-20, -4.625929e-20, 
    5.139921e-21, 1.027984e-20, 0, -2.055969e-20, -1.027984e-20, 
    -1.027984e-20, -5.139921e-21, -2.055969e-20, -4.625929e-20, 
    -2.006177e-36, 4.111937e-20, -2.055969e-20, -1.027984e-20, 2.569961e-20, 
    -1.027984e-20, 5.139921e-21, 1.027984e-20, 5.139921e-21, -3.083953e-20, 
    2.055969e-20, -2.055969e-20, -1.541976e-20, -5.139921e-21, -1.541976e-20, 
    -4.111937e-20, 3.083953e-20, 1.027984e-20, -3.083953e-20, -4.111937e-20, 
    -5.139921e-21, -5.139921e-21, 2.055969e-20, -2.569961e-20, -1.541976e-20, 
    -5.139921e-21, -5.139921e-21, 4.625929e-20, 1.541976e-20, -3.083953e-20, 
    0, -2.569961e-20, 1.541976e-20, -3.083953e-20, 2.569961e-20, 
    -1.541976e-20, 4.625929e-20, -1.027984e-20, 1.027984e-20, -2.569961e-20, 
    -3.083953e-20, 1.541976e-20, -2.006177e-36, -2.569961e-20, -2.055969e-20, 
    -2.569961e-20, -5.139921e-21, 2.055969e-20, 4.111937e-20, -3.083953e-20, 
    -1.027984e-20, 5.139921e-21, -3.597945e-20, 5.139921e-21, 5.139921e-21, 
    1.027984e-20, 1.027984e-20, -1.027984e-20, 3.083953e-20, -2.055969e-20, 
    -5.139921e-21, 3.597945e-20, 3.083953e-20, -2.055969e-20, 1.027984e-20, 
    5.139921e-21, 5.139921e-21, 1.027984e-20, 2.055969e-20, 1.541976e-20, 
    -5.139921e-21, 2.569961e-20, -5.139921e-21, 2.006177e-36, -5.139921e-21, 
    2.055969e-20, -2.006177e-36, 1.027984e-20, 5.139921e-21, -2.055969e-20, 
    -4.625929e-20, 0, 1.541976e-20, -1.541976e-20, 1.027984e-20, 
    5.139921e-21, -2.055969e-20, -1.541976e-20, -5.139921e-21, 1.541976e-20, 
    -5.139921e-21, -5.139921e-21, 2.569961e-20, -2.006177e-36, 1.541976e-20, 
    5.139921e-21, 5.139921e-21, -1.541976e-20, 2.569961e-20, 0, 1.541976e-20, 
    3.083953e-20, -1.027984e-20, 2.569961e-20, -3.083953e-20, -1.541976e-20, 
    -5.139921e-21, 2.055969e-20, -1.541976e-20, 5.139921e-21, 2.569961e-20, 
    -2.006177e-36, 2.055969e-20, 2.055969e-20, -1.027984e-20, -2.569961e-20, 
    -5.139921e-21, -1.027984e-20, 1.027984e-20, 0, 2.055969e-20, 
    -2.006177e-36, 5.139921e-21, 2.055969e-20, 0, -1.027984e-20, 
    -1.541976e-20, 1.541976e-20, 5.139921e-21, -5.139921e-21, -4.111937e-20, 
    -1.027984e-20, -2.055969e-20, 3.083953e-20, 1.027984e-20, 2.569961e-20, 
    1.027984e-20, -1.027984e-20, -2.006177e-36, -1.027984e-20, -3.083953e-20, 
    1.027984e-20, 3.597945e-20, -1.541976e-20, 0, 5.139921e-21, 
    -1.027984e-20, 0, -2.006177e-36, 2.055969e-20, -2.006177e-36, 
    1.541976e-20, 2.006177e-36, -5.139921e-21, 0, -1.541976e-20, 
    1.541976e-20, -3.597945e-20, 1.027984e-20, 1.027984e-20, 0, 2.055969e-20, 
    -2.569961e-20, 5.139921e-21, -1.541976e-20, -5.139921e-21, 1.027984e-20, 
    2.006177e-36, -2.055969e-20, 2.006177e-36, 1.027984e-20, 1.027984e-20, 
    3.083953e-20, 5.139921e-21, 1.027984e-20, -2.055969e-20, 5.139921e-21, 
    -1.027984e-20, -1.027984e-20, -3.083953e-20, 2.006177e-36, 5.139921e-21, 
    -4.111937e-20, -1.027984e-20, 1.541976e-20, 2.055969e-20, 2.055969e-20, 
    1.027984e-20, -1.541976e-20, 5.139921e-21, 5.139921e-21, -2.055969e-20, 
    1.027984e-20, 2.006177e-36, 3.083953e-20, -2.055969e-20, 1.541976e-20, 
    1.541976e-20, -1.027984e-20, -1.541976e-20, 2.055969e-20, 1.027984e-20, 
    1.027984e-20, -2.569961e-20, -1.541976e-20, 1.027984e-20, -2.569961e-20, 
    1.027984e-20, 1.027984e-20, -2.055969e-20, 2.055969e-20, 2.569961e-20, 
    -1.541976e-20, 5.139921e-21, -5.139921e-21, 0, -1.027984e-20, 
    5.139921e-21, 2.006177e-36, 5.139921e-21, -1.541976e-20, 2.569961e-20, 
    3.083953e-20, 3.597945e-20, -1.027984e-20, -3.597945e-20, 3.597945e-20, 
    -2.006177e-36, -5.139921e-21, -5.139921e-21, -5.139921e-21, 1.027984e-20, 
    1.541976e-20, -2.055969e-20, -2.055969e-20, -5.139921e-21, 3.083953e-20,
  3.083953e-20, 2.055969e-20, 1.027984e-20, -2.055969e-20, 1.027984e-20, 
    2.569961e-20, 0, 1.027984e-20, -5.139921e-21, -2.569961e-20, 
    5.139921e-21, -1.541976e-20, -1.027984e-20, -5.139921e-21, -2.006177e-36, 
    -5.139921e-21, 1.541976e-20, 1.027984e-20, 1.027984e-20, -5.139921e-21, 
    -5.139921e-21, -1.027984e-20, 0, 0, -1.541976e-20, -5.139921e-21, 
    1.027984e-20, 5.139921e-21, 2.006177e-36, -2.055969e-20, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20, -5.139921e-21, -5.139921e-21, 
    5.139921e-21, 1.541976e-20, 2.006177e-36, 1.541976e-20, -3.083953e-20, 
    2.055969e-20, 1.541976e-20, -5.139921e-21, -1.027984e-20, -5.139921e-21, 
    2.055969e-20, 5.139921e-21, 0, -2.569961e-20, 0, -5.139921e-21, 
    2.569961e-20, 1.541976e-20, -1.027984e-20, -5.139921e-21, 0, 
    4.625929e-20, 5.139921e-21, -2.569961e-20, 0, -2.569961e-20, 0, 
    -5.139921e-21, 2.055969e-20, -1.541976e-20, -1.541976e-20, 1.541976e-20, 
    1.541976e-20, 2.055969e-20, -1.541976e-20, -2.569961e-20, 2.055969e-20, 
    2.055969e-20, 2.006177e-36, -5.139921e-21, -1.027984e-20, 1.027984e-20, 
    -2.569961e-20, -1.541976e-20, 5.139921e-21, 5.139921e-21, 2.569961e-20, 
    2.006177e-36, 1.541976e-20, -3.083953e-20, 5.139921e-21, 2.055969e-20, 
    -1.541976e-20, 5.139921e-21, 0, 1.027984e-20, -2.055969e-20, 
    1.027984e-20, -2.006177e-36, 1.027984e-20, -5.139921e-21, 1.027984e-20, 
    -1.027984e-20, 1.027984e-20, -1.541976e-20, -2.055969e-20, -1.027984e-20, 
    3.083953e-20, -4.111937e-20, -1.027984e-20, 1.027984e-20, 2.055969e-20, 
    1.541976e-20, -5.139921e-21, -1.541976e-20, -1.027984e-20, 5.139921e-21, 
    2.569961e-20, -2.569961e-20, 1.027984e-20, -2.006177e-36, 1.541976e-20, 
    1.027984e-20, -2.006177e-36, -1.027984e-20, -1.027984e-20, 5.139921e-21, 
    1.027984e-20, -1.541976e-20, -1.027984e-20, 1.541976e-20, 5.139921e-21, 
    5.139921e-21, 0, 2.055969e-20, 2.569961e-20, 0, 1.027984e-20, 
    -5.139921e-21, -5.139921e-20, 5.139921e-21, 1.541976e-20, -1.027984e-20, 
    -1.541976e-20, -5.139921e-21, -5.139921e-21, -2.055969e-20, 
    -1.027984e-20, 0, -1.027984e-20, -2.006177e-36, 2.055969e-20, 
    -1.027984e-20, -3.083953e-20, 1.541976e-20, -5.139921e-21, -5.139921e-21, 
    2.006177e-36, -1.027984e-20, -5.139921e-21, -3.083953e-20, 5.139921e-21, 
    1.541976e-20, -1.027984e-20, 1.541976e-20, -5.139921e-21, 2.055969e-20, 
    0, -2.006177e-36, 5.139921e-21, -2.006177e-36, 1.027984e-20, 
    2.055969e-20, -1.541976e-20, -2.055969e-20, 5.139921e-21, -5.139921e-21, 
    -1.541976e-20, -5.139921e-21, -2.569961e-20, 1.027984e-20, -1.541976e-20, 
    5.139921e-21, 1.541976e-20, 5.139921e-21, 0, 5.139921e-21, 1.027984e-20, 
    2.569961e-20, -1.541976e-20, 1.027984e-20, 5.139921e-21, -2.055969e-20, 
    5.139921e-21, -3.083953e-20, -5.139921e-21, -1.027984e-20, 1.027984e-20, 
    1.027984e-20, -1.541976e-20, 1.027984e-20, -1.541976e-20, 1.541976e-20, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, -5.139921e-21, 3.083953e-20, 
    5.139921e-21, -5.139921e-21, 1.027984e-20, -1.027984e-20, 1.541976e-20, 
    -5.139921e-21, 1.541976e-20, 0, -1.027984e-20, 0, 1.541976e-20, 
    -2.055969e-20, -1.027984e-20, -2.006177e-36, -1.027984e-20, 
    -1.541976e-20, 2.006177e-36, 1.541976e-20, -2.569961e-20, -5.139921e-21, 
    2.569961e-20, 1.027984e-20, 1.027984e-20, -2.569961e-20, -1.027984e-20, 
    -1.541976e-20, 2.055969e-20, -5.139921e-21, 5.139921e-21, -1.541976e-20, 
    -1.027984e-20, 4.111937e-20, -2.055969e-20, -5.139921e-21, -1.027984e-20, 
    -1.027984e-20, -2.569961e-20, -5.139921e-21, 2.006177e-36, 2.569961e-20, 
    -5.139921e-21, -5.139921e-21, -1.541976e-20, -1.027984e-20, 
    -1.027984e-20, -1.541976e-20, 3.597945e-20, 5.139921e-21, 0, 
    1.541976e-20, -1.027984e-20, -5.139921e-21, 0, 1.027984e-20, 
    5.139921e-21, 0, 1.541976e-20, 5.139921e-21, 2.006177e-36, 4.111937e-20, 
    2.569961e-20, 1.541976e-20, -1.027984e-20, 2.569961e-20, 0, 0, 
    -1.027984e-20, 1.027984e-20, 1.027984e-20, 0, -2.569961e-20, 
    1.027984e-20, 1.541976e-20, -1.027984e-20, 2.055969e-20, 1.027984e-20, 
    -2.569961e-20, -2.055969e-20, 5.139921e-21, -5.139921e-21, -2.569961e-20, 
    1.027984e-20, 1.541976e-20, -1.027984e-20, 1.027984e-20, -1.541976e-20, 
    -1.027984e-20, -5.139921e-21, 0, -1.027984e-20, -2.055969e-20, 
    -2.055969e-20, -1.027984e-20, -2.006177e-36, -5.139921e-21, 
    -3.083953e-20, -1.027984e-20, 3.597945e-20, -1.541976e-20, 1.027984e-20, 
    -2.006177e-36, 5.139921e-21, 2.569961e-20, -2.055969e-20, 2.569961e-20, 
    1.027984e-20, 3.083953e-20, 1.027984e-20, 2.055969e-20, 5.139921e-21, 
    -2.055969e-20, -2.006177e-36, -1.027984e-20, 5.139921e-21, 1.541976e-20, 
    2.569961e-20, 5.139921e-21, 5.139921e-21, -5.139921e-21, 0, 
    -5.139921e-21, 5.139921e-21, -1.541976e-20, -1.541976e-20, -5.139921e-21, 
    1.027984e-20, 2.006177e-36, -1.027984e-20, 1.027984e-20, 1.027984e-20, 
    5.139921e-21, -5.139921e-21, 1.541976e-20, 1.541976e-20,
  -4.111937e-20, 2.055969e-20, 1.027984e-20, -2.055969e-20, 5.139921e-21, 
    -2.055969e-20, 3.597945e-20, 5.139921e-21, -2.569961e-20, 2.006177e-36, 
    1.027984e-20, -1.027984e-20, 0, -1.027984e-20, 0, -3.597945e-20, 
    5.139921e-21, -1.541976e-20, 2.055969e-20, 2.006177e-36, -5.139921e-21, 
    -3.597945e-20, -1.027984e-20, 2.055969e-20, -5.139921e-21, 1.027984e-20, 
    -5.139921e-21, -5.139921e-21, 0, -1.027984e-20, -2.055969e-20, 
    -1.027984e-20, 1.027984e-20, 2.569961e-20, 5.139921e-21, 5.139921e-21, 
    -1.541976e-20, -1.541976e-20, -1.027984e-20, 5.139921e-21, -5.139921e-21, 
    1.027984e-20, 5.139921e-21, -1.027984e-20, -2.055969e-20, 5.139921e-21, 
    1.541976e-20, -2.055969e-20, 5.139921e-21, 0, -5.139921e-21, 
    2.055969e-20, -5.139921e-21, 2.569961e-20, -2.055969e-20, -1.541976e-20, 
    -4.111937e-20, 1.541976e-20, 2.569961e-20, 2.055969e-20, -3.597945e-20, 
    -4.111937e-20, 3.083953e-20, 5.139921e-21, 1.541976e-20, 5.139921e-21, 
    -1.541976e-20, -2.055969e-20, -2.569961e-20, -1.027984e-20, 
    -2.055969e-20, -1.027984e-20, 5.139921e-21, 1.541976e-20, -1.027984e-20, 
    -1.541976e-20, 1.027984e-20, 2.006177e-36, 1.027984e-20, -2.569961e-20, 
    1.541976e-20, 2.055969e-20, 1.541976e-20, -5.139921e-21, -2.055969e-20, 
    -2.006177e-36, -2.055969e-20, 3.083953e-20, 3.083953e-20, -2.055969e-20, 
    0, 1.027984e-20, -1.027984e-20, 0, -5.139921e-21, -2.006177e-36, 
    -1.541976e-20, -2.055969e-20, 2.569961e-20, 2.055969e-20, 2.055969e-20, 
    5.139921e-21, 5.139921e-21, -1.541976e-20, 3.083953e-20, 2.006177e-36, 
    5.139921e-21, -2.006177e-36, -1.027984e-20, 1.541976e-20, 2.055969e-20, 
    0, 1.027984e-20, 1.027984e-20, -5.139921e-21, -2.569961e-20, 
    3.083953e-20, -1.027984e-20, -5.139921e-21, 1.541976e-20, -5.139921e-21, 
    -1.027984e-20, 2.569961e-20, 5.139921e-21, 1.541976e-20, 1.541976e-20, 
    -2.569961e-20, 5.139921e-21, -2.055969e-20, -1.027984e-20, -1.541976e-20, 
    1.027984e-20, -2.006177e-36, 0, 1.541976e-20, -1.541976e-20, 
    2.006177e-36, 1.027984e-20, 5.139921e-21, 1.541976e-20, -2.569961e-20, 
    1.027984e-20, -1.027984e-20, -1.027984e-20, -6.167906e-20, -1.541976e-20, 
    -5.139921e-21, -1.541976e-20, 5.139921e-21, -4.625929e-20, -2.055969e-20, 
    1.541976e-20, 1.027984e-20, 2.055969e-20, 3.083953e-20, 1.027984e-20, 
    -1.027984e-20, -1.027984e-20, -1.027984e-20, 1.027984e-20, -1.027984e-20, 
    -1.541976e-20, -2.006177e-36, 5.139921e-21, 2.006177e-36, -2.006177e-36, 
    0, 2.055969e-20, -1.541976e-20, -5.139921e-21, -1.027984e-20, 
    -2.055969e-20, 2.569961e-20, -5.139921e-21, 0, -1.027984e-20, 
    -2.006177e-36, 5.139921e-21, -5.139921e-21, 1.027984e-20, 2.006177e-36, 
    4.625929e-20, 2.006177e-36, -5.139921e-21, 5.139921e-21, 0, 5.139921e-21, 
    2.055969e-20, -1.027984e-20, -2.569961e-20, 5.139921e-21, 0, 
    -1.541976e-20, 2.055969e-20, 5.139921e-21, 1.027984e-20, 4.111937e-20, 0, 
    -1.541976e-20, 0, -1.541976e-20, -1.027984e-20, 1.027984e-20, 
    1.027984e-20, -2.055969e-20, 1.541976e-20, -1.027984e-20, -1.541976e-20, 
    4.111937e-20, 5.139921e-21, -2.055969e-20, -1.027984e-20, -2.055969e-20, 
    -1.027984e-20, -1.027984e-20, -5.139921e-21, 1.027984e-20, -5.139921e-21, 
    1.027984e-20, 2.055969e-20, 1.541976e-20, 3.083953e-20, 3.597945e-20, 0, 
    -1.027984e-20, 0, -2.006177e-36, -2.055969e-20, -1.027984e-20, 0, 
    1.027984e-20, 1.027984e-20, -2.006177e-36, 1.541976e-20, 2.569961e-20, 
    -5.139921e-21, -1.027984e-20, -5.139921e-21, 1.541976e-20, 5.139921e-21, 
    1.541976e-20, -2.055969e-20, 0, 1.541976e-20, 1.541976e-20, 1.541976e-20, 
    1.541976e-20, -2.055969e-20, -5.139921e-21, -1.541976e-20, -4.111937e-20, 
    2.006177e-36, -5.139921e-21, -5.139921e-21, 2.055969e-20, 1.541976e-20, 
    -2.569961e-20, 5.139921e-21, 2.006177e-36, 0, 0, -1.541976e-20, 
    -1.541976e-20, 1.541976e-20, -2.055969e-20, 2.055969e-20, -2.055969e-20, 
    -2.055969e-20, 1.541976e-20, 4.111937e-20, 1.027984e-20, 2.055969e-20, 
    5.139921e-21, -2.055969e-20, 3.083953e-20, 4.111937e-20, 5.139921e-21, 
    5.139921e-21, 1.541976e-20, 2.006177e-36, -1.027984e-20, 1.027984e-20, 0, 
    -1.541976e-20, -5.139921e-21, -5.139921e-21, 2.055969e-20, 1.541976e-20, 
    -1.027984e-20, -1.027984e-20, 5.139921e-21, 1.541976e-20, -5.139921e-21, 
    -5.139921e-21, -1.541976e-20, 1.541976e-20, -1.541976e-20, -2.569961e-20, 
    -2.006177e-36, 5.139921e-21, -5.139921e-21, 1.541976e-20, -5.139921e-21, 
    2.569961e-20, 2.569961e-20, -2.006177e-36, -1.027984e-20, -1.027984e-20, 
    -5.139921e-21, 1.541976e-20, -2.006177e-36, 2.055969e-20, 3.597945e-20, 
    -4.625929e-20, 5.139921e-21, -1.541976e-20, 5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 1.027984e-20, -5.139921e-21, 3.083953e-20, 1.027984e-20, 
    2.055969e-20, 5.139921e-21, -1.541976e-20, -1.541976e-20, 2.006177e-36, 
    1.027984e-20, -5.139921e-21, -1.541976e-20, 1.541976e-20, 2.055969e-20, 
    1.027984e-20, 1.027984e-20, -1.541976e-20, -5.139921e-21, -5.139921e-21,
  -1.027984e-20, 1.027984e-20, 4.625929e-20, 2.006177e-36, 2.006177e-36, 
    -1.541976e-20, 5.139921e-21, -5.139921e-21, -1.027984e-20, 4.111937e-20, 
    1.027984e-20, 3.083953e-20, 0, -5.139921e-21, -1.541976e-20, 
    4.625929e-20, -5.139921e-21, 3.083953e-20, -2.055969e-20, 0, 
    -1.027984e-20, 3.083953e-20, -2.055969e-20, -5.139921e-21, 1.541976e-20, 
    3.083953e-20, 1.027984e-20, -1.027984e-20, 1.541976e-20, -1.541976e-20, 
    -1.027984e-20, 1.027984e-20, 5.139921e-21, -1.027984e-20, -5.139921e-21, 
    1.027984e-20, 5.139921e-21, -4.111937e-20, -2.055969e-20, -5.139921e-21, 
    1.541976e-20, 5.139921e-20, 2.569961e-20, 1.541976e-20, -1.027984e-20, 
    -1.541976e-20, -1.027984e-20, 5.139921e-21, -1.541976e-20, -1.541976e-20, 
    3.083953e-20, 2.055969e-20, 1.541976e-20, -1.541976e-20, 2.055969e-20, 
    2.055969e-20, 2.055969e-20, 2.055969e-20, 2.055969e-20, -2.055969e-20, 
    -1.541976e-20, -1.027984e-20, -2.055969e-20, 1.027984e-20, 2.055969e-20, 
    0, 4.625929e-20, 1.541976e-20, -1.027984e-20, -1.027984e-20, 
    5.139921e-21, 5.139921e-21, -2.569961e-20, 5.139921e-21, 1.541976e-20, 
    5.139921e-21, 3.597945e-20, -5.139921e-21, 1.541976e-20, -2.006177e-36, 
    4.111937e-20, 3.597945e-20, 1.027984e-20, 5.139921e-21, -1.027984e-20, 
    1.027984e-20, -1.541976e-20, -5.139921e-21, -1.027984e-20, -1.541976e-20, 
    5.139921e-21, 1.027984e-20, 3.597945e-20, -1.027984e-20, -2.055969e-20, 
    0, 2.569961e-20, -2.055969e-20, -1.027984e-20, -1.027984e-20, 
    -4.111937e-20, -5.139921e-21, 0, -1.027984e-20, -2.055969e-20, 
    -2.006177e-36, -3.597945e-20, 0, -5.139921e-21, 0, 1.027984e-20, 
    1.027984e-20, 3.083953e-20, -2.569961e-20, 5.139921e-21, 5.139921e-21, 
    -2.055969e-20, -2.569961e-20, -3.597945e-20, 5.139921e-21, -5.139921e-21, 
    0, 1.541976e-20, 5.139921e-21, 1.541976e-20, 5.139921e-21, 3.083953e-20, 
    3.597945e-20, 1.027984e-20, -5.139921e-21, -1.541976e-20, 5.139921e-21, 
    0, -1.027984e-20, -2.055969e-20, 1.027984e-20, -4.111937e-20, 
    4.625929e-20, -5.139921e-21, -1.027984e-20, 5.139921e-21, 2.569961e-20, 
    5.139921e-21, 0, 3.597945e-20, 1.541976e-20, 5.139921e-21, -1.541976e-20, 
    -1.027984e-20, -1.027984e-20, -5.139921e-21, 2.006177e-36, -1.027984e-20, 
    -1.027984e-20, -1.541976e-20, -2.569961e-20, 5.139921e-21, 1.027984e-20, 
    -5.139921e-21, -1.541976e-20, 1.541976e-20, -1.027984e-20, -2.055969e-20, 
    -1.541976e-20, 1.027984e-20, 5.139921e-21, -2.006177e-36, 3.083953e-20, 
    0, 2.006177e-36, -1.027984e-20, 2.055969e-20, 2.006177e-36, 
    -2.569961e-20, -1.541976e-20, 2.055969e-20, 1.541976e-20, -5.139921e-21, 
    -2.006177e-36, -1.027984e-20, 1.027984e-20, -1.027984e-20, -1.027984e-20, 
    5.139921e-21, 1.541976e-20, 5.139921e-21, -3.083953e-20, 3.597945e-20, 
    2.055969e-20, 2.055969e-20, -1.541976e-20, -2.055969e-20, -1.027984e-20, 
    1.027984e-20, -1.027984e-20, -1.027984e-20, -5.139921e-21, -1.027984e-20, 
    5.139921e-21, -5.139921e-21, 1.027984e-20, -2.055969e-20, -2.006177e-36, 
    1.541976e-20, -1.541976e-20, 0, 1.541976e-20, -1.027984e-20, 
    5.139921e-21, -1.027984e-20, -1.541976e-20, 1.027984e-20, 2.006177e-36, 
    2.055969e-20, 1.027984e-20, 5.139921e-21, 1.541976e-20, -1.541976e-20, 
    1.027984e-20, 1.027984e-20, 2.055969e-20, 2.055969e-20, -1.541976e-20, 
    -1.027984e-20, -2.055969e-20, -5.139921e-21, 1.541976e-20, 1.541976e-20, 
    -4.625929e-20, -1.027984e-20, 0, -2.055969e-20, -3.597945e-20, 
    4.625929e-20, 2.569961e-20, -1.027984e-20, -1.027984e-20, -1.541976e-20, 
    5.139921e-21, 5.139921e-21, 1.541976e-20, 1.027984e-20, 2.569961e-20, 
    -5.139921e-21, -5.139921e-21, -1.541976e-20, 5.139921e-21, -5.139921e-21, 
    -2.055969e-20, 2.569961e-20, -1.027984e-20, -1.541976e-20, -1.541976e-20, 
    -1.541976e-20, 5.139921e-21, -5.139921e-21, 1.027984e-20, -5.139921e-21, 
    2.006177e-36, 4.625929e-20, 1.541976e-20, 2.055969e-20, 5.139921e-21, 
    -1.027984e-20, 2.055969e-20, 0, 1.027984e-20, -4.111937e-20, 
    2.569961e-20, -2.569961e-20, -1.541976e-20, 1.027984e-20, -1.541976e-20, 
    -1.027984e-20, -1.541976e-20, 4.625929e-20, -3.083953e-20, 4.111937e-20, 
    1.541976e-20, -5.139921e-21, 1.541976e-20, -1.541976e-20, 2.055969e-20, 
    1.027984e-20, -2.055969e-20, 3.083953e-20, -1.541976e-20, 1.541976e-20, 
    1.541976e-20, -2.006177e-36, -2.055969e-20, -5.139921e-21, 0, 
    1.027984e-20, -5.139921e-21, 3.083953e-20, 2.006177e-36, 0, 
    -2.055969e-20, 1.027984e-20, -1.027984e-20, -2.569961e-20, -1.027984e-20, 
    5.139921e-21, -1.027984e-20, 3.597945e-20, -5.139921e-21, 2.055969e-20, 
    5.139921e-21, -1.027984e-20, -5.139921e-21, 2.006177e-36, -1.541976e-20, 
    1.541976e-20, 2.055969e-20, 2.569961e-20, -5.139921e-21, 2.055969e-20, 
    1.027984e-20, 3.597945e-20, -1.027984e-20, 1.541976e-20, 5.139921e-21, 
    1.027984e-20, -1.027984e-20, -2.055969e-20, -1.027984e-20, -1.027984e-20, 
    3.083953e-20, 1.541976e-20, -5.139921e-21, 3.597945e-20, 5.139921e-21, 
    -5.139921e-21, 1.027984e-20, 1.541976e-20, -1.027984e-20, -1.541976e-20,
  1.541976e-20, -2.055969e-20, 5.139921e-21, 1.027984e-20, 1.027984e-20, 
    3.083953e-20, 5.139921e-21, -1.541976e-20, -1.541976e-20, 2.055969e-20, 
    1.027984e-20, 2.055969e-20, 5.139921e-21, 2.569961e-20, -1.541976e-20, 
    1.541976e-20, -1.027984e-20, 5.139921e-21, -1.027984e-20, 1.541976e-20, 
    -1.541976e-20, -2.006177e-36, 1.541976e-20, 5.139921e-21, -1.541976e-20, 
    2.055969e-20, 5.139921e-21, 2.569961e-20, 2.569961e-20, -1.541976e-20, 
    -4.111937e-20, 1.027984e-20, -2.569961e-20, -5.139921e-21, -2.006177e-36, 
    -1.541976e-20, -5.139921e-21, 1.027984e-20, -2.569961e-20, 1.027984e-20, 
    2.006177e-36, -2.006177e-36, -2.055969e-20, 0, -2.055969e-20, 
    1.027984e-20, -1.541976e-20, -5.139921e-21, -5.139921e-21, -1.027984e-20, 
    2.055969e-20, 2.055969e-20, 5.139921e-21, 0, -1.541976e-20, 
    -2.006177e-36, 2.569961e-20, -4.111937e-20, 2.055969e-20, -5.139921e-21, 
    -5.139921e-21, -2.055969e-20, 0, 2.006177e-36, 2.055969e-20, 0, 
    3.083953e-20, 2.569961e-20, 2.006177e-36, -1.027984e-20, -1.027984e-20, 
    1.027984e-20, 2.569961e-20, -5.139921e-21, 1.027984e-20, -2.006177e-36, 
    1.027984e-20, 2.055969e-20, 1.541976e-20, 1.027984e-20, -5.139921e-21, 
    -1.541976e-20, 2.569961e-20, -1.541976e-20, 5.139921e-21, 2.055969e-20, 
    5.139921e-21, 0, 1.541976e-20, 1.027984e-20, 1.027984e-20, 1.027984e-20, 
    -5.139921e-21, 1.027984e-20, 2.055969e-20, -1.541976e-20, -1.027984e-20, 
    -1.027984e-20, -1.027984e-20, 2.006177e-36, -5.139921e-21, -2.569961e-20, 
    -1.027984e-20, 2.055969e-20, -1.541976e-20, -2.569961e-20, -1.541976e-20, 
    3.083953e-20, 2.055969e-20, 0, -2.055969e-20, 2.055969e-20, 1.541976e-20, 
    1.541976e-20, -5.139921e-21, -1.541976e-20, 2.006177e-36, -4.625929e-20, 
    0, -5.139921e-21, 5.139921e-21, 2.055969e-20, 1.027984e-20, 0, 
    -1.027984e-20, -1.541976e-20, 2.006177e-36, 5.139921e-21, 5.139921e-21, 
    3.597945e-20, -5.139921e-21, 4.111937e-20, -5.139921e-21, 2.055969e-20, 
    5.139921e-21, 5.139921e-21, 1.541976e-20, 2.006177e-36, -2.055969e-20, 
    2.006177e-36, -1.027984e-20, -1.027984e-20, 2.055969e-20, 0, 
    5.139921e-21, -2.006177e-36, -1.541976e-20, 2.006177e-36, -2.569961e-20, 
    1.541976e-20, -3.083953e-20, 2.569961e-20, 4.625929e-20, -2.055969e-20, 
    2.569961e-20, 2.006177e-36, 1.541976e-20, 0, 2.569961e-20, 1.027984e-20, 
    -1.027984e-20, -2.055969e-20, -1.027984e-20, -2.055969e-20, 
    -2.569961e-20, -2.569961e-20, -5.139921e-21, 1.541976e-20, 0, 
    2.055969e-20, -3.597945e-20, -1.027984e-20, -3.597945e-20, 5.139921e-21, 
    -4.111937e-20, 2.055969e-20, 1.541976e-20, 2.569961e-20, -5.139921e-21, 
    -1.027984e-20, 0, 2.055969e-20, 1.541976e-20, 2.006177e-36, 2.006177e-36, 
    1.541976e-20, 2.055969e-20, -3.083953e-20, -5.139921e-21, -1.027984e-20, 
    1.541976e-20, -1.027984e-20, 4.111937e-20, -5.139921e-21, 3.597945e-20, 
    1.027984e-20, 3.083953e-20, -5.139921e-21, -5.139921e-21, 0, 
    -1.541976e-20, 1.541976e-20, 2.006177e-36, 5.139921e-21, -5.139921e-21, 
    -1.541976e-20, 1.541976e-20, 5.139921e-21, 1.027984e-20, 1.027984e-20, 
    -2.006177e-36, 2.055969e-20, 5.139921e-21, -1.027984e-20, -1.541976e-20, 
    2.569961e-20, 2.006177e-36, 0, 1.541976e-20, -1.541976e-20, 5.139921e-21, 
    1.541976e-20, 2.055969e-20, -1.541976e-20, 2.569961e-20, -2.055969e-20, 
    1.027984e-20, 2.569961e-20, 3.597945e-20, 1.027984e-20, 2.055969e-20, 0, 
    -1.541976e-20, -1.027984e-20, -1.027984e-20, -2.569961e-20, 
    -1.541976e-20, 5.139921e-21, 5.139921e-21, 1.027984e-20, 2.055969e-20, 
    -2.006177e-36, -1.541976e-20, -5.139921e-21, -1.541976e-20, 
    -1.541976e-20, -5.139921e-20, -1.541976e-20, 0, -1.027984e-20, 
    1.027984e-20, 2.569961e-20, 2.569961e-20, 1.027984e-20, 0, -1.027984e-20, 
    -2.569961e-20, 1.541976e-20, -3.083953e-20, 2.569961e-20, 5.139921e-21, 
    5.139921e-21, 2.569961e-20, -1.027984e-20, 1.541976e-20, 1.027984e-20, 
    -5.139921e-21, 1.027984e-20, -3.083953e-20, 2.569961e-20, -2.055969e-20, 
    3.083953e-20, 4.111937e-20, -3.083953e-20, 5.139921e-21, -2.055969e-20, 
    0, -2.006177e-36, 5.139921e-21, 2.006177e-36, 5.139921e-21, 2.006177e-36, 
    5.139921e-21, -1.027984e-20, 2.055969e-20, -5.139921e-21, 0, 
    2.055969e-20, -1.027984e-20, 1.541976e-20, 5.139921e-21, -1.027984e-20, 
    -2.006177e-36, 5.139921e-21, 5.139921e-21, -1.027984e-20, -5.139921e-21, 
    -1.541976e-20, -2.569961e-20, 1.541976e-20, 1.027984e-20, -1.027984e-20, 
    -3.083953e-20, -1.027984e-20, 4.111937e-20, 1.541976e-20, 1.027984e-20, 
    -2.006177e-36, 5.139921e-21, -1.027984e-20, -2.055969e-20, 1.541976e-20, 
    0, -5.139921e-21, 2.055969e-20, 5.139921e-21, -2.006177e-36, 
    3.597945e-20, 2.569961e-20, -5.139921e-21, -2.055969e-20, -5.139921e-21, 
    1.541976e-20, 1.027984e-20, 1.541976e-20, -2.006177e-36, 1.541976e-20, 
    -1.027984e-20, -2.569961e-20, 5.139921e-21, -1.027984e-20, 1.541976e-20, 
    2.055969e-20, 3.083953e-20, -1.027984e-20, -1.027984e-20, 1.541976e-20, 
    -5.139921e-21,
  8.598827e-29, 8.598799e-29, 8.598804e-29, 8.598782e-29, 8.598795e-29, 
    8.598779e-29, 8.598821e-29, 8.598798e-29, 8.598813e-29, 8.598825e-29, 
    8.598738e-29, 8.598781e-29, 8.598694e-29, 8.598721e-29, 8.598652e-29, 
    8.598698e-29, 8.598643e-29, 8.598654e-29, 8.598622e-29, 8.598631e-29, 
    8.59859e-29, 8.598618e-29, 8.59857e-29, 8.598597e-29, 8.598593e-29, 
    8.598619e-29, 8.598772e-29, 8.598743e-29, 8.598774e-29, 8.59877e-29, 
    8.598772e-29, 8.598794e-29, 8.598805e-29, 8.598829e-29, 8.598825e-29, 
    8.598807e-29, 8.598768e-29, 8.598781e-29, 8.598748e-29, 8.598749e-29, 
    8.598711e-29, 8.598728e-29, 8.598665e-29, 8.598683e-29, 8.598631e-29, 
    8.598644e-29, 8.598631e-29, 8.598635e-29, 8.598631e-29, 8.598651e-29, 
    8.598642e-29, 8.598659e-29, 8.598725e-29, 8.598705e-29, 8.598763e-29, 
    8.598798e-29, 8.59882e-29, 8.598837e-29, 8.598834e-29, 8.59883e-29, 
    8.598807e-29, 8.598786e-29, 8.59877e-29, 8.598759e-29, 8.598749e-29, 
    8.598716e-29, 8.598699e-29, 8.598661e-29, 8.598668e-29, 8.598656e-29, 
    8.598645e-29, 8.598627e-29, 8.59863e-29, 8.598621e-29, 8.598657e-29, 
    8.598633e-29, 8.598672e-29, 8.598662e-29, 8.598746e-29, 8.598778e-29, 
    8.598792e-29, 8.598804e-29, 8.598832e-29, 8.598813e-29, 8.59882e-29, 
    8.598802e-29, 8.59879e-29, 8.598796e-29, 8.598759e-29, 8.598773e-29, 
    8.598698e-29, 8.598731e-29, 8.598646e-29, 8.598667e-29, 8.598642e-29, 
    8.598654e-29, 8.598633e-29, 8.598652e-29, 8.598618e-29, 8.598611e-29, 
    8.598616e-29, 8.598597e-29, 8.598653e-29, 8.598631e-29, 8.598796e-29, 
    8.598795e-29, 8.59879e-29, 8.59881e-29, 8.598811e-29, 8.598829e-29, 
    8.598813e-29, 8.598806e-29, 8.598789e-29, 8.598778e-29, 8.598769e-29, 
    8.598747e-29, 8.598723e-29, 8.59869e-29, 8.598665e-29, 8.598649e-29, 
    8.598659e-29, 8.59865e-29, 8.59866e-29, 8.598665e-29, 8.598613e-29, 
    8.598642e-29, 8.598599e-29, 8.598601e-29, 8.598621e-29, 8.598601e-29, 
    8.598794e-29, 8.598799e-29, 8.598819e-29, 8.598804e-29, 8.598831e-29, 
    8.598816e-29, 8.598807e-29, 8.598773e-29, 8.598766e-29, 8.598758e-29, 
    8.598745e-29, 8.598727e-29, 8.598696e-29, 8.598669e-29, 8.598645e-29, 
    8.598646e-29, 8.598646e-29, 8.59864e-29, 8.598654e-29, 8.598638e-29, 
    8.598636e-29, 8.598642e-29, 8.598602e-29, 8.598613e-29, 8.598601e-29, 
    8.598609e-29, 8.598798e-29, 8.598788e-29, 8.598793e-29, 8.598784e-29, 
    8.598791e-29, 8.598761e-29, 8.598752e-29, 8.59871e-29, 8.598727e-29, 
    8.5987e-29, 8.598725e-29, 8.59872e-29, 8.598699e-29, 8.598723e-29, 
    8.598671e-29, 8.598707e-29, 8.59864e-29, 8.598676e-29, 8.598638e-29, 
    8.598645e-29, 8.598633e-29, 8.598623e-29, 8.59861e-29, 8.598586e-29, 
    8.598592e-29, 8.598572e-29, 8.598775e-29, 8.598763e-29, 8.598763e-29, 
    8.598751e-29, 8.598742e-29, 8.598721e-29, 8.598689e-29, 8.598701e-29, 
    8.598678e-29, 8.598674e-29, 8.598708e-29, 8.598687e-29, 8.598754e-29, 
    8.598743e-29, 8.59875e-29, 8.598773e-29, 8.598698e-29, 8.598737e-29, 
    8.598665e-29, 8.598686e-29, 8.598625e-29, 8.598655e-29, 8.598595e-29, 
    8.598569e-29, 8.598545e-29, 8.598516e-29, 8.598756e-29, 8.598764e-29, 
    8.598749e-29, 8.598729e-29, 8.59871e-29, 8.598685e-29, 8.598682e-29, 
    8.598677e-29, 8.598665e-29, 8.598655e-29, 8.598676e-29, 8.598652e-29, 
    8.598741e-29, 8.598695e-29, 8.598767e-29, 8.598745e-29, 8.59873e-29, 
    8.598737e-29, 8.598702e-29, 8.598694e-29, 8.598661e-29, 8.598678e-29, 
    8.598575e-29, 8.598621e-29, 8.598495e-29, 8.59853e-29, 8.598767e-29, 
    8.598756e-29, 8.598717e-29, 8.598736e-29, 8.598683e-29, 8.59867e-29, 
    8.59866e-29, 8.598646e-29, 8.598645e-29, 8.598637e-29, 8.598649e-29, 
    8.598637e-29, 8.598684e-29, 8.598663e-29, 8.598722e-29, 8.598707e-29, 
    8.598714e-29, 8.598721e-29, 8.598699e-29, 8.598675e-29, 8.598675e-29, 
    8.598668e-29, 8.598646e-29, 8.598683e-29, 8.59857e-29, 8.59864e-29, 
    8.598744e-29, 8.598722e-29, 8.598719e-29, 8.598728e-29, 8.598671e-29, 
    8.598692e-29, 8.598637e-29, 8.598652e-29, 8.598627e-29, 8.598639e-29, 
    8.598641e-29, 8.598657e-29, 8.598666e-29, 8.598691e-29, 8.598711e-29, 
    8.598727e-29, 8.598723e-29, 8.598705e-29, 8.598674e-29, 8.598645e-29, 
    8.598651e-29, 8.598629e-29, 8.598687e-29, 8.598663e-29, 8.598672e-29, 
    8.598648e-29, 8.598701e-29, 8.598655e-29, 8.598713e-29, 8.598708e-29, 
    8.598692e-29, 8.598661e-29, 8.598654e-29, 8.598647e-29, 8.598651e-29, 
    8.598674e-29, 8.598677e-29, 8.598693e-29, 8.598697e-29, 8.598708e-29, 
    8.598719e-29, 8.59871e-29, 8.5987e-29, 8.598674e-29, 8.598649e-29, 
    8.598623e-29, 8.598616e-29, 8.598586e-29, 8.598611e-29, 8.598569e-29, 
    8.598604e-29, 8.598544e-29, 8.598653e-29, 8.598606e-29, 8.598692e-29, 
    8.598682e-29, 8.598666e-29, 8.598627e-29, 8.598648e-29, 8.598624e-29, 
    8.598677e-29, 8.598705e-29, 8.598712e-29, 8.598725e-29, 8.598711e-29, 
    8.598713e-29, 8.5987e-29, 8.598704e-29, 8.598672e-29, 8.598689e-29, 
    8.598641e-29, 8.598624e-29, 8.598574e-29, 8.598544e-29, 8.598513e-29, 
    8.598499e-29, 8.598495e-29, 8.598493e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1N_TO_SOIL2N =
  1.134427e-08, 1.139429e-08, 1.138457e-08, 1.142491e-08, 1.140253e-08, 
    1.142895e-08, 1.135441e-08, 1.139627e-08, 1.136955e-08, 1.134878e-08, 
    1.15032e-08, 1.142671e-08, 1.158267e-08, 1.153388e-08, 1.165645e-08, 
    1.157508e-08, 1.167286e-08, 1.165411e-08, 1.171056e-08, 1.169439e-08, 
    1.176659e-08, 1.171802e-08, 1.180403e-08, 1.175499e-08, 1.176266e-08, 
    1.171642e-08, 1.14421e-08, 1.149367e-08, 1.143905e-08, 1.14464e-08, 
    1.14431e-08, 1.140299e-08, 1.138278e-08, 1.134045e-08, 1.134814e-08, 
    1.137922e-08, 1.144971e-08, 1.142578e-08, 1.148609e-08, 1.148473e-08, 
    1.155186e-08, 1.152159e-08, 1.163444e-08, 1.160237e-08, 1.169506e-08, 
    1.167175e-08, 1.169396e-08, 1.168723e-08, 1.169405e-08, 1.165986e-08, 
    1.167451e-08, 1.164443e-08, 1.152726e-08, 1.156169e-08, 1.1459e-08, 
    1.139725e-08, 1.135625e-08, 1.132715e-08, 1.133126e-08, 1.133911e-08, 
    1.137941e-08, 1.14173e-08, 1.144618e-08, 1.14655e-08, 1.148453e-08, 
    1.154214e-08, 1.157264e-08, 1.164093e-08, 1.162861e-08, 1.164948e-08, 
    1.166943e-08, 1.170292e-08, 1.169741e-08, 1.171216e-08, 1.164893e-08, 
    1.169095e-08, 1.162159e-08, 1.164056e-08, 1.148969e-08, 1.143224e-08, 
    1.140781e-08, 1.138643e-08, 1.133443e-08, 1.137034e-08, 1.135618e-08, 
    1.138987e-08, 1.141127e-08, 1.140069e-08, 1.146602e-08, 1.144062e-08, 
    1.157445e-08, 1.15168e-08, 1.16671e-08, 1.163114e-08, 1.167572e-08, 
    1.165297e-08, 1.169196e-08, 1.165687e-08, 1.171765e-08, 1.173088e-08, 
    1.172184e-08, 1.175659e-08, 1.165493e-08, 1.169396e-08, 1.140039e-08, 
    1.140212e-08, 1.141016e-08, 1.13748e-08, 1.137264e-08, 1.134024e-08, 
    1.136907e-08, 1.138135e-08, 1.141251e-08, 1.143095e-08, 1.144847e-08, 
    1.148701e-08, 1.153004e-08, 1.159022e-08, 1.163347e-08, 1.166245e-08, 
    1.164468e-08, 1.166037e-08, 1.164283e-08, 1.163461e-08, 1.172593e-08, 
    1.167465e-08, 1.175159e-08, 1.174733e-08, 1.171251e-08, 1.174781e-08, 
    1.140333e-08, 1.139339e-08, 1.13589e-08, 1.138589e-08, 1.133671e-08, 
    1.136424e-08, 1.138007e-08, 1.144115e-08, 1.145457e-08, 1.146702e-08, 
    1.14916e-08, 1.152314e-08, 1.157848e-08, 1.162663e-08, 1.167059e-08, 
    1.166737e-08, 1.16685e-08, 1.167832e-08, 1.1654e-08, 1.168232e-08, 
    1.168707e-08, 1.167464e-08, 1.174676e-08, 1.172616e-08, 1.174724e-08, 
    1.173383e-08, 1.139662e-08, 1.141334e-08, 1.140431e-08, 1.142129e-08, 
    1.140933e-08, 1.146254e-08, 1.14785e-08, 1.155316e-08, 1.152252e-08, 
    1.157129e-08, 1.152747e-08, 1.153524e-08, 1.157287e-08, 1.152984e-08, 
    1.162397e-08, 1.156015e-08, 1.16787e-08, 1.161496e-08, 1.16827e-08, 
    1.16704e-08, 1.169076e-08, 1.1709e-08, 1.173195e-08, 1.177428e-08, 
    1.176448e-08, 1.179989e-08, 1.143826e-08, 1.145995e-08, 1.145804e-08, 
    1.148073e-08, 1.149752e-08, 1.153389e-08, 1.159224e-08, 1.15703e-08, 
    1.161058e-08, 1.161867e-08, 1.155747e-08, 1.159504e-08, 1.147446e-08, 
    1.149394e-08, 1.148234e-08, 1.143997e-08, 1.157535e-08, 1.150587e-08, 
    1.163418e-08, 1.159654e-08, 1.17064e-08, 1.165176e-08, 1.175908e-08, 
    1.180496e-08, 1.184815e-08, 1.189861e-08, 1.147178e-08, 1.145705e-08, 
    1.148343e-08, 1.151993e-08, 1.15538e-08, 1.159883e-08, 1.160344e-08, 
    1.161188e-08, 1.163373e-08, 1.16521e-08, 1.161454e-08, 1.165671e-08, 
    1.149845e-08, 1.158139e-08, 1.145148e-08, 1.149059e-08, 1.151778e-08, 
    1.150586e-08, 1.156779e-08, 1.158239e-08, 1.164171e-08, 1.161105e-08, 
    1.179364e-08, 1.171285e-08, 1.193705e-08, 1.187439e-08, 1.14519e-08, 
    1.147173e-08, 1.154076e-08, 1.150791e-08, 1.160184e-08, 1.162496e-08, 
    1.164376e-08, 1.166778e-08, 1.167038e-08, 1.168462e-08, 1.166129e-08, 
    1.168369e-08, 1.159893e-08, 1.163681e-08, 1.153287e-08, 1.155816e-08, 
    1.154653e-08, 1.153376e-08, 1.157316e-08, 1.161513e-08, 1.161603e-08, 
    1.162949e-08, 1.166741e-08, 1.160222e-08, 1.180406e-08, 1.16794e-08, 
    1.149336e-08, 1.153156e-08, 1.153702e-08, 1.152222e-08, 1.162264e-08, 
    1.158625e-08, 1.168427e-08, 1.165778e-08, 1.170118e-08, 1.167961e-08, 
    1.167644e-08, 1.164874e-08, 1.163149e-08, 1.158792e-08, 1.155247e-08, 
    1.152436e-08, 1.15309e-08, 1.156178e-08, 1.16177e-08, 1.167061e-08, 
    1.165902e-08, 1.169788e-08, 1.159503e-08, 1.163816e-08, 1.162149e-08, 
    1.166495e-08, 1.156972e-08, 1.165081e-08, 1.154899e-08, 1.155792e-08, 
    1.158553e-08, 1.164108e-08, 1.165337e-08, 1.16665e-08, 1.16584e-08, 
    1.161912e-08, 1.161269e-08, 1.158486e-08, 1.157718e-08, 1.155597e-08, 
    1.153842e-08, 1.155446e-08, 1.15713e-08, 1.161914e-08, 1.166225e-08, 
    1.170926e-08, 1.172077e-08, 1.177568e-08, 1.173097e-08, 1.180475e-08, 
    1.174202e-08, 1.185062e-08, 1.165551e-08, 1.174018e-08, 1.158679e-08, 
    1.160331e-08, 1.16332e-08, 1.170176e-08, 1.166475e-08, 1.170803e-08, 
    1.161244e-08, 1.156284e-08, 1.155001e-08, 1.152607e-08, 1.155056e-08, 
    1.154857e-08, 1.1572e-08, 1.156447e-08, 1.162073e-08, 1.159051e-08, 
    1.167636e-08, 1.170769e-08, 1.179618e-08, 1.185042e-08, 1.190565e-08, 
    1.193003e-08, 1.193745e-08, 1.194056e-08 ;

 SOIL1N_TO_SOIL3N =
  1.346052e-10, 1.351989e-10, 1.350835e-10, 1.355623e-10, 1.352967e-10, 
    1.356103e-10, 1.347256e-10, 1.352224e-10, 1.349053e-10, 1.346587e-10, 
    1.364917e-10, 1.355837e-10, 1.37435e-10, 1.368559e-10, 1.383108e-10, 
    1.373449e-10, 1.385056e-10, 1.38283e-10, 1.389531e-10, 1.387611e-10, 
    1.396183e-10, 1.390417e-10, 1.400627e-10, 1.394806e-10, 1.395716e-10, 
    1.390227e-10, 1.357665e-10, 1.363786e-10, 1.357302e-10, 1.358175e-10, 
    1.357783e-10, 1.353022e-10, 1.350622e-10, 1.345598e-10, 1.346511e-10, 
    1.350201e-10, 1.358567e-10, 1.355727e-10, 1.362885e-10, 1.362724e-10, 
    1.370693e-10, 1.3671e-10, 1.380496e-10, 1.376688e-10, 1.387691e-10, 
    1.384924e-10, 1.387561e-10, 1.386762e-10, 1.387572e-10, 1.383513e-10, 
    1.385252e-10, 1.381681e-10, 1.367773e-10, 1.37186e-10, 1.35967e-10, 
    1.352341e-10, 1.347474e-10, 1.34402e-10, 1.344508e-10, 1.345439e-10, 
    1.350222e-10, 1.35472e-10, 1.358148e-10, 1.360441e-10, 1.362701e-10, 
    1.369539e-10, 1.373159e-10, 1.381266e-10, 1.379803e-10, 1.382281e-10, 
    1.384649e-10, 1.388624e-10, 1.38797e-10, 1.389721e-10, 1.382216e-10, 
    1.387204e-10, 1.37897e-10, 1.381222e-10, 1.363314e-10, 1.356493e-10, 
    1.353594e-10, 1.351057e-10, 1.344883e-10, 1.349146e-10, 1.347466e-10, 
    1.351464e-10, 1.354005e-10, 1.352748e-10, 1.360504e-10, 1.357489e-10, 
    1.373374e-10, 1.366531e-10, 1.384373e-10, 1.380103e-10, 1.385396e-10, 
    1.382695e-10, 1.387323e-10, 1.383158e-10, 1.390373e-10, 1.391944e-10, 
    1.39087e-10, 1.394995e-10, 1.382927e-10, 1.387561e-10, 1.352713e-10, 
    1.352918e-10, 1.353873e-10, 1.349676e-10, 1.349419e-10, 1.345573e-10, 
    1.348995e-10, 1.350453e-10, 1.354152e-10, 1.35634e-10, 1.358421e-10, 
    1.362995e-10, 1.368103e-10, 1.375247e-10, 1.38038e-10, 1.383821e-10, 
    1.381711e-10, 1.383574e-10, 1.381491e-10, 1.380515e-10, 1.391355e-10, 
    1.385268e-10, 1.394402e-10, 1.393896e-10, 1.389763e-10, 1.393953e-10, 
    1.353062e-10, 1.351883e-10, 1.347788e-10, 1.350992e-10, 1.345155e-10, 
    1.348422e-10, 1.350301e-10, 1.357551e-10, 1.359145e-10, 1.360622e-10, 
    1.363539e-10, 1.367284e-10, 1.373852e-10, 1.379568e-10, 1.384787e-10, 
    1.384404e-10, 1.384539e-10, 1.385705e-10, 1.382817e-10, 1.386179e-10, 
    1.386743e-10, 1.385268e-10, 1.393829e-10, 1.391383e-10, 1.393886e-10, 
    1.392293e-10, 1.352266e-10, 1.35425e-10, 1.353178e-10, 1.355194e-10, 
    1.353774e-10, 1.36009e-10, 1.361984e-10, 1.370847e-10, 1.36721e-10, 
    1.372999e-10, 1.367798e-10, 1.368719e-10, 1.373187e-10, 1.368079e-10, 
    1.379253e-10, 1.371677e-10, 1.38575e-10, 1.378184e-10, 1.386224e-10, 
    1.384764e-10, 1.387181e-10, 1.389346e-10, 1.39207e-10, 1.397096e-10, 
    1.395932e-10, 1.400136e-10, 1.357209e-10, 1.359782e-10, 1.359556e-10, 
    1.36225e-10, 1.364242e-10, 1.36856e-10, 1.375486e-10, 1.372882e-10, 
    1.377664e-10, 1.378623e-10, 1.371359e-10, 1.375819e-10, 1.361505e-10, 
    1.363817e-10, 1.362441e-10, 1.357412e-10, 1.373482e-10, 1.365234e-10, 
    1.380465e-10, 1.375996e-10, 1.389038e-10, 1.382552e-10, 1.395292e-10, 
    1.400738e-10, 1.405865e-10, 1.411855e-10, 1.361187e-10, 1.359439e-10, 
    1.36257e-10, 1.366903e-10, 1.370924e-10, 1.376269e-10, 1.376816e-10, 
    1.377817e-10, 1.380411e-10, 1.382592e-10, 1.378134e-10, 1.383139e-10, 
    1.364353e-10, 1.374198e-10, 1.358777e-10, 1.36342e-10, 1.366647e-10, 
    1.365232e-10, 1.372584e-10, 1.374317e-10, 1.381359e-10, 1.377719e-10, 
    1.399393e-10, 1.389803e-10, 1.416418e-10, 1.408979e-10, 1.358827e-10, 
    1.361181e-10, 1.369375e-10, 1.365476e-10, 1.376626e-10, 1.37937e-10, 
    1.381601e-10, 1.384454e-10, 1.384762e-10, 1.386452e-10, 1.383682e-10, 
    1.386342e-10, 1.37628e-10, 1.380777e-10, 1.368438e-10, 1.371441e-10, 
    1.37006e-10, 1.368544e-10, 1.373221e-10, 1.378204e-10, 1.378311e-10, 
    1.379908e-10, 1.38441e-10, 1.376671e-10, 1.400631e-10, 1.385833e-10, 
    1.363749e-10, 1.368283e-10, 1.368931e-10, 1.367174e-10, 1.379095e-10, 
    1.374776e-10, 1.38641e-10, 1.383266e-10, 1.388418e-10, 1.385858e-10, 
    1.385481e-10, 1.382193e-10, 1.380146e-10, 1.374973e-10, 1.370765e-10, 
    1.367429e-10, 1.368205e-10, 1.37187e-10, 1.378509e-10, 1.384789e-10, 
    1.383414e-10, 1.388027e-10, 1.375817e-10, 1.380937e-10, 1.378958e-10, 
    1.384118e-10, 1.372813e-10, 1.382438e-10, 1.370352e-10, 1.371412e-10, 
    1.37469e-10, 1.381284e-10, 1.382743e-10, 1.384301e-10, 1.38334e-10, 
    1.378677e-10, 1.377913e-10, 1.37461e-10, 1.373698e-10, 1.371181e-10, 
    1.369097e-10, 1.371001e-10, 1.373e-10, 1.378679e-10, 1.383797e-10, 
    1.389377e-10, 1.390743e-10, 1.397262e-10, 1.391955e-10, 1.400713e-10, 
    1.393266e-10, 1.406158e-10, 1.382997e-10, 1.393048e-10, 1.374839e-10, 
    1.376801e-10, 1.380348e-10, 1.388486e-10, 1.384093e-10, 1.389231e-10, 
    1.377884e-10, 1.371996e-10, 1.370473e-10, 1.367632e-10, 1.370538e-10, 
    1.370302e-10, 1.373083e-10, 1.37219e-10, 1.378868e-10, 1.375281e-10, 
    1.385472e-10, 1.389191e-10, 1.399695e-10, 1.406135e-10, 1.412691e-10, 
    1.415585e-10, 1.416466e-10, 1.416834e-10 ;

 SOIL1N_vr =
  2.497655, 2.497649, 2.49765, 2.497645, 2.497648, 2.497644, 2.497654, 
    2.497648, 2.497652, 2.497655, 2.497635, 2.497644, 2.497624, 2.497631, 
    2.497615, 2.497625, 2.497613, 2.497615, 2.497608, 2.49761, 2.497601, 
    2.497607, 2.497596, 2.497602, 2.497601, 2.497607, 2.497643, 2.497636, 
    2.497643, 2.497642, 2.497643, 2.497648, 2.49765, 2.497656, 2.497655, 
    2.497651, 2.497642, 2.497645, 2.497637, 2.497637, 2.497628, 2.497632, 
    2.497618, 2.497622, 2.49761, 2.497613, 2.49761, 2.497611, 2.49761, 
    2.497615, 2.497613, 2.497617, 2.497632, 2.497627, 2.49764, 2.497648, 
    2.497653, 2.497657, 2.497657, 2.497656, 2.497651, 2.497646, 2.497642, 
    2.497639, 2.497637, 2.49763, 2.497626, 2.497617, 2.497618, 2.497616, 
    2.497613, 2.497609, 2.49761, 2.497608, 2.497616, 2.497611, 2.497619, 
    2.497617, 2.497636, 2.497644, 2.497647, 2.49765, 2.497656, 2.497652, 
    2.497654, 2.497649, 2.497647, 2.497648, 2.497639, 2.497643, 2.497626, 
    2.497633, 2.497614, 2.497618, 2.497612, 2.497615, 2.49761, 2.497615, 
    2.497607, 2.497605, 2.497607, 2.497602, 2.497615, 2.49761, 2.497648, 
    2.497648, 2.497647, 2.497651, 2.497652, 2.497656, 2.497652, 2.49765, 
    2.497646, 2.497644, 2.497642, 2.497637, 2.497631, 2.497623, 2.497618, 
    2.497614, 2.497617, 2.497614, 2.497617, 2.497618, 2.497606, 2.497613, 
    2.497603, 2.497603, 2.497608, 2.497603, 2.497648, 2.497649, 2.497653, 
    2.49765, 2.497656, 2.497653, 2.497651, 2.497643, 2.497641, 2.497639, 
    2.497636, 2.497632, 2.497625, 2.497619, 2.497613, 2.497613, 2.497613, 
    2.497612, 2.497615, 2.497612, 2.497611, 2.497613, 2.497603, 2.497606, 
    2.497603, 2.497605, 2.497648, 2.497646, 2.497647, 2.497645, 2.497647, 
    2.49764, 2.497638, 2.497628, 2.497632, 2.497626, 2.497632, 2.497631, 
    2.497626, 2.497631, 2.497619, 2.497627, 2.497612, 2.49762, 2.497612, 
    2.497613, 2.497611, 2.497608, 2.497605, 2.4976, 2.497601, 2.497597, 
    2.497643, 2.49764, 2.49764, 2.497638, 2.497635, 2.497631, 2.497623, 
    2.497626, 2.497621, 2.49762, 2.497628, 2.497623, 2.497638, 2.497636, 
    2.497637, 2.497643, 2.497625, 2.497634, 2.497618, 2.497623, 2.497608, 
    2.497616, 2.497602, 2.497596, 2.49759, 2.497584, 2.497639, 2.497641, 
    2.497637, 2.497633, 2.497628, 2.497622, 2.497622, 2.497621, 2.497618, 
    2.497616, 2.49762, 2.497615, 2.497635, 2.497625, 2.497641, 2.497636, 
    2.497633, 2.497634, 2.497626, 2.497624, 2.497617, 2.497621, 2.497597, 
    2.497608, 2.497579, 2.497587, 2.497641, 2.497639, 2.49763, 2.497634, 
    2.497622, 2.497619, 2.497617, 2.497613, 2.497613, 2.497611, 2.497614, 
    2.497612, 2.497622, 2.497617, 2.497631, 2.497627, 2.497629, 2.497631, 
    2.497626, 2.49762, 2.49762, 2.497618, 2.497613, 2.497622, 2.497596, 
    2.497612, 2.497636, 2.497631, 2.49763, 2.497632, 2.497619, 2.497624, 
    2.497611, 2.497615, 2.497609, 2.497612, 2.497612, 2.497616, 2.497618, 
    2.497624, 2.497628, 2.497632, 2.497631, 2.497627, 2.49762, 2.497613, 
    2.497615, 2.49761, 2.497623, 2.497617, 2.497619, 2.497614, 2.497626, 
    2.497616, 2.497629, 2.497627, 2.497624, 2.497617, 2.497615, 2.497614, 
    2.497615, 2.49762, 2.497621, 2.497624, 2.497625, 2.497628, 2.49763, 
    2.497628, 2.497626, 2.49762, 2.497614, 2.497608, 2.497607, 2.4976, 
    2.497605, 2.497596, 2.497604, 2.49759, 2.497615, 2.497604, 2.497624, 
    2.497622, 2.497618, 2.497609, 2.497614, 2.497608, 2.497621, 2.497627, 
    2.497629, 2.497632, 2.497628, 2.497629, 2.497626, 2.497627, 2.49762, 
    2.497623, 2.497612, 2.497608, 2.497597, 2.49759, 2.497583, 2.49758, 
    2.497579, 2.497579,
  2.497912, 2.497904, 2.497906, 2.497899, 2.497903, 2.497899, 2.49791, 
    2.497904, 2.497908, 2.497911, 2.497887, 2.497899, 2.497874, 2.497882, 
    2.497863, 2.497876, 2.49786, 2.497863, 2.497854, 2.497857, 2.497845, 
    2.497853, 2.49784, 2.497847, 2.497846, 2.497853, 2.497897, 2.497889, 
    2.497897, 2.497896, 2.497896, 2.497903, 2.497906, 2.497913, 2.497911, 
    2.497907, 2.497895, 2.497899, 2.49789, 2.49789, 2.497879, 2.497884, 
    2.497866, 2.497871, 2.497857, 2.49786, 2.497857, 2.497858, 2.497857, 
    2.497862, 2.49786, 2.497865, 2.497883, 2.497878, 2.497894, 2.497904, 
    2.49791, 2.497915, 2.497914, 2.497913, 2.497907, 2.4979, 2.497896, 
    2.497893, 2.49789, 2.497881, 2.497876, 2.497865, 2.497867, 2.497864, 
    2.497861, 2.497855, 2.497856, 2.497854, 2.497864, 2.497857, 2.497868, 
    2.497865, 2.497889, 2.497898, 2.497902, 2.497905, 2.497914, 2.497908, 
    2.49791, 2.497905, 2.497901, 2.497903, 2.497893, 2.497897, 2.497876, 
    2.497885, 2.497861, 2.497867, 2.49786, 2.497863, 2.497857, 2.497863, 
    2.497853, 2.497851, 2.497853, 2.497847, 2.497863, 2.497857, 2.497903, 
    2.497903, 2.497902, 2.497907, 2.497908, 2.497913, 2.497908, 2.497906, 
    2.497901, 2.497898, 2.497896, 2.49789, 2.497883, 2.497873, 2.497866, 
    2.497862, 2.497865, 2.497862, 2.497865, 2.497866, 2.497852, 2.49786, 
    2.497848, 2.497849, 2.497854, 2.497849, 2.497903, 2.497904, 2.49791, 
    2.497905, 2.497913, 2.497909, 2.497906, 2.497897, 2.497895, 2.497893, 
    2.497889, 2.497884, 2.497875, 2.497868, 2.497861, 2.497861, 2.497861, 
    2.497859, 2.497863, 2.497859, 2.497858, 2.49786, 2.497849, 2.497852, 
    2.497849, 2.497851, 2.497904, 2.497901, 2.497903, 2.4979, 2.497902, 
    2.497893, 2.497891, 2.497879, 2.497884, 2.497876, 2.497883, 2.497882, 
    2.497876, 2.497883, 2.497868, 2.497878, 2.497859, 2.497869, 2.497859, 
    2.497861, 2.497857, 2.497854, 2.497851, 2.497844, 2.497846, 2.49784, 
    2.497897, 2.497894, 2.497894, 2.49789, 2.497888, 2.497882, 2.497873, 
    2.497876, 2.49787, 2.497869, 2.497878, 2.497873, 2.497892, 2.497889, 
    2.49789, 2.497897, 2.497876, 2.497887, 2.497866, 2.497872, 2.497855, 
    2.497864, 2.497847, 2.497839, 2.497833, 2.497825, 2.497892, 2.497894, 
    2.49789, 2.497884, 2.497879, 2.497872, 2.497871, 2.49787, 2.497866, 
    2.497864, 2.497869, 2.497863, 2.497888, 2.497875, 2.497895, 2.497889, 
    2.497885, 2.497887, 2.497877, 2.497874, 2.497865, 2.49787, 2.497841, 
    2.497854, 2.497819, 2.497828, 2.497895, 2.497892, 2.497881, 2.497886, 
    2.497871, 2.497868, 2.497865, 2.497861, 2.497861, 2.497858, 2.497862, 
    2.497859, 2.497872, 2.497866, 2.497882, 2.497878, 2.49788, 2.497882, 
    2.497876, 2.497869, 2.497869, 2.497867, 2.497861, 2.497871, 2.49784, 
    2.497859, 2.497889, 2.497883, 2.497882, 2.497884, 2.497868, 2.497874, 
    2.497859, 2.497863, 2.497856, 2.497859, 2.49786, 2.497864, 2.497867, 
    2.497874, 2.497879, 2.497884, 2.497883, 2.497878, 2.497869, 2.497861, 
    2.497862, 2.497856, 2.497873, 2.497866, 2.497868, 2.497861, 2.497876, 
    2.497864, 2.49788, 2.497878, 2.497874, 2.497865, 2.497863, 2.497861, 
    2.497863, 2.497869, 2.49787, 2.497874, 2.497875, 2.497879, 2.497881, 
    2.497879, 2.497876, 2.497869, 2.497862, 2.497854, 2.497853, 2.497844, 
    2.497851, 2.497839, 2.497849, 2.497832, 2.497863, 2.49785, 2.497874, 
    2.497871, 2.497866, 2.497856, 2.497862, 2.497855, 2.49787, 2.497878, 
    2.49788, 2.497883, 2.49788, 2.49788, 2.497876, 2.497877, 2.497869, 
    2.497873, 2.49786, 2.497855, 2.497841, 2.497832, 2.497824, 2.49782, 
    2.497819, 2.497818,
  2.498032, 2.498024, 2.498025, 2.498018, 2.498022, 2.498017, 2.49803, 
    2.498023, 2.498028, 2.498031, 2.498004, 2.498018, 2.497991, 2.497999, 
    2.497978, 2.497992, 2.497975, 2.497978, 2.497968, 2.497971, 2.497959, 
    2.497967, 2.497952, 2.497961, 2.497959, 2.497967, 2.498015, 2.498006, 
    2.498016, 2.498014, 2.498015, 2.498022, 2.498025, 2.498033, 2.498031, 
    2.498026, 2.498014, 2.498018, 2.498008, 2.498008, 2.497996, 2.498001, 
    2.497982, 2.497987, 2.497971, 2.497975, 2.497971, 2.497972, 2.497971, 
    2.497977, 2.497975, 2.49798, 2.498, 2.497994, 2.498012, 2.498023, 
    2.49803, 2.498035, 2.498034, 2.498033, 2.498026, 2.498019, 2.498014, 
    2.498011, 2.498008, 2.497998, 2.497992, 2.497981, 2.497983, 2.497979, 
    2.497976, 2.49797, 2.497971, 2.497968, 2.497979, 2.497972, 2.497984, 
    2.497981, 2.498007, 2.498017, 2.498021, 2.498025, 2.498034, 2.498028, 
    2.49803, 2.498024, 2.49802, 2.498022, 2.498011, 2.498015, 2.497992, 
    2.498002, 2.497976, 2.497982, 2.497974, 2.497978, 2.497972, 2.497978, 
    2.497967, 2.497965, 2.497967, 2.49796, 2.497978, 2.497971, 2.498022, 
    2.498022, 2.498021, 2.498027, 2.498027, 2.498033, 2.498028, 2.498026, 
    2.49802, 2.498017, 2.498014, 2.498007, 2.498, 2.497989, 2.497982, 
    2.497977, 2.49798, 2.497977, 2.49798, 2.497982, 2.497966, 2.497975, 
    2.497961, 2.497962, 2.497968, 2.497962, 2.498022, 2.498024, 2.498029, 
    2.498025, 2.498034, 2.498029, 2.498026, 2.498015, 2.498013, 2.498011, 
    2.498006, 2.498001, 2.497991, 2.497983, 2.497975, 2.497976, 2.497976, 
    2.497974, 2.497978, 2.497973, 2.497972, 2.497975, 2.497962, 2.497966, 
    2.497962, 2.497964, 2.498023, 2.49802, 2.498022, 2.498019, 2.498021, 
    2.498012, 2.498009, 2.497996, 2.498001, 2.497993, 2.498, 2.497999, 
    2.497992, 2.498, 2.497983, 2.497994, 2.497974, 2.497985, 2.497973, 
    2.497975, 2.497972, 2.497969, 2.497965, 2.497957, 2.497959, 2.497953, 
    2.498016, 2.498012, 2.498012, 2.498008, 2.498005, 2.497999, 2.497989, 
    2.497993, 2.497986, 2.497984, 2.497995, 2.497988, 2.498009, 2.498006, 
    2.498008, 2.498015, 2.497992, 2.498004, 2.497982, 2.497988, 2.497969, 
    2.497979, 2.49796, 2.497952, 2.497945, 2.497936, 2.49801, 2.498013, 
    2.498008, 2.498002, 2.497996, 2.497988, 2.497987, 2.497986, 2.497982, 
    2.497978, 2.497985, 2.497978, 2.498005, 2.497991, 2.498013, 2.498007, 
    2.498002, 2.498004, 2.497993, 2.497991, 2.49798, 2.497986, 2.497954, 
    2.497968, 2.497929, 2.49794, 2.498013, 2.49801, 2.497998, 2.498004, 
    2.497987, 2.497983, 2.49798, 2.497976, 2.497975, 2.497973, 2.497977, 
    2.497973, 2.497988, 2.497981, 2.497999, 2.497995, 2.497997, 2.497999, 
    2.497992, 2.497985, 2.497985, 2.497983, 2.497976, 2.497987, 2.497952, 
    2.497974, 2.498006, 2.497999, 2.497998, 2.498001, 2.497984, 2.49799, 
    2.497973, 2.497977, 2.49797, 2.497974, 2.497974, 2.497979, 2.497982, 
    2.49799, 2.497996, 2.498001, 2.498, 2.497994, 2.497984, 2.497975, 
    2.497977, 2.497971, 2.497988, 2.497981, 2.497984, 2.497976, 2.497993, 
    2.497979, 2.497997, 2.497995, 2.49799, 2.49798, 2.497978, 2.497976, 
    2.497977, 2.497984, 2.497985, 2.49799, 2.497992, 2.497995, 2.497998, 
    2.497996, 2.497993, 2.497984, 2.497977, 2.497969, 2.497967, 2.497957, 
    2.497965, 2.497952, 2.497963, 2.497944, 2.497978, 2.497963, 2.49799, 
    2.497987, 2.497982, 2.49797, 2.497976, 2.497969, 2.497985, 2.497994, 
    2.497996, 2.498, 2.497996, 2.497997, 2.497993, 2.497994, 2.497984, 
    2.497989, 2.497974, 2.497969, 2.497954, 2.497944, 2.497935, 2.49793, 
    2.497929, 2.497929,
  2.498126, 2.498117, 2.498119, 2.498111, 2.498116, 2.498111, 2.498124, 
    2.498116, 2.498121, 2.498125, 2.498098, 2.498111, 2.498083, 2.498092, 
    2.49807, 2.498085, 2.498067, 2.498071, 2.498061, 2.498064, 2.498051, 
    2.498059, 2.498044, 2.498053, 2.498051, 2.49806, 2.498108, 2.498099, 
    2.498109, 2.498108, 2.498108, 2.498115, 2.498119, 2.498127, 2.498125, 
    2.49812, 2.498107, 2.498111, 2.498101, 2.498101, 2.498089, 2.498094, 
    2.498074, 2.49808, 2.498064, 2.498068, 2.498064, 2.498065, 2.498064, 
    2.49807, 2.498067, 2.498072, 2.498093, 2.498087, 2.498105, 2.498116, 
    2.498124, 2.498129, 2.498128, 2.498127, 2.49812, 2.498113, 2.498108, 
    2.498104, 2.498101, 2.498091, 2.498085, 2.498073, 2.498075, 2.498071, 
    2.498068, 2.498062, 2.498063, 2.49806, 2.498072, 2.498064, 2.498076, 
    2.498073, 2.4981, 2.49811, 2.498115, 2.498118, 2.498127, 2.498121, 
    2.498124, 2.498118, 2.498114, 2.498116, 2.498104, 2.498109, 2.498085, 
    2.498095, 2.498068, 2.498075, 2.498067, 2.498071, 2.498064, 2.49807, 
    2.49806, 2.498057, 2.498059, 2.498053, 2.49807, 2.498064, 2.498116, 
    2.498116, 2.498114, 2.49812, 2.498121, 2.498127, 2.498122, 2.498119, 
    2.498114, 2.49811, 2.498107, 2.498101, 2.498093, 2.498082, 2.498074, 
    2.498069, 2.498072, 2.49807, 2.498073, 2.498074, 2.498058, 2.498067, 
    2.498053, 2.498054, 2.49806, 2.498054, 2.498115, 2.498117, 2.498123, 
    2.498118, 2.498127, 2.498122, 2.498119, 2.498109, 2.498106, 2.498104, 
    2.4981, 2.498094, 2.498084, 2.498075, 2.498068, 2.498068, 2.498068, 
    2.498066, 2.498071, 2.498066, 2.498065, 2.498067, 2.498054, 2.498058, 
    2.498054, 2.498057, 2.498116, 2.498114, 2.498115, 2.498112, 2.498114, 
    2.498105, 2.498102, 2.498089, 2.498094, 2.498085, 2.498093, 2.498092, 
    2.498085, 2.498093, 2.498076, 2.498087, 2.498066, 2.498078, 2.498066, 
    2.498068, 2.498064, 2.498061, 2.498057, 2.498049, 2.498051, 2.498045, 
    2.498109, 2.498105, 2.498106, 2.498101, 2.498099, 2.498092, 2.498082, 
    2.498085, 2.498078, 2.498077, 2.498088, 2.498081, 2.498103, 2.498099, 
    2.498101, 2.498109, 2.498085, 2.498097, 2.498074, 2.498081, 2.498061, 
    2.498071, 2.498052, 2.498044, 2.498036, 2.498027, 2.498103, 2.498106, 
    2.498101, 2.498095, 2.498089, 2.49808, 2.49808, 2.498078, 2.498074, 
    2.498071, 2.498078, 2.49807, 2.498098, 2.498084, 2.498107, 2.4981, 
    2.498095, 2.498097, 2.498086, 2.498083, 2.498073, 2.498078, 2.498046, 
    2.49806, 2.49802, 2.498032, 2.498107, 2.498103, 2.498091, 2.498097, 
    2.49808, 2.498076, 2.498073, 2.498068, 2.498068, 2.498065, 2.49807, 
    2.498065, 2.49808, 2.498074, 2.498092, 2.498088, 2.49809, 2.498092, 
    2.498085, 2.498078, 2.498077, 2.498075, 2.498068, 2.49808, 2.498044, 
    2.498066, 2.498099, 2.498092, 2.498091, 2.498094, 2.498076, 2.498083, 
    2.498065, 2.49807, 2.498062, 2.498066, 2.498067, 2.498072, 2.498075, 
    2.498082, 2.498089, 2.498094, 2.498093, 2.498087, 2.498077, 2.498068, 
    2.49807, 2.498063, 2.498081, 2.498074, 2.498076, 2.498069, 2.498086, 
    2.498071, 2.498089, 2.498088, 2.498083, 2.498073, 2.498071, 2.498069, 
    2.49807, 2.498077, 2.498078, 2.498083, 2.498084, 2.498088, 2.498091, 
    2.498088, 2.498085, 2.498077, 2.498069, 2.498061, 2.498059, 2.498049, 
    2.498057, 2.498044, 2.498055, 2.498036, 2.49807, 2.498055, 2.498083, 
    2.49808, 2.498075, 2.498062, 2.498069, 2.498061, 2.498078, 2.498087, 
    2.498089, 2.498093, 2.498089, 2.49809, 2.498085, 2.498087, 2.498077, 
    2.498082, 2.498067, 2.498061, 2.498045, 2.498036, 2.498026, 2.498022, 
    2.49802, 2.49802,
  2.498261, 2.498253, 2.498254, 2.498248, 2.498251, 2.498247, 2.498259, 
    2.498252, 2.498256, 2.49826, 2.498235, 2.498247, 2.498222, 2.49823, 
    2.49821, 2.498223, 2.498207, 2.49821, 2.498201, 2.498204, 2.498192, 
    2.4982, 2.498186, 2.498194, 2.498193, 2.4982, 2.498245, 2.498236, 
    2.498245, 2.498244, 2.498245, 2.498251, 2.498254, 2.498261, 2.49826, 
    2.498255, 2.498244, 2.498247, 2.498238, 2.498238, 2.498227, 2.498232, 
    2.498214, 2.498219, 2.498204, 2.498208, 2.498204, 2.498205, 2.498204, 
    2.498209, 2.498207, 2.498212, 2.498231, 2.498225, 2.498242, 2.498252, 
    2.498259, 2.498263, 2.498263, 2.498261, 2.498255, 2.498249, 2.498244, 
    2.498241, 2.498238, 2.498229, 2.498224, 2.498213, 2.498214, 2.498211, 
    2.498208, 2.498202, 2.498203, 2.498201, 2.498211, 2.498204, 2.498216, 
    2.498213, 2.498237, 2.498246, 2.49825, 2.498254, 2.498262, 2.498256, 
    2.498259, 2.498253, 2.49825, 2.498251, 2.498241, 2.498245, 2.498223, 
    2.498233, 2.498208, 2.498214, 2.498207, 2.49821, 2.498204, 2.49821, 
    2.4982, 2.498198, 2.498199, 2.498194, 2.49821, 2.498204, 2.498251, 
    2.498251, 2.49825, 2.498256, 2.498256, 2.498261, 2.498257, 2.498255, 
    2.49825, 2.498247, 2.498244, 2.498237, 2.49823, 2.498221, 2.498214, 
    2.498209, 2.498212, 2.498209, 2.498212, 2.498214, 2.498199, 2.498207, 
    2.498194, 2.498195, 2.498201, 2.498195, 2.498251, 2.498253, 2.498258, 
    2.498254, 2.498262, 2.498257, 2.498255, 2.498245, 2.498243, 2.498241, 
    2.498237, 2.498232, 2.498223, 2.498215, 2.498208, 2.498208, 2.498208, 
    2.498206, 2.49821, 2.498206, 2.498205, 2.498207, 2.498195, 2.498199, 
    2.498195, 2.498197, 2.498252, 2.49825, 2.498251, 2.498248, 2.49825, 
    2.498241, 2.498239, 2.498227, 2.498232, 2.498224, 2.498231, 2.49823, 
    2.498224, 2.49823, 2.498215, 2.498226, 2.498206, 2.498217, 2.498206, 
    2.498208, 2.498204, 2.498201, 2.498198, 2.498191, 2.498192, 2.498187, 
    2.498245, 2.498242, 2.498242, 2.498239, 2.498236, 2.49823, 2.49822, 
    2.498224, 2.498217, 2.498216, 2.498226, 2.49822, 2.49824, 2.498236, 
    2.498238, 2.498245, 2.498223, 2.498235, 2.498214, 2.49822, 2.498202, 
    2.498211, 2.498193, 2.498186, 2.498179, 2.49817, 2.49824, 2.498242, 
    2.498238, 2.498232, 2.498227, 2.498219, 2.498219, 2.498217, 2.498214, 
    2.498211, 2.498217, 2.49821, 2.498236, 2.498222, 2.498243, 2.498237, 
    2.498232, 2.498235, 2.498224, 2.498222, 2.498212, 2.498217, 2.498188, 
    2.498201, 2.498164, 2.498174, 2.498243, 2.49824, 2.498229, 2.498234, 
    2.498219, 2.498215, 2.498212, 2.498208, 2.498208, 2.498205, 2.498209, 
    2.498205, 2.498219, 2.498213, 2.49823, 2.498226, 2.498228, 2.49823, 
    2.498224, 2.498217, 2.498217, 2.498214, 2.498208, 2.498219, 2.498186, 
    2.498206, 2.498236, 2.49823, 2.498229, 2.498232, 2.498215, 2.498221, 
    2.498205, 2.49821, 2.498203, 2.498206, 2.498207, 2.498211, 2.498214, 
    2.498221, 2.498227, 2.498231, 2.49823, 2.498225, 2.498216, 2.498208, 
    2.498209, 2.498203, 2.49822, 2.498213, 2.498216, 2.498209, 2.498224, 
    2.498211, 2.498227, 2.498226, 2.498221, 2.498212, 2.49821, 2.498208, 
    2.49821, 2.498216, 2.498217, 2.498222, 2.498223, 2.498226, 2.498229, 
    2.498227, 2.498224, 2.498216, 2.498209, 2.498201, 2.498199, 2.498191, 
    2.498198, 2.498186, 2.498196, 2.498178, 2.49821, 2.498196, 2.498221, 
    2.498219, 2.498214, 2.498203, 2.498209, 2.498202, 2.498217, 2.498225, 
    2.498227, 2.498231, 2.498227, 2.498228, 2.498224, 2.498225, 2.498216, 
    2.498221, 2.498207, 2.498202, 2.498187, 2.498178, 2.498169, 2.498165, 
    2.498164, 2.498164,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL1_HR_S2 =
  5.978543e-08, 6.004907e-08, 5.999782e-08, 6.021046e-08, 6.009251e-08, 
    6.023175e-08, 5.983888e-08, 6.005953e-08, 5.991868e-08, 5.980917e-08, 
    6.062314e-08, 6.021995e-08, 6.104205e-08, 6.078488e-08, 6.143096e-08, 
    6.100203e-08, 6.151746e-08, 6.14186e-08, 6.171618e-08, 6.163093e-08, 
    6.201154e-08, 6.175553e-08, 6.220887e-08, 6.195041e-08, 6.199083e-08, 
    6.174708e-08, 6.03011e-08, 6.057294e-08, 6.0285e-08, 6.032376e-08, 
    6.030637e-08, 6.009494e-08, 5.998839e-08, 5.976528e-08, 5.980579e-08, 
    5.996966e-08, 6.034119e-08, 6.021508e-08, 6.053295e-08, 6.052576e-08, 
    6.087966e-08, 6.072009e-08, 6.131496e-08, 6.114588e-08, 6.163449e-08, 
    6.15116e-08, 6.162871e-08, 6.159321e-08, 6.162917e-08, 6.144895e-08, 
    6.152617e-08, 6.136759e-08, 6.074998e-08, 6.093147e-08, 6.039016e-08, 
    6.006469e-08, 5.984855e-08, 5.969518e-08, 5.971686e-08, 5.975819e-08, 
    5.997062e-08, 6.017036e-08, 6.032258e-08, 6.042441e-08, 6.052473e-08, 
    6.082841e-08, 6.098917e-08, 6.134913e-08, 6.128419e-08, 6.139423e-08, 
    6.149938e-08, 6.16759e-08, 6.164684e-08, 6.172461e-08, 6.139133e-08, 
    6.161283e-08, 6.124719e-08, 6.134719e-08, 6.055196e-08, 6.02491e-08, 
    6.012034e-08, 6.000767e-08, 5.973353e-08, 5.992284e-08, 5.984821e-08, 
    6.002577e-08, 6.013859e-08, 6.008279e-08, 6.042718e-08, 6.029329e-08, 
    6.09987e-08, 6.069484e-08, 6.148711e-08, 6.129752e-08, 6.153256e-08, 
    6.141263e-08, 6.161812e-08, 6.143318e-08, 6.175356e-08, 6.182332e-08, 
    6.177565e-08, 6.19588e-08, 6.142292e-08, 6.16287e-08, 6.008123e-08, 
    6.009033e-08, 6.013273e-08, 5.994635e-08, 5.993495e-08, 5.976418e-08, 
    5.991613e-08, 5.998084e-08, 6.014513e-08, 6.024231e-08, 6.033468e-08, 
    6.053779e-08, 6.076464e-08, 6.108188e-08, 6.130981e-08, 6.14626e-08, 
    6.136892e-08, 6.145162e-08, 6.135916e-08, 6.131582e-08, 6.179718e-08, 
    6.152688e-08, 6.193246e-08, 6.191001e-08, 6.172647e-08, 6.191254e-08, 
    6.009672e-08, 6.004435e-08, 5.986252e-08, 6.000482e-08, 5.974557e-08, 
    5.989068e-08, 5.997411e-08, 6.029608e-08, 6.036683e-08, 6.043243e-08, 
    6.056199e-08, 6.072826e-08, 6.101995e-08, 6.127377e-08, 6.15055e-08, 
    6.148852e-08, 6.14945e-08, 6.154626e-08, 6.141804e-08, 6.156731e-08, 
    6.159236e-08, 6.152685e-08, 6.190701e-08, 6.17984e-08, 6.190954e-08, 
    6.183883e-08, 6.006137e-08, 6.014949e-08, 6.010188e-08, 6.019141e-08, 
    6.012833e-08, 6.040883e-08, 6.049293e-08, 6.088649e-08, 6.072499e-08, 
    6.098205e-08, 6.07511e-08, 6.079202e-08, 6.099041e-08, 6.076358e-08, 
    6.125977e-08, 6.092335e-08, 6.154827e-08, 6.121228e-08, 6.156932e-08, 
    6.150449e-08, 6.161184e-08, 6.170797e-08, 6.182893e-08, 6.20521e-08, 
    6.200042e-08, 6.218706e-08, 6.028086e-08, 6.039516e-08, 6.03851e-08, 
    6.050472e-08, 6.059319e-08, 6.078494e-08, 6.109251e-08, 6.097685e-08, 
    6.118919e-08, 6.123182e-08, 6.090923e-08, 6.110728e-08, 6.047166e-08, 
    6.057434e-08, 6.051321e-08, 6.028988e-08, 6.100349e-08, 6.063724e-08, 
    6.131357e-08, 6.111515e-08, 6.169426e-08, 6.140624e-08, 6.197197e-08, 
    6.221381e-08, 6.244147e-08, 6.270748e-08, 6.045754e-08, 6.037988e-08, 
    6.051895e-08, 6.071134e-08, 6.088989e-08, 6.112725e-08, 6.115155e-08, 
    6.119601e-08, 6.131121e-08, 6.140805e-08, 6.121006e-08, 6.143233e-08, 
    6.059813e-08, 6.103529e-08, 6.035052e-08, 6.055669e-08, 6.070001e-08, 
    6.063715e-08, 6.096364e-08, 6.104058e-08, 6.135328e-08, 6.119164e-08, 
    6.215411e-08, 6.172827e-08, 6.291007e-08, 6.257977e-08, 6.035275e-08, 
    6.045728e-08, 6.082111e-08, 6.0648e-08, 6.11431e-08, 6.126498e-08, 
    6.136406e-08, 6.149071e-08, 6.150439e-08, 6.157943e-08, 6.145646e-08, 
    6.157457e-08, 6.112776e-08, 6.132743e-08, 6.077953e-08, 6.091287e-08, 
    6.085153e-08, 6.078425e-08, 6.099192e-08, 6.121318e-08, 6.121792e-08, 
    6.128886e-08, 6.148876e-08, 6.114511e-08, 6.220905e-08, 6.155194e-08, 
    6.057127e-08, 6.077262e-08, 6.08014e-08, 6.072339e-08, 6.125276e-08, 
    6.106094e-08, 6.15776e-08, 6.143797e-08, 6.166676e-08, 6.155307e-08, 
    6.153633e-08, 6.139032e-08, 6.12994e-08, 6.106973e-08, 6.088288e-08, 
    6.073471e-08, 6.076917e-08, 6.093192e-08, 6.122671e-08, 6.150562e-08, 
    6.144452e-08, 6.164937e-08, 6.11072e-08, 6.133453e-08, 6.124666e-08, 
    6.147578e-08, 6.097378e-08, 6.140122e-08, 6.086452e-08, 6.091157e-08, 
    6.105714e-08, 6.134994e-08, 6.141475e-08, 6.148391e-08, 6.144123e-08, 
    6.12342e-08, 6.120029e-08, 6.10536e-08, 6.101309e-08, 6.090133e-08, 
    6.080879e-08, 6.089333e-08, 6.098212e-08, 6.123429e-08, 6.146155e-08, 
    6.170934e-08, 6.176998e-08, 6.205948e-08, 6.18238e-08, 6.221271e-08, 
    6.188203e-08, 6.245448e-08, 6.142601e-08, 6.187233e-08, 6.106377e-08, 
    6.115087e-08, 6.130841e-08, 6.166979e-08, 6.14747e-08, 6.170286e-08, 
    6.119896e-08, 6.093753e-08, 6.086991e-08, 6.074372e-08, 6.087279e-08, 
    6.086229e-08, 6.09858e-08, 6.094611e-08, 6.124267e-08, 6.108337e-08, 
    6.153591e-08, 6.170107e-08, 6.21675e-08, 6.245345e-08, 6.274457e-08, 
    6.287309e-08, 6.291221e-08, 6.292857e-08 ;

 SOIL1_HR_S3 =
  7.095174e-10, 7.126475e-10, 7.12039e-10, 7.145636e-10, 7.131633e-10, 
    7.148163e-10, 7.101521e-10, 7.127717e-10, 7.110994e-10, 7.097993e-10, 
    7.194632e-10, 7.146763e-10, 7.244367e-10, 7.213833e-10, 7.290542e-10, 
    7.239614e-10, 7.300812e-10, 7.289074e-10, 7.324406e-10, 7.314284e-10, 
    7.359474e-10, 7.329078e-10, 7.382904e-10, 7.352216e-10, 7.357016e-10, 
    7.328075e-10, 7.156398e-10, 7.188671e-10, 7.154485e-10, 7.159087e-10, 
    7.157022e-10, 7.131921e-10, 7.119271e-10, 7.092784e-10, 7.097593e-10, 
    7.117047e-10, 7.161157e-10, 7.146184e-10, 7.183922e-10, 7.18307e-10, 
    7.225087e-10, 7.206142e-10, 7.276769e-10, 7.256695e-10, 7.314706e-10, 
    7.300116e-10, 7.314021e-10, 7.309805e-10, 7.314075e-10, 7.292678e-10, 
    7.301845e-10, 7.283018e-10, 7.20969e-10, 7.231238e-10, 7.166971e-10, 
    7.12833e-10, 7.10267e-10, 7.08446e-10, 7.087035e-10, 7.091941e-10, 
    7.117161e-10, 7.140875e-10, 7.158947e-10, 7.171036e-10, 7.182948e-10, 
    7.219002e-10, 7.238089e-10, 7.280827e-10, 7.273115e-10, 7.286181e-10, 
    7.298665e-10, 7.319623e-10, 7.316174e-10, 7.325408e-10, 7.285837e-10, 
    7.312135e-10, 7.268722e-10, 7.280596e-10, 7.186181e-10, 7.150224e-10, 
    7.134936e-10, 7.12156e-10, 7.089014e-10, 7.111489e-10, 7.102628e-10, 
    7.123709e-10, 7.137103e-10, 7.130479e-10, 7.171366e-10, 7.15547e-10, 
    7.23922e-10, 7.203144e-10, 7.297208e-10, 7.274698e-10, 7.302605e-10, 
    7.288365e-10, 7.312764e-10, 7.290805e-10, 7.328845e-10, 7.337128e-10, 
    7.331467e-10, 7.353212e-10, 7.289587e-10, 7.31402e-10, 7.130293e-10, 
    7.131373e-10, 7.136407e-10, 7.11428e-10, 7.112926e-10, 7.092651e-10, 
    7.110693e-10, 7.118375e-10, 7.13788e-10, 7.149417e-10, 7.160384e-10, 
    7.184499e-10, 7.211431e-10, 7.249095e-10, 7.276157e-10, 7.294298e-10, 
    7.283175e-10, 7.292995e-10, 7.282017e-10, 7.276872e-10, 7.334023e-10, 
    7.301931e-10, 7.350085e-10, 7.34742e-10, 7.325627e-10, 7.347721e-10, 
    7.132132e-10, 7.125915e-10, 7.104328e-10, 7.121221e-10, 7.090444e-10, 
    7.107671e-10, 7.117576e-10, 7.155801e-10, 7.164201e-10, 7.171989e-10, 
    7.187371e-10, 7.207112e-10, 7.241743e-10, 7.271879e-10, 7.299391e-10, 
    7.297375e-10, 7.298085e-10, 7.304231e-10, 7.289007e-10, 7.30673e-10, 
    7.309705e-10, 7.301927e-10, 7.347064e-10, 7.334168e-10, 7.347364e-10, 
    7.338968e-10, 7.127936e-10, 7.138397e-10, 7.132744e-10, 7.143374e-10, 
    7.135885e-10, 7.169187e-10, 7.179172e-10, 7.225898e-10, 7.206722e-10, 
    7.237243e-10, 7.209823e-10, 7.214681e-10, 7.238236e-10, 7.211305e-10, 
    7.270216e-10, 7.230274e-10, 7.30447e-10, 7.264578e-10, 7.306969e-10, 
    7.299272e-10, 7.312017e-10, 7.323431e-10, 7.337792e-10, 7.36429e-10, 
    7.358154e-10, 7.380315e-10, 7.153995e-10, 7.167564e-10, 7.16637e-10, 
    7.180572e-10, 7.191075e-10, 7.213841e-10, 7.250358e-10, 7.236626e-10, 
    7.261836e-10, 7.266897e-10, 7.228597e-10, 7.252111e-10, 7.176646e-10, 
    7.188837e-10, 7.181579e-10, 7.155064e-10, 7.239789e-10, 7.196305e-10, 
    7.276604e-10, 7.253046e-10, 7.321804e-10, 7.287607e-10, 7.354776e-10, 
    7.38349e-10, 7.410522e-10, 7.442107e-10, 7.174971e-10, 7.16575e-10, 
    7.182261e-10, 7.205103e-10, 7.226301e-10, 7.254483e-10, 7.257367e-10, 
    7.262646e-10, 7.276323e-10, 7.287822e-10, 7.264315e-10, 7.290705e-10, 
    7.191662e-10, 7.243564e-10, 7.162264e-10, 7.186742e-10, 7.203757e-10, 
    7.196294e-10, 7.235057e-10, 7.244192e-10, 7.281319e-10, 7.262128e-10, 
    7.376402e-10, 7.32584e-10, 7.466162e-10, 7.426943e-10, 7.162529e-10, 
    7.17494e-10, 7.218135e-10, 7.197583e-10, 7.256364e-10, 7.270834e-10, 
    7.282598e-10, 7.297635e-10, 7.29926e-10, 7.308169e-10, 7.293569e-10, 
    7.307593e-10, 7.254543e-10, 7.278249e-10, 7.213199e-10, 7.22903e-10, 
    7.221748e-10, 7.213758e-10, 7.238415e-10, 7.264684e-10, 7.265247e-10, 
    7.273671e-10, 7.297404e-10, 7.256603e-10, 7.382925e-10, 7.304906e-10, 
    7.188473e-10, 7.212378e-10, 7.215795e-10, 7.206534e-10, 7.269383e-10, 
    7.24661e-10, 7.307952e-10, 7.291373e-10, 7.318538e-10, 7.305039e-10, 
    7.303053e-10, 7.285716e-10, 7.274922e-10, 7.247654e-10, 7.225468e-10, 
    7.207878e-10, 7.211968e-10, 7.231291e-10, 7.266291e-10, 7.299406e-10, 
    7.292152e-10, 7.316474e-10, 7.252102e-10, 7.279092e-10, 7.26866e-10, 
    7.295863e-10, 7.236261e-10, 7.28701e-10, 7.223289e-10, 7.228876e-10, 
    7.246158e-10, 7.280922e-10, 7.288616e-10, 7.296829e-10, 7.291761e-10, 
    7.267181e-10, 7.263154e-10, 7.245738e-10, 7.240929e-10, 7.22766e-10, 
    7.216673e-10, 7.22671e-10, 7.237251e-10, 7.267191e-10, 7.294174e-10, 
    7.323593e-10, 7.330794e-10, 7.365167e-10, 7.337184e-10, 7.383359e-10, 
    7.344098e-10, 7.412067e-10, 7.289954e-10, 7.342946e-10, 7.246945e-10, 
    7.257287e-10, 7.275991e-10, 7.318898e-10, 7.295735e-10, 7.322825e-10, 
    7.262996e-10, 7.231957e-10, 7.223929e-10, 7.208947e-10, 7.224271e-10, 
    7.223025e-10, 7.237689e-10, 7.232977e-10, 7.268185e-10, 7.249273e-10, 
    7.303003e-10, 7.322611e-10, 7.377992e-10, 7.411944e-10, 7.446511e-10, 
    7.461771e-10, 7.466416e-10, 7.468358e-10 ;

 SOIL2C =
  5.783956, 5.783962, 5.78396, 5.783966, 5.783963, 5.783966, 5.783957, 
    5.783962, 5.783959, 5.783956, 5.783975, 5.783966, 5.783984, 5.783978, 
    5.783993, 5.783983, 5.783995, 5.783993, 5.784, 5.783998, 5.784007, 
    5.784001, 5.784011, 5.784005, 5.784006, 5.784, 5.783967, 5.783974, 
    5.783967, 5.783968, 5.783967, 5.783963, 5.78396, 5.783955, 5.783956, 
    5.78396, 5.783968, 5.783966, 5.783973, 5.783973, 5.783981, 5.783977, 
    5.78399, 5.783987, 5.783998, 5.783995, 5.783998, 5.783997, 5.783998, 
    5.783994, 5.783996, 5.783992, 5.783978, 5.783982, 5.783969, 5.783962, 
    5.783957, 5.783954, 5.783954, 5.783955, 5.78396, 5.783965, 5.783968, 
    5.78397, 5.783973, 5.783979, 5.783983, 5.783991, 5.78399, 5.783992, 
    5.783995, 5.783999, 5.783998, 5.784, 5.783992, 5.783998, 5.783989, 
    5.783991, 5.783973, 5.783966, 5.783963, 5.783961, 5.783955, 5.783959, 
    5.783957, 5.783961, 5.783964, 5.783963, 5.78397, 5.783967, 5.783983, 
    5.783977, 5.783995, 5.78399, 5.783996, 5.783993, 5.783998, 5.783993, 
    5.784, 5.784002, 5.784001, 5.784005, 5.783993, 5.783998, 5.783962, 
    5.783963, 5.783964, 5.783959, 5.783959, 5.783955, 5.783959, 5.78396, 
    5.783964, 5.783966, 5.783968, 5.783973, 5.783978, 5.783985, 5.78399, 
    5.783994, 5.783992, 5.783994, 5.783992, 5.78399, 5.784001, 5.783996, 
    5.784005, 5.784004, 5.784, 5.784004, 5.783963, 5.783962, 5.783957, 
    5.783961, 5.783955, 5.783958, 5.78396, 5.783967, 5.783969, 5.78397, 
    5.783973, 5.783977, 5.783984, 5.783989, 5.783995, 5.783995, 5.783995, 
    5.783996, 5.783993, 5.783997, 5.783997, 5.783996, 5.784004, 5.784002, 
    5.784004, 5.784002, 5.783962, 5.783964, 5.783963, 5.783965, 5.783964, 
    5.78397, 5.783972, 5.783981, 5.783977, 5.783983, 5.783978, 5.783978, 
    5.783983, 5.783978, 5.783989, 5.783982, 5.783996, 5.783988, 5.783997, 
    5.783995, 5.783998, 5.783999, 5.784002, 5.784008, 5.784006, 5.78401, 
    5.783967, 5.783969, 5.783969, 5.783972, 5.783974, 5.783978, 5.783986, 
    5.783983, 5.783988, 5.783988, 5.783981, 5.783986, 5.783971, 5.783974, 
    5.783972, 5.783967, 5.783984, 5.783975, 5.78399, 5.783986, 5.783999, 
    5.783993, 5.784006, 5.784011, 5.784016, 5.784022, 5.783971, 5.783969, 
    5.783972, 5.783977, 5.783981, 5.783986, 5.783987, 5.783988, 5.78399, 
    5.783993, 5.783988, 5.783993, 5.783974, 5.783984, 5.783968, 5.783973, 
    5.783977, 5.783975, 5.783983, 5.783984, 5.783991, 5.783988, 5.78401, 
    5.784, 5.784027, 5.784019, 5.783968, 5.783971, 5.783979, 5.783976, 
    5.783987, 5.783989, 5.783992, 5.783995, 5.783995, 5.783997, 5.783994, 
    5.783997, 5.783986, 5.783991, 5.783978, 5.783981, 5.78398, 5.783978, 
    5.783983, 5.783988, 5.783988, 5.78399, 5.783995, 5.783987, 5.784011, 
    5.783996, 5.783974, 5.783978, 5.783979, 5.783977, 5.783989, 5.783985, 
    5.783997, 5.783993, 5.783998, 5.783996, 5.783996, 5.783992, 5.78399, 
    5.783985, 5.783981, 5.783978, 5.783978, 5.783982, 5.783988, 5.783995, 
    5.783994, 5.783998, 5.783986, 5.783991, 5.783989, 5.783994, 5.783983, 
    5.783993, 5.78398, 5.783981, 5.783985, 5.783991, 5.783993, 5.783995, 
    5.783993, 5.783989, 5.783988, 5.783985, 5.783984, 5.783981, 5.783979, 
    5.783981, 5.783983, 5.783989, 5.783994, 5.783999, 5.784001, 5.784008, 
    5.784002, 5.784011, 5.784004, 5.784017, 5.783993, 5.784003, 5.783985, 
    5.783987, 5.78399, 5.783998, 5.783994, 5.783999, 5.783988, 5.783982, 
    5.78398, 5.783978, 5.78398, 5.78398, 5.783983, 5.783982, 5.783989, 
    5.783985, 5.783996, 5.783999, 5.78401, 5.784017, 5.784023, 5.784026, 
    5.784027, 5.784028 ;

 SOIL2C_TO_SOIL1C =
  1.057659e-09, 1.062326e-09, 1.061419e-09, 1.065184e-09, 1.063096e-09, 
    1.065561e-09, 1.058605e-09, 1.062512e-09, 1.060018e-09, 1.058079e-09, 
    1.07249e-09, 1.065352e-09, 1.079906e-09, 1.075353e-09, 1.086791e-09, 
    1.079198e-09, 1.088323e-09, 1.086573e-09, 1.091841e-09, 1.090332e-09, 
    1.09707e-09, 1.092538e-09, 1.100564e-09, 1.095988e-09, 1.096703e-09, 
    1.092388e-09, 1.066788e-09, 1.071601e-09, 1.066503e-09, 1.06719e-09, 
    1.066882e-09, 1.063139e-09, 1.061252e-09, 1.057302e-09, 1.05802e-09, 
    1.060921e-09, 1.067498e-09, 1.065265e-09, 1.070893e-09, 1.070766e-09, 
    1.077031e-09, 1.074206e-09, 1.084738e-09, 1.081744e-09, 1.090395e-09, 
    1.088219e-09, 1.090292e-09, 1.089664e-09, 1.090301e-09, 1.08711e-09, 
    1.088477e-09, 1.085669e-09, 1.074735e-09, 1.077948e-09, 1.068365e-09, 
    1.062603e-09, 1.058777e-09, 1.056061e-09, 1.056445e-09, 1.057177e-09, 
    1.060938e-09, 1.064474e-09, 1.067169e-09, 1.068971e-09, 1.070748e-09, 
    1.076124e-09, 1.07897e-09, 1.085343e-09, 1.084193e-09, 1.086141e-09, 
    1.088003e-09, 1.091128e-09, 1.090613e-09, 1.09199e-09, 1.08609e-09, 
    1.090011e-09, 1.083538e-09, 1.085308e-09, 1.07123e-09, 1.065868e-09, 
    1.063588e-09, 1.061593e-09, 1.05674e-09, 1.060092e-09, 1.058771e-09, 
    1.061914e-09, 1.063911e-09, 1.062924e-09, 1.069021e-09, 1.06665e-09, 
    1.079139e-09, 1.073759e-09, 1.087786e-09, 1.084429e-09, 1.08859e-09, 
    1.086467e-09, 1.090105e-09, 1.086831e-09, 1.092503e-09, 1.093738e-09, 
    1.092894e-09, 1.096136e-09, 1.086649e-09, 1.090292e-09, 1.062896e-09, 
    1.063057e-09, 1.063807e-09, 1.060508e-09, 1.060306e-09, 1.057283e-09, 
    1.059973e-09, 1.061119e-09, 1.064027e-09, 1.065747e-09, 1.067383e-09, 
    1.070979e-09, 1.074995e-09, 1.080611e-09, 1.084646e-09, 1.087352e-09, 
    1.085693e-09, 1.087157e-09, 1.08552e-09, 1.084753e-09, 1.093275e-09, 
    1.08849e-09, 1.09567e-09, 1.095273e-09, 1.092023e-09, 1.095317e-09, 
    1.06317e-09, 1.062243e-09, 1.059024e-09, 1.061543e-09, 1.056954e-09, 
    1.059522e-09, 1.061e-09, 1.0667e-09, 1.067952e-09, 1.069113e-09, 
    1.071407e-09, 1.074351e-09, 1.079515e-09, 1.084009e-09, 1.088111e-09, 
    1.08781e-09, 1.087916e-09, 1.088833e-09, 1.086563e-09, 1.089205e-09, 
    1.089649e-09, 1.088489e-09, 1.095219e-09, 1.093297e-09, 1.095264e-09, 
    1.094012e-09, 1.062544e-09, 1.064104e-09, 1.063261e-09, 1.064847e-09, 
    1.06373e-09, 1.068696e-09, 1.070185e-09, 1.077152e-09, 1.074293e-09, 
    1.078844e-09, 1.074755e-09, 1.07548e-09, 1.078992e-09, 1.074976e-09, 
    1.083761e-09, 1.077805e-09, 1.088868e-09, 1.08292e-09, 1.089241e-09, 
    1.088093e-09, 1.089994e-09, 1.091696e-09, 1.093837e-09, 1.097788e-09, 
    1.096873e-09, 1.100178e-09, 1.06643e-09, 1.068454e-09, 1.068276e-09, 
    1.070393e-09, 1.07196e-09, 1.075354e-09, 1.080799e-09, 1.078752e-09, 
    1.082511e-09, 1.083266e-09, 1.077555e-09, 1.081061e-09, 1.069808e-09, 
    1.071626e-09, 1.070544e-09, 1.06659e-09, 1.079223e-09, 1.072739e-09, 
    1.084713e-09, 1.0812e-09, 1.091453e-09, 1.086354e-09, 1.096369e-09, 
    1.100651e-09, 1.104682e-09, 1.109391e-09, 1.069558e-09, 1.068183e-09, 
    1.070645e-09, 1.074051e-09, 1.077212e-09, 1.081415e-09, 1.081845e-09, 
    1.082632e-09, 1.084671e-09, 1.086386e-09, 1.082881e-09, 1.086816e-09, 
    1.072047e-09, 1.079786e-09, 1.067663e-09, 1.071313e-09, 1.073851e-09, 
    1.072738e-09, 1.078518e-09, 1.07988e-09, 1.085416e-09, 1.082554e-09, 
    1.099594e-09, 1.092055e-09, 1.112978e-09, 1.10713e-09, 1.067703e-09, 
    1.069553e-09, 1.075995e-09, 1.07293e-09, 1.081695e-09, 1.083853e-09, 
    1.085607e-09, 1.087849e-09, 1.088091e-09, 1.08942e-09, 1.087243e-09, 
    1.089334e-09, 1.081424e-09, 1.084958e-09, 1.075259e-09, 1.077619e-09, 
    1.076533e-09, 1.075342e-09, 1.079019e-09, 1.082936e-09, 1.08302e-09, 
    1.084276e-09, 1.087815e-09, 1.081731e-09, 1.100567e-09, 1.088933e-09, 
    1.071572e-09, 1.075136e-09, 1.075646e-09, 1.074265e-09, 1.083637e-09, 
    1.080241e-09, 1.089387e-09, 1.086915e-09, 1.090966e-09, 1.088953e-09, 
    1.088657e-09, 1.086072e-09, 1.084462e-09, 1.080396e-09, 1.077088e-09, 
    1.074465e-09, 1.075075e-09, 1.077956e-09, 1.083175e-09, 1.088113e-09, 
    1.087031e-09, 1.090658e-09, 1.08106e-09, 1.085084e-09, 1.083529e-09, 
    1.087585e-09, 1.078697e-09, 1.086265e-09, 1.076763e-09, 1.077596e-09, 
    1.080173e-09, 1.085357e-09, 1.086504e-09, 1.087729e-09, 1.086973e-09, 
    1.083308e-09, 1.082708e-09, 1.080111e-09, 1.079393e-09, 1.077415e-09, 
    1.075777e-09, 1.077273e-09, 1.078845e-09, 1.08331e-09, 1.087333e-09, 
    1.09172e-09, 1.092794e-09, 1.097919e-09, 1.093746e-09, 1.100631e-09, 
    1.094777e-09, 1.104912e-09, 1.086704e-09, 1.094605e-09, 1.080291e-09, 
    1.081833e-09, 1.084622e-09, 1.09102e-09, 1.087566e-09, 1.091605e-09, 
    1.082684e-09, 1.078056e-09, 1.076858e-09, 1.074625e-09, 1.07691e-09, 
    1.076724e-09, 1.07891e-09, 1.078208e-09, 1.083458e-09, 1.080638e-09, 
    1.08865e-09, 1.091573e-09, 1.099831e-09, 1.104894e-09, 1.110048e-09, 
    1.112323e-09, 1.113016e-09, 1.113305e-09 ;

 SOIL2C_TO_SOIL3C =
  7.554707e-11, 7.588046e-11, 7.581565e-11, 7.608456e-11, 7.59354e-11, 
    7.611147e-11, 7.561467e-11, 7.589369e-11, 7.571557e-11, 7.557709e-11, 
    7.660642e-11, 7.609656e-11, 7.713615e-11, 7.681093e-11, 7.762796e-11, 
    7.708553e-11, 7.773734e-11, 7.761233e-11, 7.798864e-11, 7.788083e-11, 
    7.836214e-11, 7.80384e-11, 7.861169e-11, 7.828484e-11, 7.833596e-11, 
    7.802772e-11, 7.619918e-11, 7.654293e-11, 7.617881e-11, 7.622782e-11, 
    7.620583e-11, 7.593847e-11, 7.580372e-11, 7.55216e-11, 7.557283e-11, 
    7.578004e-11, 7.624987e-11, 7.609039e-11, 7.649235e-11, 7.648328e-11, 
    7.69308e-11, 7.672901e-11, 7.748126e-11, 7.726746e-11, 7.788533e-11, 
    7.772993e-11, 7.787803e-11, 7.783313e-11, 7.787861e-11, 7.765071e-11, 
    7.774835e-11, 7.754782e-11, 7.67668e-11, 7.699632e-11, 7.63118e-11, 
    7.590022e-11, 7.56269e-11, 7.543295e-11, 7.546037e-11, 7.551264e-11, 
    7.578126e-11, 7.603384e-11, 7.622633e-11, 7.63551e-11, 7.648197e-11, 
    7.686598e-11, 7.706928e-11, 7.752449e-11, 7.744235e-11, 7.758151e-11, 
    7.771447e-11, 7.79377e-11, 7.790096e-11, 7.799931e-11, 7.757785e-11, 
    7.785794e-11, 7.739556e-11, 7.752202e-11, 7.65164e-11, 7.613342e-11, 
    7.597058e-11, 7.582811e-11, 7.548145e-11, 7.572084e-11, 7.562647e-11, 
    7.5851e-11, 7.599367e-11, 7.592311e-11, 7.635861e-11, 7.61893e-11, 
    7.708133e-11, 7.669709e-11, 7.769897e-11, 7.745921e-11, 7.775643e-11, 
    7.760477e-11, 7.786464e-11, 7.763076e-11, 7.803591e-11, 7.812413e-11, 
    7.806385e-11, 7.829545e-11, 7.761779e-11, 7.787802e-11, 7.592113e-11, 
    7.593264e-11, 7.598625e-11, 7.575057e-11, 7.573615e-11, 7.552019e-11, 
    7.571236e-11, 7.579419e-11, 7.600194e-11, 7.612482e-11, 7.624164e-11, 
    7.649849e-11, 7.678535e-11, 7.718651e-11, 7.747475e-11, 7.766796e-11, 
    7.754949e-11, 7.765408e-11, 7.753716e-11, 7.748236e-11, 7.809108e-11, 
    7.774926e-11, 7.826214e-11, 7.823376e-11, 7.800165e-11, 7.823696e-11, 
    7.594072e-11, 7.587449e-11, 7.564457e-11, 7.582451e-11, 7.549668e-11, 
    7.568017e-11, 7.578568e-11, 7.619282e-11, 7.628229e-11, 7.636524e-11, 
    7.652908e-11, 7.673934e-11, 7.710821e-11, 7.742918e-11, 7.772221e-11, 
    7.770074e-11, 7.770831e-11, 7.777376e-11, 7.761161e-11, 7.780038e-11, 
    7.783205e-11, 7.774922e-11, 7.822996e-11, 7.809262e-11, 7.823316e-11, 
    7.814373e-11, 7.589603e-11, 7.600745e-11, 7.594724e-11, 7.606046e-11, 
    7.598069e-11, 7.63354e-11, 7.644176e-11, 7.693944e-11, 7.67352e-11, 
    7.706027e-11, 7.676822e-11, 7.681997e-11, 7.707085e-11, 7.678401e-11, 
    7.741147e-11, 7.698604e-11, 7.77763e-11, 7.735142e-11, 7.780293e-11, 
    7.772095e-11, 7.785669e-11, 7.797826e-11, 7.813122e-11, 7.841343e-11, 
    7.834808e-11, 7.858411e-11, 7.617358e-11, 7.631811e-11, 7.63054e-11, 
    7.645666e-11, 7.656854e-11, 7.681102e-11, 7.719995e-11, 7.70537e-11, 
    7.732222e-11, 7.737612e-11, 7.696819e-11, 7.721863e-11, 7.641485e-11, 
    7.654469e-11, 7.646739e-11, 7.618497e-11, 7.708739e-11, 7.662424e-11, 
    7.747951e-11, 7.722859e-11, 7.796092e-11, 7.75967e-11, 7.831211e-11, 
    7.861793e-11, 7.890583e-11, 7.924222e-11, 7.639701e-11, 7.62988e-11, 
    7.647466e-11, 7.671795e-11, 7.694374e-11, 7.724389e-11, 7.727462e-11, 
    7.733084e-11, 7.747652e-11, 7.759899e-11, 7.734861e-11, 7.762969e-11, 
    7.657479e-11, 7.71276e-11, 7.626166e-11, 7.652238e-11, 7.670362e-11, 
    7.662412e-11, 7.703699e-11, 7.71343e-11, 7.752973e-11, 7.732532e-11, 
    7.854244e-11, 7.800392e-11, 7.949841e-11, 7.908072e-11, 7.626448e-11, 
    7.639667e-11, 7.685676e-11, 7.663785e-11, 7.726394e-11, 7.741806e-11, 
    7.754335e-11, 7.770351e-11, 7.772081e-11, 7.781571e-11, 7.76602e-11, 
    7.780956e-11, 7.724454e-11, 7.749703e-11, 7.680418e-11, 7.69728e-11, 
    7.689523e-11, 7.681014e-11, 7.707276e-11, 7.735255e-11, 7.735855e-11, 
    7.744826e-11, 7.770105e-11, 7.726648e-11, 7.861191e-11, 7.778094e-11, 
    7.654082e-11, 7.679544e-11, 7.683183e-11, 7.67332e-11, 7.740261e-11, 
    7.716004e-11, 7.781339e-11, 7.763681e-11, 7.792614e-11, 7.778237e-11, 
    7.776121e-11, 7.757656e-11, 7.74616e-11, 7.717116e-11, 7.693486e-11, 
    7.67475e-11, 7.679107e-11, 7.699688e-11, 7.736967e-11, 7.772237e-11, 
    7.764511e-11, 7.790416e-11, 7.721854e-11, 7.750602e-11, 7.73949e-11, 
    7.768464e-11, 7.704981e-11, 7.759034e-11, 7.691165e-11, 7.697116e-11, 
    7.715523e-11, 7.75255e-11, 7.760745e-11, 7.769492e-11, 7.764095e-11, 
    7.737914e-11, 7.733626e-11, 7.715076e-11, 7.709954e-11, 7.69582e-11, 
    7.684119e-11, 7.694809e-11, 7.706037e-11, 7.737926e-11, 7.766664e-11, 
    7.797998e-11, 7.805668e-11, 7.842277e-11, 7.812473e-11, 7.861654e-11, 
    7.819837e-11, 7.892228e-11, 7.762169e-11, 7.81861e-11, 7.716361e-11, 
    7.727376e-11, 7.747299e-11, 7.792997e-11, 7.768328e-11, 7.79718e-11, 
    7.733458e-11, 7.700398e-11, 7.691846e-11, 7.675889e-11, 7.692211e-11, 
    7.690884e-11, 7.706503e-11, 7.701484e-11, 7.738984e-11, 7.718841e-11, 
    7.776068e-11, 7.796952e-11, 7.855937e-11, 7.892098e-11, 7.928912e-11, 
    7.945165e-11, 7.950113e-11, 7.952181e-11 ;

 SOIL2C_vr =
  20.00587, 20.00588, 20.00588, 20.00589, 20.00588, 20.00589, 20.00587, 
    20.00588, 20.00587, 20.00587, 20.00592, 20.00589, 20.00594, 20.00593, 
    20.00597, 20.00594, 20.00597, 20.00597, 20.00598, 20.00598, 20.006, 
    20.00599, 20.00601, 20.006, 20.006, 20.00599, 20.0059, 20.00591, 20.0059, 
    20.0059, 20.0059, 20.00588, 20.00588, 20.00587, 20.00587, 20.00588, 
    20.0059, 20.00589, 20.00591, 20.00591, 20.00593, 20.00592, 20.00596, 
    20.00595, 20.00598, 20.00597, 20.00598, 20.00598, 20.00598, 20.00597, 
    20.00597, 20.00596, 20.00592, 20.00594, 20.0059, 20.00588, 20.00587, 
    20.00586, 20.00586, 20.00587, 20.00588, 20.00589, 20.0059, 20.00591, 
    20.00591, 20.00593, 20.00594, 20.00596, 20.00596, 20.00596, 20.00597, 
    20.00598, 20.00598, 20.00598, 20.00596, 20.00598, 20.00595, 20.00596, 
    20.00591, 20.00589, 20.00589, 20.00588, 20.00586, 20.00587, 20.00587, 
    20.00588, 20.00589, 20.00588, 20.00591, 20.0059, 20.00594, 20.00592, 
    20.00597, 20.00596, 20.00597, 20.00597, 20.00598, 20.00597, 20.00599, 
    20.00599, 20.00599, 20.006, 20.00597, 20.00598, 20.00588, 20.00588, 
    20.00589, 20.00588, 20.00587, 20.00587, 20.00587, 20.00588, 20.00589, 
    20.00589, 20.0059, 20.00591, 20.00593, 20.00595, 20.00596, 20.00597, 
    20.00596, 20.00597, 20.00596, 20.00596, 20.00599, 20.00597, 20.006, 
    20.00599, 20.00599, 20.00599, 20.00588, 20.00588, 20.00587, 20.00588, 
    20.00586, 20.00587, 20.00588, 20.0059, 20.0059, 20.00591, 20.00591, 
    20.00592, 20.00594, 20.00596, 20.00597, 20.00597, 20.00597, 20.00597, 
    20.00597, 20.00597, 20.00598, 20.00597, 20.00599, 20.00599, 20.00599, 
    20.00599, 20.00588, 20.00589, 20.00589, 20.00589, 20.00589, 20.0059, 
    20.00591, 20.00593, 20.00592, 20.00594, 20.00592, 20.00593, 20.00594, 
    20.00593, 20.00596, 20.00594, 20.00597, 20.00595, 20.00598, 20.00597, 
    20.00598, 20.00598, 20.00599, 20.006, 20.006, 20.00601, 20.0059, 20.0059, 
    20.0059, 20.00591, 20.00591, 20.00593, 20.00595, 20.00594, 20.00595, 
    20.00595, 20.00593, 20.00595, 20.00591, 20.00591, 20.00591, 20.0059, 
    20.00594, 20.00592, 20.00596, 20.00595, 20.00598, 20.00596, 20.006, 
    20.00601, 20.00603, 20.00604, 20.00591, 20.0059, 20.00591, 20.00592, 
    20.00593, 20.00595, 20.00595, 20.00595, 20.00596, 20.00596, 20.00595, 
    20.00597, 20.00591, 20.00594, 20.0059, 20.00591, 20.00592, 20.00592, 
    20.00594, 20.00594, 20.00596, 20.00595, 20.00601, 20.00599, 20.00606, 
    20.00604, 20.0059, 20.00591, 20.00593, 20.00592, 20.00595, 20.00596, 
    20.00596, 20.00597, 20.00597, 20.00598, 20.00597, 20.00598, 20.00595, 
    20.00596, 20.00593, 20.00594, 20.00593, 20.00593, 20.00594, 20.00595, 
    20.00595, 20.00596, 20.00597, 20.00595, 20.00601, 20.00597, 20.00591, 
    20.00593, 20.00593, 20.00592, 20.00595, 20.00594, 20.00598, 20.00597, 
    20.00598, 20.00597, 20.00597, 20.00596, 20.00596, 20.00595, 20.00593, 
    20.00592, 20.00593, 20.00594, 20.00595, 20.00597, 20.00597, 20.00598, 
    20.00595, 20.00596, 20.00595, 20.00597, 20.00594, 20.00596, 20.00593, 
    20.00593, 20.00594, 20.00596, 20.00597, 20.00597, 20.00597, 20.00595, 
    20.00595, 20.00594, 20.00594, 20.00593, 20.00593, 20.00593, 20.00594, 
    20.00595, 20.00597, 20.00598, 20.00599, 20.006, 20.00599, 20.00601, 
    20.00599, 20.00603, 20.00597, 20.00599, 20.00594, 20.00595, 20.00596, 
    20.00598, 20.00597, 20.00598, 20.00595, 20.00594, 20.00593, 20.00592, 
    20.00593, 20.00593, 20.00594, 20.00594, 20.00595, 20.00595, 20.00597, 
    20.00598, 20.00601, 20.00603, 20.00605, 20.00605, 20.00606, 20.00606,
  20.00534, 20.00536, 20.00535, 20.00537, 20.00536, 20.00537, 20.00534, 
    20.00536, 20.00535, 20.00534, 20.0054, 20.00537, 20.00543, 20.00541, 
    20.00546, 20.00543, 20.00547, 20.00546, 20.00549, 20.00548, 20.00551, 
    20.00549, 20.00552, 20.0055, 20.00551, 20.00549, 20.00538, 20.0054, 
    20.00537, 20.00538, 20.00538, 20.00536, 20.00535, 20.00534, 20.00534, 
    20.00535, 20.00538, 20.00537, 20.00539, 20.00539, 20.00542, 20.00541, 
    20.00546, 20.00544, 20.00548, 20.00547, 20.00548, 20.00548, 20.00548, 
    20.00546, 20.00547, 20.00546, 20.00541, 20.00542, 20.00538, 20.00536, 
    20.00534, 20.00533, 20.00533, 20.00533, 20.00535, 20.00537, 20.00538, 
    20.00539, 20.00539, 20.00542, 20.00543, 20.00546, 20.00545, 20.00546, 
    20.00547, 20.00548, 20.00548, 20.00549, 20.00546, 20.00548, 20.00545, 
    20.00546, 20.0054, 20.00537, 20.00536, 20.00535, 20.00533, 20.00535, 
    20.00534, 20.00536, 20.00537, 20.00536, 20.00539, 20.00538, 20.00543, 
    20.00541, 20.00547, 20.00545, 20.00547, 20.00546, 20.00548, 20.00546, 
    20.00549, 20.00549, 20.00549, 20.0055, 20.00546, 20.00548, 20.00536, 
    20.00536, 20.00536, 20.00535, 20.00535, 20.00533, 20.00535, 20.00535, 
    20.00537, 20.00537, 20.00538, 20.0054, 20.00541, 20.00544, 20.00546, 
    20.00547, 20.00546, 20.00546, 20.00546, 20.00546, 20.00549, 20.00547, 
    20.0055, 20.0055, 20.00549, 20.0055, 20.00536, 20.00536, 20.00534, 
    20.00535, 20.00533, 20.00535, 20.00535, 20.00538, 20.00538, 20.00539, 
    20.0054, 20.00541, 20.00543, 20.00545, 20.00547, 20.00547, 20.00547, 
    20.00547, 20.00546, 20.00547, 20.00548, 20.00547, 20.0055, 20.00549, 
    20.0055, 20.0055, 20.00536, 20.00537, 20.00536, 20.00537, 20.00536, 
    20.00538, 20.00539, 20.00542, 20.00541, 20.00543, 20.00541, 20.00541, 
    20.00543, 20.00541, 20.00545, 20.00542, 20.00547, 20.00545, 20.00547, 
    20.00547, 20.00548, 20.00549, 20.00549, 20.00551, 20.00551, 20.00552, 
    20.00537, 20.00538, 20.00538, 20.00539, 20.0054, 20.00541, 20.00544, 
    20.00543, 20.00545, 20.00545, 20.00542, 20.00544, 20.00539, 20.0054, 
    20.00539, 20.00538, 20.00543, 20.0054, 20.00546, 20.00544, 20.00548, 
    20.00546, 20.0055, 20.00552, 20.00554, 20.00556, 20.00539, 20.00538, 
    20.00539, 20.00541, 20.00542, 20.00544, 20.00544, 20.00545, 20.00546, 
    20.00546, 20.00545, 20.00546, 20.0054, 20.00543, 20.00538, 20.0054, 
    20.00541, 20.0054, 20.00543, 20.00543, 20.00546, 20.00545, 20.00552, 
    20.00549, 20.00558, 20.00555, 20.00538, 20.00539, 20.00542, 20.0054, 
    20.00544, 20.00545, 20.00546, 20.00547, 20.00547, 20.00547, 20.00546, 
    20.00547, 20.00544, 20.00546, 20.00541, 20.00542, 20.00542, 20.00541, 
    20.00543, 20.00545, 20.00545, 20.00545, 20.00547, 20.00544, 20.00552, 
    20.00547, 20.0054, 20.00541, 20.00541, 20.00541, 20.00545, 20.00544, 
    20.00547, 20.00546, 20.00548, 20.00547, 20.00547, 20.00546, 20.00545, 
    20.00544, 20.00542, 20.00541, 20.00541, 20.00542, 20.00545, 20.00547, 
    20.00546, 20.00548, 20.00544, 20.00546, 20.00545, 20.00547, 20.00543, 
    20.00546, 20.00542, 20.00542, 20.00543, 20.00546, 20.00546, 20.00547, 
    20.00546, 20.00545, 20.00545, 20.00543, 20.00543, 20.00542, 20.00542, 
    20.00542, 20.00543, 20.00545, 20.00547, 20.00549, 20.00549, 20.00551, 
    20.00549, 20.00552, 20.0055, 20.00554, 20.00546, 20.0055, 20.00544, 
    20.00544, 20.00546, 20.00548, 20.00547, 20.00548, 20.00545, 20.00543, 
    20.00542, 20.00541, 20.00542, 20.00542, 20.00543, 20.00543, 20.00545, 
    20.00544, 20.00547, 20.00548, 20.00552, 20.00554, 20.00556, 20.00557, 
    20.00558, 20.00558,
  20.00503, 20.00505, 20.00505, 20.00507, 20.00506, 20.00507, 20.00504, 
    20.00505, 20.00504, 20.00503, 20.0051, 20.00507, 20.00514, 20.00512, 
    20.00517, 20.00513, 20.00518, 20.00517, 20.00519, 20.00519, 20.00522, 
    20.0052, 20.00524, 20.00521, 20.00522, 20.0052, 20.00507, 20.0051, 
    20.00507, 20.00508, 20.00508, 20.00506, 20.00505, 20.00503, 20.00503, 
    20.00505, 20.00508, 20.00507, 20.00509, 20.00509, 20.00512, 20.00511, 
    20.00516, 20.00515, 20.00519, 20.00518, 20.00519, 20.00518, 20.00519, 
    20.00517, 20.00518, 20.00517, 20.00511, 20.00513, 20.00508, 20.00505, 
    20.00504, 20.00502, 20.00502, 20.00503, 20.00505, 20.00506, 20.00508, 
    20.00508, 20.00509, 20.00512, 20.00513, 20.00516, 20.00516, 20.00517, 
    20.00517, 20.00519, 20.00519, 20.00519, 20.00517, 20.00518, 20.00515, 
    20.00516, 20.0051, 20.00507, 20.00506, 20.00505, 20.00503, 20.00504, 
    20.00504, 20.00505, 20.00506, 20.00506, 20.00508, 20.00507, 20.00513, 
    20.00511, 20.00517, 20.00516, 20.00518, 20.00517, 20.00519, 20.00517, 
    20.0052, 20.0052, 20.0052, 20.00521, 20.00517, 20.00519, 20.00506, 
    20.00506, 20.00506, 20.00504, 20.00504, 20.00503, 20.00504, 20.00505, 
    20.00506, 20.00507, 20.00508, 20.00509, 20.00511, 20.00514, 20.00516, 
    20.00517, 20.00517, 20.00517, 20.00516, 20.00516, 20.0052, 20.00518, 
    20.00521, 20.00521, 20.00519, 20.00521, 20.00506, 20.00505, 20.00504, 
    20.00505, 20.00503, 20.00504, 20.00505, 20.00507, 20.00508, 20.00508, 
    20.0051, 20.00511, 20.00513, 20.00516, 20.00518, 20.00517, 20.00517, 
    20.00518, 20.00517, 20.00518, 20.00518, 20.00518, 20.00521, 20.0052, 
    20.00521, 20.0052, 20.00505, 20.00506, 20.00506, 20.00507, 20.00506, 
    20.00508, 20.00509, 20.00512, 20.00511, 20.00513, 20.00511, 20.00512, 
    20.00513, 20.00511, 20.00516, 20.00513, 20.00518, 20.00515, 20.00518, 
    20.00518, 20.00518, 20.00519, 20.0052, 20.00522, 20.00522, 20.00523, 
    20.00507, 20.00508, 20.00508, 20.00509, 20.0051, 20.00512, 20.00514, 
    20.00513, 20.00515, 20.00515, 20.00513, 20.00514, 20.00509, 20.0051, 
    20.00509, 20.00507, 20.00513, 20.0051, 20.00516, 20.00514, 20.00519, 
    20.00517, 20.00521, 20.00524, 20.00525, 20.00528, 20.00509, 20.00508, 
    20.00509, 20.00511, 20.00512, 20.00514, 20.00515, 20.00515, 20.00516, 
    20.00517, 20.00515, 20.00517, 20.0051, 20.00514, 20.00508, 20.0051, 
    20.00511, 20.0051, 20.00513, 20.00514, 20.00516, 20.00515, 20.00523, 
    20.0052, 20.00529, 20.00527, 20.00508, 20.00509, 20.00512, 20.0051, 
    20.00515, 20.00516, 20.00516, 20.00517, 20.00518, 20.00518, 20.00517, 
    20.00518, 20.00514, 20.00516, 20.00512, 20.00513, 20.00512, 20.00512, 
    20.00513, 20.00515, 20.00515, 20.00516, 20.00517, 20.00515, 20.00524, 
    20.00518, 20.0051, 20.00511, 20.00512, 20.00511, 20.00516, 20.00514, 
    20.00518, 20.00517, 20.00519, 20.00518, 20.00518, 20.00517, 20.00516, 
    20.00514, 20.00512, 20.00511, 20.00511, 20.00513, 20.00515, 20.00518, 
    20.00517, 20.00519, 20.00514, 20.00516, 20.00515, 20.00517, 20.00513, 
    20.00517, 20.00512, 20.00513, 20.00514, 20.00516, 20.00517, 20.00517, 
    20.00517, 20.00515, 20.00515, 20.00514, 20.00513, 20.00513, 20.00512, 
    20.00513, 20.00513, 20.00515, 20.00517, 20.00519, 20.0052, 20.00522, 
    20.0052, 20.00524, 20.00521, 20.00526, 20.00517, 20.00521, 20.00514, 
    20.00515, 20.00516, 20.00519, 20.00517, 20.00519, 20.00515, 20.00513, 
    20.00512, 20.00511, 20.00512, 20.00512, 20.00513, 20.00513, 20.00515, 
    20.00514, 20.00518, 20.00519, 20.00523, 20.00525, 20.00528, 20.00529, 
    20.00529, 20.00529,
  20.00479, 20.00481, 20.00481, 20.00483, 20.00482, 20.00483, 20.0048, 
    20.00481, 20.0048, 20.00479, 20.00486, 20.00483, 20.0049, 20.00488, 
    20.00493, 20.0049, 20.00494, 20.00493, 20.00496, 20.00495, 20.00498, 
    20.00496, 20.005, 20.00498, 20.00498, 20.00496, 20.00484, 20.00486, 
    20.00484, 20.00484, 20.00484, 20.00482, 20.00481, 20.00479, 20.00479, 
    20.00481, 20.00484, 20.00483, 20.00486, 20.00485, 20.00488, 20.00487, 
    20.00492, 20.00491, 20.00495, 20.00494, 20.00495, 20.00495, 20.00495, 
    20.00493, 20.00494, 20.00493, 20.00488, 20.00489, 20.00484, 20.00482, 
    20.0048, 20.00478, 20.00479, 20.00479, 20.00481, 20.00482, 20.00484, 
    20.00485, 20.00485, 20.00488, 20.00489, 20.00493, 20.00492, 20.00493, 
    20.00494, 20.00495, 20.00495, 20.00496, 20.00493, 20.00495, 20.00492, 
    20.00493, 20.00486, 20.00483, 20.00482, 20.00481, 20.00479, 20.0048, 
    20.0048, 20.00481, 20.00482, 20.00482, 20.00485, 20.00484, 20.0049, 
    20.00487, 20.00494, 20.00492, 20.00494, 20.00493, 20.00495, 20.00493, 
    20.00496, 20.00497, 20.00496, 20.00498, 20.00493, 20.00495, 20.00482, 
    20.00482, 20.00482, 20.0048, 20.0048, 20.00479, 20.0048, 20.00481, 
    20.00482, 20.00483, 20.00484, 20.00486, 20.00488, 20.0049, 20.00492, 
    20.00494, 20.00493, 20.00493, 20.00493, 20.00492, 20.00496, 20.00494, 
    20.00498, 20.00497, 20.00496, 20.00497, 20.00482, 20.00481, 20.0048, 
    20.00481, 20.00479, 20.0048, 20.00481, 20.00484, 20.00484, 20.00485, 
    20.00486, 20.00487, 20.0049, 20.00492, 20.00494, 20.00494, 20.00494, 
    20.00494, 20.00493, 20.00495, 20.00495, 20.00494, 20.00497, 20.00496, 
    20.00497, 20.00497, 20.00481, 20.00482, 20.00482, 20.00483, 20.00482, 
    20.00484, 20.00485, 20.00489, 20.00487, 20.00489, 20.00488, 20.00488, 
    20.00489, 20.00488, 20.00492, 20.00489, 20.00494, 20.00492, 20.00495, 
    20.00494, 20.00495, 20.00496, 20.00497, 20.00499, 20.00498, 20.005, 
    20.00483, 20.00484, 20.00484, 20.00485, 20.00486, 20.00488, 20.0049, 
    20.00489, 20.00491, 20.00492, 20.00489, 20.00491, 20.00485, 20.00486, 
    20.00485, 20.00484, 20.0049, 20.00487, 20.00492, 20.00491, 20.00496, 
    20.00493, 20.00498, 20.005, 20.00502, 20.00504, 20.00485, 20.00484, 
    20.00485, 20.00487, 20.00489, 20.00491, 20.00491, 20.00491, 20.00492, 
    20.00493, 20.00491, 20.00493, 20.00486, 20.0049, 20.00484, 20.00486, 
    20.00487, 20.00487, 20.00489, 20.0049, 20.00493, 20.00491, 20.005, 
    20.00496, 20.00506, 20.00503, 20.00484, 20.00485, 20.00488, 20.00487, 
    20.00491, 20.00492, 20.00493, 20.00494, 20.00494, 20.00495, 20.00494, 
    20.00495, 20.00491, 20.00492, 20.00488, 20.00489, 20.00488, 20.00488, 
    20.0049, 20.00492, 20.00492, 20.00492, 20.00494, 20.00491, 20.005, 
    20.00494, 20.00486, 20.00488, 20.00488, 20.00487, 20.00492, 20.0049, 
    20.00495, 20.00493, 20.00495, 20.00494, 20.00494, 20.00493, 20.00492, 
    20.0049, 20.00489, 20.00487, 20.00488, 20.00489, 20.00492, 20.00494, 
    20.00493, 20.00495, 20.00491, 20.00492, 20.00492, 20.00494, 20.00489, 
    20.00493, 20.00488, 20.00489, 20.0049, 20.00493, 20.00493, 20.00494, 
    20.00493, 20.00492, 20.00491, 20.0049, 20.0049, 20.00489, 20.00488, 
    20.00489, 20.00489, 20.00492, 20.00494, 20.00496, 20.00496, 20.00499, 
    20.00497, 20.005, 20.00497, 20.00502, 20.00493, 20.00497, 20.0049, 
    20.00491, 20.00492, 20.00495, 20.00494, 20.00496, 20.00491, 20.00489, 
    20.00488, 20.00487, 20.00488, 20.00488, 20.00489, 20.00489, 20.00492, 
    20.0049, 20.00494, 20.00496, 20.005, 20.00502, 20.00505, 20.00506, 
    20.00506, 20.00506,
  20.00426, 20.00427, 20.00427, 20.00429, 20.00428, 20.00429, 20.00426, 
    20.00428, 20.00426, 20.00426, 20.00432, 20.00429, 20.00435, 20.00433, 
    20.00438, 20.00435, 20.00438, 20.00438, 20.0044, 20.00439, 20.00442, 
    20.0044, 20.00444, 20.00442, 20.00442, 20.0044, 20.00429, 20.00431, 
    20.00429, 20.0043, 20.00429, 20.00428, 20.00427, 20.00425, 20.00426, 
    20.00427, 20.0043, 20.00429, 20.00431, 20.00431, 20.00434, 20.00433, 
    20.00437, 20.00436, 20.00439, 20.00438, 20.00439, 20.00439, 20.00439, 
    20.00438, 20.00439, 20.00437, 20.00433, 20.00434, 20.0043, 20.00428, 
    20.00426, 20.00425, 20.00425, 20.00425, 20.00427, 20.00428, 20.0043, 
    20.0043, 20.00431, 20.00433, 20.00434, 20.00437, 20.00437, 20.00438, 
    20.00438, 20.0044, 20.00439, 20.0044, 20.00438, 20.00439, 20.00437, 
    20.00437, 20.00431, 20.00429, 20.00428, 20.00427, 20.00425, 20.00426, 
    20.00426, 20.00427, 20.00428, 20.00428, 20.0043, 20.00429, 20.00435, 
    20.00432, 20.00438, 20.00437, 20.00439, 20.00438, 20.00439, 20.00438, 
    20.0044, 20.00441, 20.00441, 20.00442, 20.00438, 20.00439, 20.00428, 
    20.00428, 20.00428, 20.00427, 20.00427, 20.00425, 20.00426, 20.00427, 
    20.00428, 20.00429, 20.0043, 20.00431, 20.00433, 20.00435, 20.00437, 
    20.00438, 20.00437, 20.00438, 20.00437, 20.00437, 20.00441, 20.00439, 
    20.00442, 20.00442, 20.0044, 20.00442, 20.00428, 20.00427, 20.00426, 
    20.00427, 20.00425, 20.00426, 20.00427, 20.00429, 20.0043, 20.0043, 
    20.00431, 20.00433, 20.00435, 20.00437, 20.00438, 20.00438, 20.00438, 
    20.00439, 20.00438, 20.00439, 20.00439, 20.00439, 20.00442, 20.00441, 
    20.00442, 20.00441, 20.00428, 20.00428, 20.00428, 20.00429, 20.00428, 
    20.0043, 20.00431, 20.00434, 20.00433, 20.00434, 20.00433, 20.00433, 
    20.00434, 20.00433, 20.00437, 20.00434, 20.00439, 20.00436, 20.00439, 
    20.00438, 20.00439, 20.0044, 20.00441, 20.00443, 20.00442, 20.00444, 
    20.00429, 20.0043, 20.0043, 20.00431, 20.00432, 20.00433, 20.00435, 
    20.00434, 20.00436, 20.00436, 20.00434, 20.00435, 20.00431, 20.00431, 
    20.00431, 20.00429, 20.00435, 20.00432, 20.00437, 20.00435, 20.0044, 
    20.00438, 20.00442, 20.00444, 20.00446, 20.00448, 20.0043, 20.0043, 
    20.00431, 20.00432, 20.00434, 20.00436, 20.00436, 20.00436, 20.00437, 
    20.00438, 20.00436, 20.00438, 20.00432, 20.00435, 20.0043, 20.00431, 
    20.00432, 20.00432, 20.00434, 20.00435, 20.00437, 20.00436, 20.00443, 
    20.0044, 20.00449, 20.00447, 20.0043, 20.0043, 20.00433, 20.00432, 
    20.00436, 20.00437, 20.00437, 20.00438, 20.00438, 20.00439, 20.00438, 
    20.00439, 20.00436, 20.00437, 20.00433, 20.00434, 20.00434, 20.00433, 
    20.00435, 20.00436, 20.00436, 20.00437, 20.00438, 20.00436, 20.00444, 
    20.00439, 20.00431, 20.00433, 20.00433, 20.00433, 20.00437, 20.00435, 
    20.00439, 20.00438, 20.0044, 20.00439, 20.00439, 20.00438, 20.00437, 
    20.00435, 20.00434, 20.00433, 20.00433, 20.00434, 20.00436, 20.00438, 
    20.00438, 20.0044, 20.00435, 20.00437, 20.00437, 20.00438, 20.00434, 
    20.00438, 20.00434, 20.00434, 20.00435, 20.00437, 20.00438, 20.00438, 
    20.00438, 20.00436, 20.00436, 20.00435, 20.00435, 20.00434, 20.00433, 
    20.00434, 20.00434, 20.00436, 20.00438, 20.0044, 20.0044, 20.00443, 
    20.00441, 20.00444, 20.00441, 20.00446, 20.00438, 20.00441, 20.00435, 
    20.00436, 20.00437, 20.0044, 20.00438, 20.0044, 20.00436, 20.00434, 
    20.00434, 20.00433, 20.00434, 20.00434, 20.00434, 20.00434, 20.00436, 
    20.00435, 20.00439, 20.0044, 20.00443, 20.00446, 20.00448, 20.00449, 
    20.00449, 20.00449,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N =
  0.5258142, 0.5258147, 0.5258146, 0.525815, 0.5258148, 0.5258151, 0.5258143, 
    0.5258147, 0.5258144, 0.5258142, 0.5258159, 0.5258151, 0.5258167, 
    0.5258162, 0.5258176, 0.5258167, 0.5258178, 0.5258175, 0.5258182, 
    0.525818, 0.5258188, 0.5258182, 0.5258192, 0.5258186, 0.5258187, 
    0.5258182, 0.5258152, 0.5258158, 0.5258152, 0.5258152, 0.5258152, 
    0.5258148, 0.5258146, 0.5258141, 0.5258142, 0.5258145, 0.5258153, 
    0.5258151, 0.5258157, 0.5258157, 0.5258164, 0.5258161, 0.5258173, 
    0.525817, 0.525818, 0.5258178, 0.525818, 0.5258179, 0.525818, 0.5258176, 
    0.5258178, 0.5258175, 0.5258161, 0.5258166, 0.5258154, 0.5258147, 
    0.5258143, 0.525814, 0.525814, 0.5258141, 0.5258145, 0.525815, 0.5258152, 
    0.5258155, 0.5258157, 0.5258163, 0.5258167, 0.5258174, 0.5258173, 
    0.5258175, 0.5258177, 0.525818, 0.525818, 0.5258182, 0.5258175, 
    0.5258179, 0.5258172, 0.5258174, 0.5258157, 0.5258151, 0.5258148, 
    0.5258146, 0.5258141, 0.5258144, 0.5258143, 0.5258147, 0.5258149, 
    0.5258148, 0.5258155, 0.5258152, 0.5258167, 0.525816, 0.5258177, 
    0.5258173, 0.5258178, 0.5258175, 0.5258179, 0.5258176, 0.5258182, 
    0.5258184, 0.5258183, 0.5258186, 0.5258176, 0.525818, 0.5258148, 
    0.5258148, 0.5258149, 0.5258145, 0.5258145, 0.5258141, 0.5258144, 
    0.5258145, 0.5258149, 0.5258151, 0.5258153, 0.5258157, 0.5258162, 
    0.5258169, 0.5258173, 0.5258176, 0.5258175, 0.5258176, 0.5258174, 
    0.5258173, 0.5258183, 0.5258178, 0.5258186, 0.5258186, 0.5258182, 
    0.5258186, 0.5258148, 0.5258147, 0.5258143, 0.5258146, 0.5258141, 
    0.5258144, 0.5258145, 0.5258152, 0.5258154, 0.5258155, 0.5258158, 
    0.5258161, 0.5258167, 0.5258172, 0.5258177, 0.5258177, 0.5258177, 
    0.5258178, 0.5258175, 0.5258179, 0.5258179, 0.5258178, 0.5258185, 
    0.5258183, 0.5258186, 0.5258184, 0.5258147, 0.5258149, 0.5258148, 
    0.525815, 0.5258149, 0.5258154, 0.5258156, 0.5258164, 0.5258161, 
    0.5258166, 0.5258161, 0.5258163, 0.5258167, 0.5258162, 0.5258172, 
    0.5258165, 0.5258178, 0.5258171, 0.5258179, 0.5258177, 0.5258179, 
    0.5258182, 0.5258184, 0.5258188, 0.5258188, 0.5258191, 0.5258152, 
    0.5258154, 0.5258154, 0.5258157, 0.5258158, 0.5258162, 0.5258169, 
    0.5258166, 0.525817, 0.5258172, 0.5258165, 0.5258169, 0.5258156, 
    0.5258158, 0.5258157, 0.5258152, 0.5258167, 0.5258159, 0.5258173, 
    0.5258169, 0.5258181, 0.5258175, 0.5258187, 0.5258192, 0.5258197, 
    0.5258202, 0.5258155, 0.5258154, 0.5258157, 0.5258161, 0.5258164, 
    0.5258169, 0.525817, 0.5258171, 0.5258173, 0.5258175, 0.5258171, 
    0.5258176, 0.5258158, 0.5258167, 0.5258153, 0.5258158, 0.525816, 
    0.5258159, 0.5258166, 0.5258167, 0.5258174, 0.5258171, 0.5258191, 
    0.5258182, 0.5258206, 0.52582, 0.5258153, 0.5258155, 0.5258163, 0.525816, 
    0.525817, 0.5258172, 0.5258175, 0.5258177, 0.5258177, 0.5258179, 
    0.5258176, 0.5258179, 0.5258169, 0.5258173, 0.5258162, 0.5258165, 
    0.5258164, 0.5258162, 0.5258167, 0.5258171, 0.5258171, 0.5258173, 
    0.5258177, 0.525817, 0.5258192, 0.5258178, 0.5258158, 0.5258162, 
    0.5258163, 0.5258161, 0.5258172, 0.5258168, 0.5258179, 0.5258176, 
    0.525818, 0.5258178, 0.5258178, 0.5258175, 0.5258173, 0.5258168, 
    0.5258164, 0.5258161, 0.5258162, 0.5258166, 0.5258172, 0.5258177, 
    0.5258176, 0.525818, 0.5258169, 0.5258174, 0.5258172, 0.5258176, 
    0.5258166, 0.5258175, 0.5258164, 0.5258165, 0.5258168, 0.5258174, 
    0.5258175, 0.5258177, 0.5258176, 0.5258172, 0.5258171, 0.5258168, 
    0.5258167, 0.5258164, 0.5258163, 0.5258164, 0.5258166, 0.5258172, 
    0.5258176, 0.5258182, 0.5258183, 0.5258189, 0.5258184, 0.5258192, 
    0.5258185, 0.5258197, 0.5258176, 0.5258185, 0.5258168, 0.525817, 
    0.5258173, 0.525818, 0.5258176, 0.5258181, 0.5258171, 0.5258166, 
    0.5258164, 0.5258161, 0.5258164, 0.5258164, 0.5258166, 0.5258166, 
    0.5258172, 0.5258169, 0.5258178, 0.5258181, 0.5258191, 0.5258197, 
    0.5258203, 0.5258206, 0.5258206, 0.5258207 ;

 SOIL2N_TNDNCY_VERT_TRANS =
  -2.569961e-21, -1.027984e-20, 2.569961e-21, 2.569961e-21, -1.541976e-20, 
    -5.139921e-21, 2.569961e-21, -7.709882e-21, -2.569961e-21, 1.28498e-20, 
    -7.709882e-21, -5.139921e-21, 1.027984e-20, -1.027984e-20, 1.541976e-20, 
    -1.027984e-20, 2.569961e-21, -1.027984e-20, -2.569961e-21, -1.027984e-20, 
    -7.709882e-21, 1.003089e-36, -1.28498e-20, 1.003089e-36, 1.027984e-20, 
    -2.569961e-21, -5.139921e-21, -7.709882e-21, -1.003089e-36, 
    -2.569961e-21, 1.798972e-20, -7.709882e-21, -1.003089e-36, 0, 
    7.709882e-21, -5.139921e-21, -1.28498e-20, -1.541976e-20, 1.541976e-20, 
    0, 5.139921e-21, -1.027984e-20, 5.139921e-21, -2.569961e-21, 
    -1.28498e-20, -5.139921e-21, -1.28498e-20, 1.28498e-20, 5.139921e-21, 
    -7.709882e-21, 2.569961e-21, -1.027984e-20, -1.798972e-20, -1.798972e-20, 
    5.139921e-21, 1.003089e-36, 1.003089e-36, 7.709882e-21, 1.027984e-20, 
    7.709882e-21, -1.798972e-20, -1.28498e-20, 2.569961e-21, 1.003089e-36, 
    -2.569961e-21, -2.569961e-21, 7.709882e-21, 1.027984e-20, 2.055969e-20, 
    -7.709882e-21, 1.28498e-20, -5.139921e-21, 1.003089e-36, 1.28498e-20, 
    2.569961e-21, 1.027984e-20, 1.027984e-20, 2.569961e-21, -7.709882e-21, 
    -1.027984e-20, 7.709882e-21, -5.139921e-21, 1.027984e-20, 1.798972e-20, 
    5.139921e-21, -1.003089e-36, -2.569961e-21, -1.28498e-20, 2.569961e-21, 
    0, -5.139921e-21, -1.541976e-20, -1.28498e-20, 7.709882e-21, 
    5.139921e-21, -7.709882e-21, -1.28498e-20, -2.569961e-21, -2.569961e-21, 
    -5.139921e-21, 1.798972e-20, -2.569961e-21, -1.798972e-20, 7.709882e-21, 
    5.139921e-21, -2.569961e-21, -5.139921e-21, 1.28498e-20, 0, 1.027984e-20, 
    -2.569961e-21, 2.569961e-21, 1.28498e-20, 5.139921e-21, 2.569961e-21, 
    2.569961e-21, -2.569961e-21, -2.569961e-20, 1.798972e-20, -7.709882e-21, 
    2.569961e-21, 1.027984e-20, -2.569961e-21, 7.709882e-21, -7.709882e-21, 
    -5.139921e-21, -1.027984e-20, 1.28498e-20, -1.28498e-20, 1.027984e-20, 
    -5.139921e-21, 2.569961e-21, -1.28498e-20, 1.027984e-20, 1.027984e-20, 
    -7.709882e-21, 2.569961e-21, -5.139921e-21, -2.569961e-21, 2.569961e-21, 
    1.541976e-20, 5.139921e-21, -5.139921e-21, 1.28498e-20, -1.28498e-20, 0, 
    1.003089e-36, -1.28498e-20, 2.569961e-21, -2.569961e-20, -1.003089e-36, 
    2.569961e-21, 0, -7.709882e-21, 1.541976e-20, 1.027984e-20, 
    -2.569961e-21, 1.027984e-20, 7.709882e-21, -5.139921e-21, 7.709882e-21, 
    2.569961e-21, 2.569961e-21, 5.139921e-21, -7.709882e-21, 2.312965e-20, 
    2.569961e-21, -1.541976e-20, -1.003089e-36, 2.569961e-21, -2.569961e-21, 
    -2.569961e-21, -1.027984e-20, 0, 2.569961e-21, 1.541976e-20, 
    -2.569961e-21, -2.569961e-21, 1.541976e-20, 7.709882e-21, 1.027984e-20, 
    7.709882e-21, 5.139921e-21, 7.709882e-21, -1.28498e-20, -1.003089e-36, 
    -2.569961e-21, 2.312965e-20, 5.139921e-21, 1.28498e-20, 7.709882e-21, 
    5.139921e-21, 1.003089e-36, -1.798972e-20, 2.569961e-21, 0, 
    -2.569961e-21, -7.709882e-21, -2.312965e-20, -1.003089e-36, 
    -7.709882e-21, 1.027984e-20, -2.569961e-21, -1.798972e-20, 7.709882e-21, 
    -1.28498e-20, 1.027984e-20, 5.139921e-21, -5.139921e-21, -5.139921e-21, 
    1.28498e-20, 5.139921e-21, -1.28498e-20, 2.569961e-21, 7.709882e-21, 
    1.541976e-20, -1.003089e-36, -5.139921e-21, 5.139921e-21, -1.027984e-20, 
    5.139921e-21, 7.709882e-21, 1.003089e-36, 5.139921e-21, 1.28498e-20, 
    -1.027984e-20, -1.003089e-36, -2.569961e-21, 1.28498e-20, -7.709882e-21, 
    5.139921e-21, -7.709882e-21, 5.139921e-21, 0, 7.709882e-21, 0, 
    1.541976e-20, -1.28498e-20, 5.139921e-21, 5.139921e-21, -2.569961e-21, 
    -5.139921e-21, -1.027984e-20, -1.027984e-20, -5.139921e-21, 
    -7.709882e-21, 1.003089e-36, 2.826957e-20, 1.798972e-20, 0, -1.28498e-20, 
    7.709882e-21, 0, -2.569961e-21, 2.569961e-21, 2.569961e-21, 
    -1.003089e-36, -2.569961e-21, 5.139921e-21, -1.003089e-36, -5.139921e-21, 
    7.709882e-21, -2.569961e-21, -1.28498e-20, -1.027984e-20, -1.003089e-36, 
    1.798972e-20, 2.569961e-21, -1.798972e-20, -1.027984e-20, 0, 
    2.569961e-21, 2.312965e-20, -7.709882e-21, -1.541976e-20, 1.003089e-36, 
    -2.569961e-21, 1.28498e-20, 2.569961e-21, 2.569961e-21, 1.027984e-20, 
    2.569961e-21, -1.027984e-20, 2.569961e-21, 1.798972e-20, 7.709882e-21, 
    -1.027984e-20, -7.709882e-21, 5.139921e-21, -5.139921e-21, 1.003089e-36, 
    -7.709882e-21, 2.569961e-21, 5.139921e-21, -2.569961e-21, 5.139921e-21, 
    5.139921e-21, 2.569961e-21, -2.569961e-21, -1.541976e-20, 7.709882e-21, 
    2.569961e-21, 5.139921e-21, -1.798972e-20, -1.28498e-20, -2.569961e-21, 
    -1.28498e-20, -1.541976e-20, -2.569961e-21, -2.569961e-20, -7.709882e-21, 
    -2.569961e-21, 0, -5.139921e-21, 7.709882e-21, 2.569961e-21, 
    -1.28498e-20, 7.709882e-21, 1.798972e-20, 1.027984e-20, -1.541976e-20, 
    5.139921e-21, 2.569961e-21, 5.139921e-21, 2.569961e-21, 1.027984e-20, 
    2.055969e-20, 5.139921e-21, 5.139921e-21, -2.569961e-21, -5.139921e-21, 
    -1.027984e-20, 5.139921e-21, -2.569961e-21, -1.28498e-20, -2.569961e-21, 
    -1.28498e-20, 5.139921e-21,
  -5.139921e-21, 2.569961e-21, -2.569961e-21, -5.139921e-21, -7.709882e-21, 
    -7.709882e-21, -7.709882e-21, 0, -7.709882e-21, 1.027984e-20, 
    7.709882e-21, -7.709882e-21, 7.709882e-21, 2.569961e-21, 2.569961e-21, 
    2.569961e-21, -7.709882e-21, 2.569961e-21, -2.569961e-21, 0, 1.28498e-20, 
    -7.709882e-21, -2.569961e-21, 1.027984e-20, 7.709882e-21, 7.709882e-21, 
    -5.139921e-21, 7.709882e-21, -5.139921e-21, 0, 2.569961e-21, 
    2.569961e-21, 5.139921e-21, 2.569961e-21, 7.709882e-21, 2.569961e-21, 
    2.569961e-21, 5.139921e-21, -5.139921e-21, -5.139921e-21, -2.569961e-21, 
    -1.027984e-20, -2.569961e-21, 2.569961e-21, 2.569961e-21, -2.569961e-21, 
    1.003089e-36, 7.709882e-21, -5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, 1.027984e-20, -5.139921e-21, 2.569961e-21, -1.027984e-20, 
    2.569961e-21, 1.541976e-20, -1.027984e-20, -1.027984e-20, 7.709882e-21, 
    -5.139921e-21, -7.709882e-21, -1.541976e-20, -7.709882e-21, 
    -7.709882e-21, -2.569961e-21, -2.569961e-21, 7.709882e-21, -1.027984e-20, 
    2.569961e-21, 0, -5.139921e-21, 1.027984e-20, -7.709882e-21, 
    2.569961e-21, 2.569961e-21, -7.709882e-21, -5.139921e-21, 2.569961e-21, 
    -5.139921e-21, -2.569961e-21, -2.569961e-21, -1.027984e-20, 0, 
    -1.027984e-20, 7.709882e-21, 5.139921e-21, -1.28498e-20, 1.541976e-20, 
    5.139921e-21, 1.28498e-20, -5.139921e-21, 2.569961e-21, 5.139921e-21, 
    7.709882e-21, -5.139921e-21, -1.027984e-20, 2.569961e-21, 5.139921e-21, 
    -7.709882e-21, 1.003089e-36, 7.709882e-21, -7.709882e-21, -1.027984e-20, 
    -2.569961e-21, -2.055969e-20, -5.139921e-21, 0, 7.709882e-21, 
    -1.027984e-20, 2.569961e-21, 2.569961e-21, 7.709882e-21, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, -7.709882e-21, -2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 5.139921e-21, 1.027984e-20, 2.569961e-21, 0, 
    -5.139921e-21, 0, 5.139921e-21, -2.569961e-21, 1.027984e-20, 
    -5.139921e-21, 7.709882e-21, 1.541976e-20, -2.569961e-21, 2.569961e-21, 
    -7.709882e-21, -2.312965e-20, -1.28498e-20, -2.569961e-21, -2.569961e-21, 
    7.709882e-21, -1.541976e-20, 2.569961e-21, 5.139921e-21, 1.28498e-20, 
    2.569961e-21, -7.709882e-21, -7.709882e-21, 7.709882e-21, 2.569961e-21, 
    5.139921e-21, -2.569961e-21, -7.709882e-21, 1.027984e-20, 5.139921e-21, 
    2.569961e-21, 2.569961e-21, 0, 1.027984e-20, -1.003089e-36, -1.28498e-20, 
    5.139921e-21, -5.139921e-21, 1.003089e-36, 5.139921e-21, 7.709882e-21, 
    -2.569961e-21, 2.569961e-21, -7.709882e-21, -1.28498e-20, -7.709882e-21, 
    0, 7.709882e-21, -5.139921e-21, 0, -1.027984e-20, 1.28498e-20, 
    -2.569961e-21, -5.139921e-21, 7.709882e-21, -1.027984e-20, 2.569961e-21, 
    -5.139921e-21, -1.003089e-36, 2.569961e-21, -2.569961e-21, 0, 
    -2.569961e-21, -7.709882e-21, -2.569961e-21, -2.569961e-21, 
    -5.139921e-21, 1.541976e-20, 7.709882e-21, 2.569961e-21, -2.569961e-21, 
    2.569961e-21, 0, -1.541976e-20, 2.569961e-21, 0, 2.569961e-21, 0, 
    1.798972e-20, 0, -2.569961e-21, 7.709882e-21, -5.139921e-21, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, 2.569961e-21, 0, 0, 
    1.541976e-20, 7.709882e-21, -2.569961e-21, -5.139921e-21, 2.569961e-21, 
    2.569961e-21, -2.569961e-21, 2.569961e-21, 2.569961e-21, -7.709882e-21, 
    0, -2.569961e-21, 1.003089e-36, 0, -5.139921e-21, -1.027984e-20, 
    -7.709882e-21, -1.28498e-20, -2.569961e-21, 5.139921e-21, -5.139921e-21, 
    -2.569961e-21, -1.28498e-20, 2.569961e-21, -2.569961e-21, 5.139921e-21, 
    -2.569961e-21, -2.569961e-21, 1.541976e-20, 0, 5.139921e-21, 
    1.541976e-20, 2.569961e-21, 5.139921e-21, -1.28498e-20, -7.709882e-21, 
    -5.139921e-21, -2.569961e-21, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, 1.027984e-20, -1.027984e-20, 5.139921e-21, -2.569961e-21, 
    -2.569961e-21, 5.139921e-21, -2.569961e-21, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, 0, -7.709882e-21, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, -1.28498e-20, -2.569961e-21, 0, 
    -7.709882e-21, -1.541976e-20, -2.569961e-21, 0, 2.569961e-21, 
    2.569961e-21, -1.027984e-20, -2.569961e-21, -1.003089e-36, 1.027984e-20, 
    0, -7.709882e-21, -2.569961e-21, -5.139921e-21, 5.139921e-21, 
    -7.709882e-21, 7.709882e-21, -2.569961e-21, -2.569961e-21, -1.28498e-20, 
    2.569961e-21, -2.569961e-21, 5.139921e-21, -5.139921e-21, 1.027984e-20, 
    -1.027984e-20, 7.709882e-21, -7.709882e-21, -7.709882e-21, 5.139921e-21, 
    0, -5.139921e-21, 1.28498e-20, -5.139921e-21, -1.027984e-20, 
    -1.027984e-20, 5.139921e-21, -7.709882e-21, -1.28498e-20, 1.027984e-20, 
    5.139921e-21, 2.569961e-21, -5.139921e-21, 2.569961e-21, -1.027984e-20, 
    -1.28498e-20, 2.569961e-21, -2.569961e-21, 2.569961e-21, 0, 2.569961e-21, 
    -7.709882e-21, -1.28498e-20, -7.709882e-21, 5.139921e-21, 0, 
    1.541976e-20, 1.28498e-20, 2.569961e-21, 2.569961e-21, -2.569961e-21, 
    1.798972e-20, 1.798972e-20,
  1.003089e-36, -2.569961e-21, -1.027984e-20, -5.139921e-21, 1.003089e-36, 
    2.569961e-21, -5.139921e-21, 5.139921e-21, 2.569961e-21, 1.28498e-20, 
    2.569961e-21, -5.139921e-21, -7.709882e-21, 1.027984e-20, -5.139921e-21, 
    -5.139921e-21, 2.055969e-20, -7.709882e-21, 2.569961e-21, -5.139921e-21, 
    -2.569961e-21, 5.139921e-21, 1.027984e-20, 2.569961e-21, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, -5.139921e-21, -5.139921e-21, 
    -1.798972e-20, 5.139921e-21, -7.709882e-21, -5.139921e-21, 2.569961e-21, 
    -7.709882e-21, 2.569961e-21, 1.027984e-20, 1.003089e-36, 2.569961e-21, 
    2.569961e-21, 5.139921e-21, -2.569961e-21, 1.027984e-20, -1.541976e-20, 
    1.027984e-20, 5.139921e-21, -1.027984e-20, -1.027984e-20, 5.139921e-21, 
    5.139921e-21, 7.709882e-21, 2.569961e-21, -2.569961e-21, -5.139921e-21, 
    -2.569961e-21, 0, -1.003089e-36, 2.569961e-21, 1.027984e-20, 
    -5.139921e-21, -1.027984e-20, -5.139921e-21, 2.569961e-21, -1.798972e-20, 
    2.569961e-21, 2.569961e-21, -7.709882e-21, -7.709882e-21, -1.027984e-20, 
    1.28498e-20, -1.003089e-36, -2.569961e-21, 2.569961e-21, -5.139921e-21, 
    0, -1.28498e-20, 1.027984e-20, 2.569961e-21, 1.027984e-20, 1.027984e-20, 
    1.541976e-20, 7.709882e-21, 1.003089e-36, -5.139921e-21, -5.139921e-21, 
    -7.709882e-21, 0, 5.139921e-21, 5.139921e-21, 2.569961e-20, 2.569961e-21, 
    1.541976e-20, 5.139921e-21, 1.003089e-36, 7.709882e-21, 7.709882e-21, 
    5.139921e-21, 7.709882e-21, -1.28498e-20, -5.139921e-21, 2.569961e-21, 
    2.569961e-21, -5.139921e-21, -2.569961e-21, -2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 2.569961e-21, 1.541976e-20, 5.139921e-21, -7.709882e-21, 
    -1.798972e-20, 5.139921e-21, 2.569961e-21, -7.709882e-21, 2.569961e-21, 
    -1.003089e-36, -2.569961e-21, -1.28498e-20, -2.312965e-20, 7.709882e-21, 
    2.569961e-21, -2.569961e-21, 1.003089e-36, -2.569961e-21, -2.569961e-21, 
    5.139921e-21, 7.709882e-21, -2.569961e-21, 1.027984e-20, -1.027984e-20, 
    -2.569961e-21, -2.569961e-21, -1.798972e-20, -5.139921e-21, 
    -7.709882e-21, -2.569961e-21, 2.569961e-21, -1.027984e-20, 1.28498e-20, 
    1.28498e-20, -1.003089e-36, 2.569961e-21, 2.569961e-21, -2.569961e-21, 
    2.055969e-20, 1.003089e-36, -1.541976e-20, 5.139921e-21, -2.569961e-21, 
    0, -1.798972e-20, 1.28498e-20, 7.709882e-21, -2.569961e-21, -1.28498e-20, 
    -1.003089e-36, -5.139921e-21, -2.569961e-21, -5.139921e-21, 7.709882e-21, 
    -5.139921e-21, -5.139921e-21, -5.139921e-21, -5.139921e-21, 
    -1.027984e-20, 2.569961e-21, 1.003089e-36, 1.28498e-20, 2.569961e-21, 
    -1.541976e-20, -1.027984e-20, -2.569961e-21, -7.709882e-21, 0, 
    1.027984e-20, -7.709882e-21, -1.027984e-20, -5.139921e-21, 1.541976e-20, 
    -1.003089e-36, -7.709882e-21, 2.569961e-21, 7.709882e-21, -2.569961e-21, 
    5.139921e-21, 1.027984e-20, 5.139921e-21, -5.139921e-21, 5.139921e-21, 
    5.139921e-21, 7.709882e-21, -5.139921e-21, 1.28498e-20, 7.709882e-21, 
    5.139921e-21, -5.139921e-21, 5.139921e-21, -5.139921e-21, 7.709882e-21, 
    -2.569961e-21, 5.139921e-21, 2.569961e-21, -7.709882e-21, -1.027984e-20, 
    5.139921e-21, -7.709882e-21, 0, 1.28498e-20, 1.027984e-20, -1.798972e-20, 
    1.541976e-20, -5.139921e-21, 1.027984e-20, 7.709882e-21, -7.709882e-21, 
    -5.139921e-21, -1.027984e-20, -2.569961e-21, 2.569961e-21, -5.139921e-21, 
    7.709882e-21, -2.569961e-21, 2.569961e-21, -7.709882e-21, 1.798972e-20, 
    2.569961e-21, -7.709882e-21, 7.709882e-21, 1.027984e-20, -1.541976e-20, 
    2.569961e-21, 2.569961e-21, -7.709882e-21, -7.709882e-21, -7.709882e-21, 
    0, 0, -2.569961e-21, 5.139921e-21, -2.569961e-21, -1.003089e-36, 
    -2.569961e-21, 5.139921e-21, 7.709882e-21, 7.709882e-21, 1.027984e-20, 
    5.139921e-21, -5.139921e-21, 7.709882e-21, 0, -7.709882e-21, 
    7.709882e-21, -2.569961e-21, 5.139921e-21, 1.003089e-36, -1.28498e-20, 
    5.139921e-21, -7.709882e-21, 0, -7.709882e-21, 1.28498e-20, 1.28498e-20, 
    1.027984e-20, -5.139921e-21, -2.569961e-21, -7.709882e-21, 5.139921e-21, 
    -7.709882e-21, 1.28498e-20, 7.709882e-21, -1.541976e-20, -2.569961e-21, 
    -2.569961e-21, -2.569961e-21, -5.139921e-21, 0, 5.139921e-21, 0, 
    -5.139921e-21, -2.569961e-21, 2.569961e-21, -7.709882e-21, 5.139921e-21, 
    1.541976e-20, -2.569961e-21, -5.139921e-21, 0, -7.709882e-21, 
    1.027984e-20, 2.569961e-21, -1.027984e-20, 1.28498e-20, -1.28498e-20, 
    -5.139921e-21, 1.28498e-20, -7.709882e-21, -2.569961e-21, 1.28498e-20, 
    2.569961e-21, -5.139921e-21, 5.139921e-21, -1.027984e-20, -2.569961e-21, 
    2.569961e-21, 7.709882e-21, -1.027984e-20, -5.139921e-21, 1.541976e-20, 
    5.139921e-21, 5.139921e-21, 5.139921e-21, 7.709882e-21, -5.139921e-21, 
    2.569961e-21, -7.709882e-21, -1.027984e-20, 2.569961e-21, -1.798972e-20, 
    5.139921e-21, 2.569961e-21, -2.569961e-21, -2.569961e-20, 7.709882e-21, 
    5.139921e-21, 1.027984e-20, 0, 1.027984e-20, -5.139921e-21, 2.569961e-21, 
    -7.709882e-21, 0, 2.312965e-20, 2.569961e-21, -5.139921e-21, 
    -1.541976e-20, -5.139921e-21, -1.541976e-20,
  2.569961e-21, -5.139921e-21, -2.055969e-20, -2.569961e-21, 2.569961e-21, 
    -1.28498e-20, 1.027984e-20, -5.139921e-21, 2.569961e-21, -2.569961e-21, 
    -5.139921e-21, 1.541976e-20, -2.569961e-21, -1.027984e-20, 0, 
    5.139921e-21, 2.569961e-21, -1.027984e-20, -5.139921e-21, 2.569961e-21, 
    -1.541976e-20, -7.709882e-21, 2.569961e-21, -1.003089e-36, -2.569961e-21, 
    2.569961e-21, -7.709882e-21, 2.569961e-21, 2.569961e-21, 7.709882e-21, 
    1.798972e-20, 5.139921e-21, -5.139921e-21, -1.027984e-20, 7.709882e-21, 
    -1.003089e-36, -7.709882e-21, -1.28498e-20, -1.003089e-36, -1.28498e-20, 
    0, -2.569961e-21, -5.139921e-21, 0, -7.709882e-21, -2.055969e-20, 
    2.569961e-21, 7.709882e-21, 0, 7.709882e-21, 1.28498e-20, -5.139921e-21, 
    -1.541976e-20, -2.569961e-21, -2.569961e-21, 5.139921e-21, -2.569961e-21, 
    -1.027984e-20, -1.027984e-20, 2.569961e-21, -1.003089e-36, 1.28498e-20, 
    -1.003089e-36, 1.027984e-20, 5.139921e-21, -2.569961e-21, 7.709882e-21, 
    -2.569961e-21, -2.569961e-21, -2.312965e-20, 1.28498e-20, -2.569961e-21, 
    -2.569961e-21, -2.569961e-21, 1.027984e-20, 1.28498e-20, 1.027984e-20, 0, 
    -1.027984e-20, -1.28498e-20, -5.139921e-21, 5.139921e-21, 7.709882e-21, 
    -7.709882e-21, -7.709882e-21, -1.541976e-20, 2.055969e-20, -7.709882e-21, 
    1.003089e-36, 1.027984e-20, -5.139921e-21, 0, 5.139921e-21, 
    -1.541976e-20, -7.709882e-21, 5.139921e-21, 7.709882e-21, 7.709882e-21, 
    1.003089e-36, -1.027984e-20, -1.798972e-20, 0, -1.027984e-20, 
    1.027984e-20, -5.139921e-21, 2.055969e-20, 0, 1.027984e-20, 1.28498e-20, 
    -7.709882e-21, 1.027984e-20, 0, -7.709882e-21, -5.139921e-21, 
    1.003089e-36, 7.709882e-21, 5.139921e-21, 2.569961e-21, 1.003089e-36, 0, 
    2.569961e-21, -2.569961e-21, -2.312965e-20, 2.569961e-21, 1.027984e-20, 
    1.28498e-20, 2.569961e-21, -2.569961e-21, -1.28498e-20, 0, 2.569961e-21, 
    -2.569961e-21, -7.709882e-21, 7.709882e-21, 2.569961e-21, 5.139921e-21, 
    2.569961e-21, 2.312965e-20, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    1.003089e-36, -7.709882e-21, -1.28498e-20, 1.28498e-20, -1.541976e-20, 
    1.798972e-20, -1.003089e-36, 2.569961e-21, -7.709882e-21, -5.139921e-21, 
    2.569961e-21, 1.28498e-20, -5.139921e-21, -7.709882e-21, -7.709882e-21, 
    5.139921e-21, -1.027984e-20, 1.28498e-20, -5.139921e-21, 2.569961e-21, 
    7.709882e-21, -7.709882e-21, -7.709882e-21, 0, -1.027984e-20, 
    -5.139921e-21, 1.28498e-20, -5.139921e-21, -1.027984e-20, -1.027984e-20, 
    -7.709882e-21, 1.798972e-20, 7.709882e-21, -5.139921e-21, 7.709882e-21, 
    -1.541976e-20, -1.541976e-20, -1.027984e-20, 7.709882e-21, 5.139921e-21, 
    1.003089e-36, 1.027984e-20, 7.709882e-21, -5.139921e-21, 1.027984e-20, 
    -7.709882e-21, 1.28498e-20, -1.541976e-20, -5.139921e-21, -1.28498e-20, 
    -2.569961e-21, -1.541976e-20, -1.027984e-20, -2.569961e-21, 
    -7.709882e-21, 2.569961e-21, 1.798972e-20, 5.139921e-21, -1.541976e-20, 
    1.28498e-20, -2.055969e-20, -1.541976e-20, -5.139921e-21, 1.003089e-36, 
    -1.28498e-20, -1.28498e-20, 7.709882e-21, 2.569961e-21, -2.569961e-21, 
    -2.569961e-21, 0, -1.28498e-20, 7.709882e-21, -5.139921e-21, 
    -1.027984e-20, 2.569961e-21, 7.709882e-21, -1.003089e-36, -1.28498e-20, 
    1.027984e-20, 2.569961e-21, 5.139921e-21, -2.569961e-21, -7.709882e-21, 
    1.28498e-20, -1.003089e-36, -5.139921e-21, 5.139921e-21, 2.569961e-21, 
    1.027984e-20, 7.709882e-21, 2.055969e-20, -5.139921e-21, 0, 
    -5.139921e-21, -7.709882e-21, 0, 3.340949e-20, 7.709882e-21, 
    -5.139921e-21, 5.139921e-21, -1.541976e-20, -1.28498e-20, 5.139921e-21, 
    5.139921e-21, 5.139921e-21, -7.709882e-21, -2.569961e-21, 1.027984e-20, 
    -1.28498e-20, -5.139921e-21, -2.569961e-21, 1.541976e-20, -2.569961e-21, 
    -7.709882e-21, 2.569961e-21, -2.569961e-21, 1.027984e-20, 1.027984e-20, 
    1.798972e-20, 0, -2.569961e-21, -1.28498e-20, 2.569961e-21, 
    -1.003089e-36, 1.027984e-20, -7.709882e-21, -2.569961e-21, -2.569961e-21, 
    -1.28498e-20, 2.569961e-21, -7.709882e-21, -1.003089e-36, 1.541976e-20, 
    -5.139921e-21, 1.28498e-20, -1.28498e-20, 0, 1.027984e-20, -1.28498e-20, 
    0, 7.709882e-21, -1.027984e-20, -1.541976e-20, -2.569961e-21, 
    1.027984e-20, 1.28498e-20, -5.139921e-21, 5.139921e-21, -1.003089e-36, 
    -1.003089e-36, -7.709882e-21, 7.709882e-21, -2.569961e-21, 1.28498e-20, 
    0, 2.569961e-21, -3.083953e-20, -5.139921e-21, -7.709882e-21, 
    2.569961e-21, 7.709882e-21, 5.139921e-21, 0, 2.569961e-21, -2.569961e-20, 
    5.139921e-21, 2.569961e-21, -1.003089e-36, -2.569961e-21, 2.569961e-21, 
    1.541976e-20, 1.027984e-20, -1.027984e-20, -5.139921e-21, 7.709882e-21, 
    -7.709882e-21, 5.139921e-21, 5.139921e-21, -2.569961e-21, -1.003089e-36, 
    0, -2.569961e-21, -2.569961e-21, 1.027984e-20, 2.569961e-21, 
    1.003089e-36, -2.569961e-21, 5.139921e-21, -2.569961e-21, 1.541976e-20, 
    1.027984e-20, -5.139921e-21, 2.569961e-21, 1.003089e-36, 5.139921e-21, 
    -5.139921e-21,
  5.139921e-21, 1.027984e-20, 1.027984e-20, 5.139921e-21, -1.28498e-20, 
    -1.541976e-20, -1.003089e-36, -2.569961e-21, -1.003089e-36, 1.541976e-20, 
    7.709882e-21, 1.003089e-36, 1.541976e-20, 7.709882e-21, 1.003089e-36, 
    1.28498e-20, 7.709882e-21, 5.139921e-21, 2.569961e-21, 7.709882e-21, 
    -1.003089e-36, -1.798972e-20, -1.003089e-36, 1.541976e-20, -5.139921e-21, 
    -1.798972e-20, -1.027984e-20, -1.003089e-36, -1.003089e-36, 
    -5.139921e-21, 0, 1.28498e-20, -2.569961e-21, 7.709882e-21, 5.139921e-21, 
    -5.139921e-21, 2.569961e-21, -1.027984e-20, -1.027984e-20, 2.569961e-21, 
    -2.569961e-21, -5.139921e-21, -1.541976e-20, -1.003089e-36, 
    -2.569961e-21, -5.139921e-21, 1.28498e-20, -2.569961e-20, -1.28498e-20, 
    1.027984e-20, -5.139921e-21, -1.541976e-20, -5.139921e-21, 7.709882e-21, 
    -1.027984e-20, 1.003089e-36, 2.569961e-21, 1.541976e-20, 0, 
    -7.709882e-21, 2.569961e-21, -1.798972e-20, 5.139921e-21, -7.709882e-21, 
    1.027984e-20, -2.569961e-21, 1.027984e-20, -2.569961e-21, -5.139921e-21, 
    2.055969e-20, 5.139921e-21, -1.28498e-20, 1.28498e-20, 1.541976e-20, 
    1.003089e-36, -2.569961e-21, -5.139921e-21, -7.709882e-21, 7.709882e-21, 
    -1.027984e-20, -2.055969e-20, -1.28498e-20, 1.003089e-36, 5.139921e-21, 
    1.541976e-20, 1.027984e-20, 7.709882e-21, -7.709882e-21, 5.139921e-21, 
    -7.709882e-21, -1.28498e-20, 7.709882e-21, 5.139921e-21, -7.709882e-21, 
    -7.709882e-21, -2.826957e-20, 1.027984e-20, 0, -5.139921e-21, 
    -1.027984e-20, 7.709882e-21, 2.569961e-21, -1.28498e-20, 1.798972e-20, 
    -1.798972e-20, -2.569961e-21, 1.027984e-20, 2.569961e-21, 2.569961e-21, 
    -1.541976e-20, -2.312965e-20, -1.003089e-36, 5.139921e-21, 5.139921e-21, 
    -2.569961e-21, 2.569961e-21, -2.569961e-21, 2.569961e-21, -7.709882e-21, 
    1.541976e-20, -1.798972e-20, -2.569961e-21, 2.055969e-20, 1.003089e-36, 
    2.569961e-21, -2.055969e-20, -1.003089e-36, -1.027984e-20, 1.541976e-20, 
    1.027984e-20, -5.139921e-21, 2.569961e-21, -7.709882e-21, -1.541976e-20, 
    2.569961e-21, -5.139921e-21, -1.798972e-20, -1.798972e-20, 2.569961e-21, 
    -2.569961e-21, 1.541976e-20, -2.569961e-21, -7.709882e-21, 1.541976e-20, 
    -2.569961e-21, 1.541976e-20, -1.541976e-20, -5.139921e-21, 5.139921e-21, 
    -2.569961e-21, 7.709882e-21, -1.28498e-20, 2.569961e-21, -7.709882e-21, 
    -2.569961e-21, -1.798972e-20, -7.709882e-21, 7.709882e-21, 1.027984e-20, 
    -2.312965e-20, 1.798972e-20, -2.055969e-20, -1.541976e-20, 2.569961e-21, 
    2.826957e-20, -1.003089e-36, 5.139921e-21, -1.027984e-20, 5.139921e-21, 
    -7.709882e-21, -2.055969e-20, -5.139921e-21, 7.709882e-21, 1.027984e-20, 
    -1.28498e-20, 0, -5.139921e-21, 1.027984e-20, -2.569961e-21, 
    7.709882e-21, 7.709882e-21, 2.569961e-21, -2.055969e-20, 2.569961e-21, 
    -1.28498e-20, -1.28498e-20, -5.139921e-21, -1.28498e-20, 1.027984e-20, 
    -1.027984e-20, 1.027984e-20, 1.28498e-20, 2.569961e-21, -7.709882e-21, 
    -5.139921e-21, 7.709882e-21, 1.28498e-20, 1.027984e-20, 1.541976e-20, 
    1.027984e-20, 7.709882e-21, -1.798972e-20, -1.003089e-36, 5.139921e-21, 
    1.541976e-20, 2.569961e-21, 5.139921e-21, -2.569961e-21, 1.541976e-20, 
    -7.709882e-21, -1.003089e-36, 2.569961e-21, 1.28498e-20, 2.569961e-20, 
    -7.709882e-21, 5.139921e-21, 2.569961e-21, 1.798972e-20, 2.569961e-21, 
    5.139921e-21, 1.027984e-20, -5.139921e-21, -1.28498e-20, -1.541976e-20, 
    -5.139921e-21, 2.569961e-20, 1.541976e-20, 7.709882e-21, -5.139921e-21, 
    1.027984e-20, 7.709882e-21, -1.003089e-36, -5.139921e-21, -2.569961e-21, 
    -5.139921e-21, -2.569961e-21, 5.139921e-21, -1.027984e-20, -2.569961e-21, 
    -5.139921e-21, 2.569961e-21, -2.569961e-21, 1.28498e-20, 7.709882e-21, 
    -5.139921e-21, 7.709882e-21, 7.709882e-21, -1.027984e-20, -1.003089e-36, 
    -1.28498e-20, 1.003089e-36, 2.569961e-20, 2.569961e-21, -5.139921e-21, 
    5.139921e-21, -2.055969e-20, 1.541976e-20, 2.569961e-21, 2.569961e-21, 
    5.139921e-21, -2.569961e-21, 1.027984e-20, -5.139921e-21, -1.027984e-20, 
    7.709882e-21, 1.28498e-20, -1.003089e-36, 2.569961e-21, -1.28498e-20, 
    -1.027984e-20, -2.569961e-21, 5.139921e-21, -1.027984e-20, 7.709882e-21, 
    2.569961e-21, 1.541976e-20, -1.541976e-20, 5.139921e-21, -2.569961e-21, 
    -7.709882e-21, -7.709882e-21, -1.003089e-36, -1.003089e-36, 7.709882e-21, 
    -1.027984e-20, 2.055969e-20, 2.312965e-20, -1.003089e-36, 1.003089e-36, 
    0, 7.709882e-21, 2.569961e-21, 2.569961e-21, 1.541976e-20, -2.569961e-21, 
    2.569961e-21, 7.709882e-21, -1.28498e-20, -5.139921e-21, 5.139921e-21, 
    -2.569961e-21, 7.709882e-21, 5.139921e-21, -1.027984e-20, 5.139921e-21, 
    -1.541976e-20, -5.139921e-21, -1.798972e-20, -1.28498e-20, 7.709882e-21, 
    1.027984e-20, 7.709882e-21, -2.569961e-21, 1.027984e-20, -1.027984e-20, 
    2.569961e-21, 7.709882e-21, 1.003089e-36, 2.569961e-21, -2.569961e-21, 
    -1.003089e-36, 2.569961e-21, -2.312965e-20, -2.569961e-21, 2.569961e-21, 
    2.312965e-20, -2.569961e-21, -5.139921e-21, -1.28498e-20, 1.027984e-20, 
    1.541976e-20, 2.569961e-21, 2.569961e-21, 0, -1.28498e-20, 2.055969e-20, 
    -1.541976e-20, 5.139921e-21,
  6.259378e-29, 6.259384e-29, 6.259383e-29, 6.259388e-29, 6.259385e-29, 
    6.259388e-29, 6.259379e-29, 6.259384e-29, 6.259381e-29, 6.259378e-29, 
    6.259398e-29, 6.259388e-29, 6.259407e-29, 6.259401e-29, 6.259417e-29, 
    6.259407e-29, 6.259419e-29, 6.259416e-29, 6.259423e-29, 6.259421e-29, 
    6.25943e-29, 6.259424e-29, 6.259435e-29, 6.259429e-29, 6.25943e-29, 
    6.259424e-29, 6.25939e-29, 6.259396e-29, 6.25939e-29, 6.25939e-29, 
    6.25939e-29, 6.259385e-29, 6.259382e-29, 6.259377e-29, 6.259378e-29, 
    6.259382e-29, 6.259391e-29, 6.259388e-29, 6.259395e-29, 6.259395e-29, 
    6.259404e-29, 6.2594e-29, 6.259414e-29, 6.25941e-29, 6.259422e-29, 
    6.259419e-29, 6.259421e-29, 6.25942e-29, 6.259421e-29, 6.259417e-29, 
    6.259419e-29, 6.259415e-29, 6.259401e-29, 6.259405e-29, 6.259392e-29, 
    6.259384e-29, 6.259379e-29, 6.259376e-29, 6.259376e-29, 6.259377e-29, 
    6.259382e-29, 6.259387e-29, 6.25939e-29, 6.259393e-29, 6.259395e-29, 
    6.259402e-29, 6.259406e-29, 6.259414e-29, 6.259413e-29, 6.259416e-29, 
    6.259418e-29, 6.259422e-29, 6.259422e-29, 6.259423e-29, 6.259416e-29, 
    6.259421e-29, 6.259412e-29, 6.259414e-29, 6.259396e-29, 6.259388e-29, 
    6.259385e-29, 6.259383e-29, 6.259376e-29, 6.259381e-29, 6.259379e-29, 
    6.259384e-29, 6.259386e-29, 6.259385e-29, 6.259393e-29, 6.25939e-29, 
    6.259407e-29, 6.259399e-29, 6.259418e-29, 6.259413e-29, 6.259419e-29, 
    6.259416e-29, 6.259421e-29, 6.259417e-29, 6.259424e-29, 6.259426e-29, 
    6.259425e-29, 6.259429e-29, 6.259416e-29, 6.259421e-29, 6.259385e-29, 
    6.259385e-29, 6.259386e-29, 6.259381e-29, 6.259381e-29, 6.259377e-29, 
    6.259381e-29, 6.259382e-29, 6.259386e-29, 6.259388e-29, 6.259391e-29, 
    6.259396e-29, 6.259401e-29, 6.259408e-29, 6.259414e-29, 6.259417e-29, 
    6.259415e-29, 6.259417e-29, 6.259415e-29, 6.259414e-29, 6.259425e-29, 
    6.259419e-29, 6.259428e-29, 6.259428e-29, 6.259423e-29, 6.259428e-29, 
    6.259385e-29, 6.259384e-29, 6.259379e-29, 6.259383e-29, 6.259377e-29, 
    6.25938e-29, 6.259382e-29, 6.25939e-29, 6.259391e-29, 6.259393e-29, 
    6.259396e-29, 6.2594e-29, 6.259407e-29, 6.259413e-29, 6.259419e-29, 
    6.259418e-29, 6.259418e-29, 6.259419e-29, 6.259416e-29, 6.25942e-29, 
    6.25942e-29, 6.259419e-29, 6.259428e-29, 6.259425e-29, 6.259428e-29, 
    6.259426e-29, 6.259384e-29, 6.259386e-29, 6.259385e-29, 6.259387e-29, 
    6.259386e-29, 6.259393e-29, 6.259394e-29, 6.259404e-29, 6.2594e-29, 
    6.259406e-29, 6.259401e-29, 6.259402e-29, 6.259406e-29, 6.259401e-29, 
    6.259413e-29, 6.259405e-29, 6.259419e-29, 6.259411e-29, 6.25942e-29, 
    6.259419e-29, 6.259421e-29, 6.259423e-29, 6.259426e-29, 6.259431e-29, 
    6.25943e-29, 6.259434e-29, 6.25939e-29, 6.259392e-29, 6.259392e-29, 
    6.259394e-29, 6.259397e-29, 6.259401e-29, 6.259408e-29, 6.259406e-29, 
    6.259411e-29, 6.259412e-29, 6.259404e-29, 6.259409e-29, 6.259394e-29, 
    6.259396e-29, 6.259395e-29, 6.25939e-29, 6.259407e-29, 6.259398e-29, 
    6.259414e-29, 6.259409e-29, 6.259423e-29, 6.259416e-29, 6.259429e-29, 
    6.259435e-29, 6.25944e-29, 6.259447e-29, 6.259393e-29, 6.259391e-29, 
    6.259395e-29, 6.259399e-29, 6.259404e-29, 6.25941e-29, 6.25941e-29, 
    6.259411e-29, 6.259414e-29, 6.259416e-29, 6.259411e-29, 6.259417e-29, 
    6.259397e-29, 6.259407e-29, 6.259391e-29, 6.259396e-29, 6.259399e-29, 
    6.259398e-29, 6.259405e-29, 6.259407e-29, 6.259415e-29, 6.259411e-29, 
    6.259434e-29, 6.259423e-29, 6.259452e-29, 6.259444e-29, 6.259391e-29, 
    6.259393e-29, 6.259402e-29, 6.259398e-29, 6.25941e-29, 6.259413e-29, 
    6.259415e-29, 6.259418e-29, 6.259419e-29, 6.25942e-29, 6.259417e-29, 
    6.25942e-29, 6.25941e-29, 6.259414e-29, 6.259401e-29, 6.259404e-29, 
    6.259403e-29, 6.259401e-29, 6.259406e-29, 6.259411e-29, 6.259411e-29, 
    6.259413e-29, 6.259418e-29, 6.25941e-29, 6.259435e-29, 6.259419e-29, 
    6.259396e-29, 6.259401e-29, 6.259402e-29, 6.2594e-29, 6.259413e-29, 
    6.259408e-29, 6.25942e-29, 6.259417e-29, 6.259422e-29, 6.259419e-29, 
    6.259419e-29, 6.259416e-29, 6.259413e-29, 6.259408e-29, 6.259404e-29, 
    6.2594e-29, 6.259401e-29, 6.259405e-29, 6.259412e-29, 6.259419e-29, 
    6.259417e-29, 6.259422e-29, 6.259409e-29, 6.259414e-29, 6.259412e-29, 
    6.259417e-29, 6.259406e-29, 6.259416e-29, 6.259403e-29, 6.259404e-29, 
    6.259408e-29, 6.259414e-29, 6.259416e-29, 6.259418e-29, 6.259417e-29, 
    6.259412e-29, 6.259411e-29, 6.259408e-29, 6.259407e-29, 6.259404e-29, 
    6.259402e-29, 6.259404e-29, 6.259406e-29, 6.259412e-29, 6.259417e-29, 
    6.259423e-29, 6.259425e-29, 6.259431e-29, 6.259426e-29, 6.259435e-29, 
    6.259427e-29, 6.259441e-29, 6.259416e-29, 6.259427e-29, 6.259408e-29, 
    6.25941e-29, 6.259414e-29, 6.259422e-29, 6.259417e-29, 6.259423e-29, 
    6.259411e-29, 6.259405e-29, 6.259404e-29, 6.259401e-29, 6.259404e-29, 
    6.259403e-29, 6.259406e-29, 6.259405e-29, 6.259412e-29, 6.259408e-29, 
    6.259419e-29, 6.259423e-29, 6.259434e-29, 6.259441e-29, 6.259447e-29, 
    6.25945e-29, 6.259452e-29, 6.259452e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2N_TO_SOIL1N =
  2.136685e-10, 2.146114e-10, 2.144281e-10, 2.151886e-10, 2.147668e-10, 
    2.152648e-10, 2.138597e-10, 2.146488e-10, 2.14145e-10, 2.137534e-10, 
    2.166646e-10, 2.152226e-10, 2.181628e-10, 2.17243e-10, 2.195538e-10, 
    2.180197e-10, 2.198632e-10, 2.195096e-10, 2.205739e-10, 2.20269e-10, 
    2.216303e-10, 2.207147e-10, 2.223361e-10, 2.214117e-10, 2.215562e-10, 
    2.206844e-10, 2.155128e-10, 2.164851e-10, 2.154552e-10, 2.155938e-10, 
    2.155316e-10, 2.147755e-10, 2.143944e-10, 2.135964e-10, 2.137413e-10, 
    2.143274e-10, 2.156562e-10, 2.152051e-10, 2.16342e-10, 2.163163e-10, 
    2.17582e-10, 2.170114e-10, 2.191389e-10, 2.185342e-10, 2.202818e-10, 
    2.198422e-10, 2.202611e-10, 2.201341e-10, 2.202628e-10, 2.196182e-10, 
    2.198943e-10, 2.193272e-10, 2.171182e-10, 2.177674e-10, 2.158314e-10, 
    2.146673e-10, 2.138943e-10, 2.133457e-10, 2.134233e-10, 2.135711e-10, 
    2.143308e-10, 2.150452e-10, 2.155896e-10, 2.159538e-10, 2.163126e-10, 
    2.173987e-10, 2.179737e-10, 2.192612e-10, 2.190289e-10, 2.194225e-10, 
    2.197985e-10, 2.204299e-10, 2.20326e-10, 2.206041e-10, 2.194121e-10, 
    2.202043e-10, 2.188965e-10, 2.192542e-10, 2.1641e-10, 2.153268e-10, 
    2.148663e-10, 2.144633e-10, 2.134829e-10, 2.1416e-10, 2.13893e-10, 
    2.145281e-10, 2.149316e-10, 2.14732e-10, 2.159638e-10, 2.154849e-10, 
    2.180078e-10, 2.169211e-10, 2.197546e-10, 2.190765e-10, 2.199172e-10, 
    2.194882e-10, 2.202232e-10, 2.195617e-10, 2.207076e-10, 2.209571e-10, 
    2.207866e-10, 2.214417e-10, 2.195251e-10, 2.202611e-10, 2.147264e-10, 
    2.14759e-10, 2.149106e-10, 2.14244e-10, 2.142033e-10, 2.135925e-10, 
    2.14136e-10, 2.143674e-10, 2.14955e-10, 2.153025e-10, 2.156329e-10, 
    2.163594e-10, 2.171707e-10, 2.183053e-10, 2.191205e-10, 2.19667e-10, 
    2.193319e-10, 2.196277e-10, 2.19297e-10, 2.19142e-10, 2.208636e-10, 
    2.198969e-10, 2.213475e-10, 2.212672e-10, 2.206107e-10, 2.212762e-10, 
    2.147818e-10, 2.145945e-10, 2.139442e-10, 2.144531e-10, 2.13526e-10, 
    2.140449e-10, 2.143433e-10, 2.154948e-10, 2.157479e-10, 2.159825e-10, 
    2.164459e-10, 2.170406e-10, 2.180838e-10, 2.189916e-10, 2.198204e-10, 
    2.197597e-10, 2.197811e-10, 2.199662e-10, 2.195076e-10, 2.200415e-10, 
    2.201311e-10, 2.198968e-10, 2.212565e-10, 2.20868e-10, 2.212655e-10, 
    2.210126e-10, 2.146554e-10, 2.149706e-10, 2.148003e-10, 2.151205e-10, 
    2.148949e-10, 2.158981e-10, 2.161989e-10, 2.176065e-10, 2.170289e-10, 
    2.179482e-10, 2.171223e-10, 2.172686e-10, 2.179782e-10, 2.171669e-10, 
    2.189415e-10, 2.177383e-10, 2.199734e-10, 2.187717e-10, 2.200487e-10, 
    2.198168e-10, 2.202007e-10, 2.205446e-10, 2.209772e-10, 2.217754e-10, 
    2.215905e-10, 2.222581e-10, 2.154404e-10, 2.158492e-10, 2.158133e-10, 
    2.162411e-10, 2.165575e-10, 2.172433e-10, 2.183433e-10, 2.179297e-10, 
    2.186891e-10, 2.188416e-10, 2.176878e-10, 2.183961e-10, 2.161228e-10, 
    2.1649e-10, 2.162714e-10, 2.154727e-10, 2.180249e-10, 2.16715e-10, 
    2.19134e-10, 2.184243e-10, 2.204955e-10, 2.194654e-10, 2.214888e-10, 
    2.223537e-10, 2.23168e-10, 2.241194e-10, 2.160723e-10, 2.157946e-10, 
    2.16292e-10, 2.169801e-10, 2.176186e-10, 2.184676e-10, 2.185545e-10, 
    2.187135e-10, 2.191255e-10, 2.194719e-10, 2.187638e-10, 2.195587e-10, 
    2.165752e-10, 2.181387e-10, 2.156895e-10, 2.164269e-10, 2.169395e-10, 
    2.167147e-10, 2.178824e-10, 2.181576e-10, 2.19276e-10, 2.186979e-10, 
    2.221402e-10, 2.206171e-10, 2.24844e-10, 2.236626e-10, 2.156975e-10, 
    2.160714e-10, 2.173726e-10, 2.167535e-10, 2.185243e-10, 2.189602e-10, 
    2.193145e-10, 2.197675e-10, 2.198164e-10, 2.200848e-10, 2.19645e-10, 
    2.200675e-10, 2.184694e-10, 2.191835e-10, 2.172239e-10, 2.177008e-10, 
    2.174815e-10, 2.172408e-10, 2.179836e-10, 2.187749e-10, 2.187919e-10, 
    2.190456e-10, 2.197605e-10, 2.185315e-10, 2.223367e-10, 2.199865e-10, 
    2.164791e-10, 2.171992e-10, 2.173021e-10, 2.170232e-10, 2.189165e-10, 
    2.182304e-10, 2.200783e-10, 2.195789e-10, 2.203972e-10, 2.199905e-10, 
    2.199307e-10, 2.194085e-10, 2.190833e-10, 2.182619e-10, 2.175936e-10, 
    2.170636e-10, 2.171869e-10, 2.17769e-10, 2.188233e-10, 2.198208e-10, 
    2.196023e-10, 2.20335e-10, 2.183959e-10, 2.192089e-10, 2.188947e-10, 
    2.197141e-10, 2.179187e-10, 2.194474e-10, 2.175279e-10, 2.176962e-10, 
    2.182168e-10, 2.19264e-10, 2.194958e-10, 2.197432e-10, 2.195906e-10, 
    2.188501e-10, 2.187288e-10, 2.182042e-10, 2.180593e-10, 2.176596e-10, 
    2.173286e-10, 2.17631e-10, 2.179485e-10, 2.188504e-10, 2.196632e-10, 
    2.205495e-10, 2.207664e-10, 2.218018e-10, 2.209588e-10, 2.223498e-10, 
    2.211671e-10, 2.232145e-10, 2.195361e-10, 2.211324e-10, 2.182405e-10, 
    2.185521e-10, 2.191155e-10, 2.20408e-10, 2.197103e-10, 2.205263e-10, 
    2.187241e-10, 2.17789e-10, 2.175472e-10, 2.170959e-10, 2.175575e-10, 
    2.175199e-10, 2.179617e-10, 2.178197e-10, 2.188804e-10, 2.183106e-10, 
    2.199292e-10, 2.205199e-10, 2.221881e-10, 2.232109e-10, 2.242521e-10, 
    2.247117e-10, 2.248517e-10, 2.249102e-10 ;

 SOIL2N_TO_SOIL3N =
  1.526203e-11, 1.532939e-11, 1.531629e-11, 1.537062e-11, 1.534048e-11, 
    1.537605e-11, 1.527569e-11, 1.533206e-11, 1.529608e-11, 1.52681e-11, 
    1.547604e-11, 1.537304e-11, 1.558306e-11, 1.551736e-11, 1.568242e-11, 
    1.557283e-11, 1.570451e-11, 1.567926e-11, 1.575528e-11, 1.57335e-11, 
    1.583074e-11, 1.576533e-11, 1.588115e-11, 1.581512e-11, 1.582545e-11, 
    1.576318e-11, 1.539377e-11, 1.546322e-11, 1.538966e-11, 1.539956e-11, 
    1.539512e-11, 1.534111e-11, 1.531388e-11, 1.525689e-11, 1.526724e-11, 
    1.53091e-11, 1.540401e-11, 1.53718e-11, 1.5453e-11, 1.545117e-11, 
    1.554157e-11, 1.550081e-11, 1.565278e-11, 1.560959e-11, 1.573441e-11, 
    1.570302e-11, 1.573294e-11, 1.572386e-11, 1.573305e-11, 1.568701e-11, 
    1.570674e-11, 1.566623e-11, 1.550845e-11, 1.555481e-11, 1.541653e-11, 
    1.533338e-11, 1.527816e-11, 1.523898e-11, 1.524452e-11, 1.525508e-11, 
    1.530935e-11, 1.536037e-11, 1.539926e-11, 1.542527e-11, 1.54509e-11, 
    1.552848e-11, 1.556955e-11, 1.566151e-11, 1.564492e-11, 1.567303e-11, 
    1.569989e-11, 1.574499e-11, 1.573757e-11, 1.575744e-11, 1.567229e-11, 
    1.572888e-11, 1.563547e-11, 1.566101e-11, 1.545786e-11, 1.538049e-11, 
    1.534759e-11, 1.531881e-11, 1.524878e-11, 1.529714e-11, 1.527807e-11, 
    1.532343e-11, 1.535226e-11, 1.5338e-11, 1.542598e-11, 1.539178e-11, 
    1.557199e-11, 1.549436e-11, 1.569676e-11, 1.564832e-11, 1.570837e-11, 
    1.567773e-11, 1.573023e-11, 1.568298e-11, 1.576483e-11, 1.578265e-11, 
    1.577047e-11, 1.581726e-11, 1.568036e-11, 1.573293e-11, 1.53376e-11, 
    1.533993e-11, 1.535076e-11, 1.530314e-11, 1.530023e-11, 1.525661e-11, 
    1.529543e-11, 1.531196e-11, 1.535393e-11, 1.537875e-11, 1.540235e-11, 
    1.545424e-11, 1.551219e-11, 1.559324e-11, 1.565146e-11, 1.56905e-11, 
    1.566656e-11, 1.568769e-11, 1.566407e-11, 1.5653e-11, 1.577597e-11, 
    1.570692e-11, 1.581053e-11, 1.58048e-11, 1.575791e-11, 1.580545e-11, 
    1.534156e-11, 1.532818e-11, 1.528173e-11, 1.531808e-11, 1.525185e-11, 
    1.528892e-11, 1.531024e-11, 1.539249e-11, 1.541057e-11, 1.542732e-11, 
    1.546042e-11, 1.55029e-11, 1.557742e-11, 1.564226e-11, 1.570146e-11, 
    1.569712e-11, 1.569865e-11, 1.571187e-11, 1.567911e-11, 1.571725e-11, 
    1.572365e-11, 1.570691e-11, 1.580403e-11, 1.577629e-11, 1.580468e-11, 
    1.578661e-11, 1.533253e-11, 1.535504e-11, 1.534288e-11, 1.536575e-11, 
    1.534963e-11, 1.542129e-11, 1.544278e-11, 1.554332e-11, 1.550206e-11, 
    1.556773e-11, 1.550873e-11, 1.551918e-11, 1.556987e-11, 1.551192e-11, 
    1.563868e-11, 1.555274e-11, 1.571238e-11, 1.562655e-11, 1.571776e-11, 
    1.57012e-11, 1.572862e-11, 1.575318e-11, 1.578408e-11, 1.58411e-11, 
    1.582789e-11, 1.587558e-11, 1.53886e-11, 1.54178e-11, 1.541523e-11, 
    1.544579e-11, 1.546839e-11, 1.551738e-11, 1.559595e-11, 1.55664e-11, 
    1.562065e-11, 1.563154e-11, 1.554913e-11, 1.559972e-11, 1.543734e-11, 
    1.546357e-11, 1.544796e-11, 1.53909e-11, 1.557321e-11, 1.547965e-11, 
    1.565243e-11, 1.560174e-11, 1.574968e-11, 1.56761e-11, 1.582063e-11, 
    1.588241e-11, 1.594057e-11, 1.600853e-11, 1.543374e-11, 1.54139e-11, 
    1.544943e-11, 1.549858e-11, 1.554419e-11, 1.560483e-11, 1.561103e-11, 
    1.562239e-11, 1.565182e-11, 1.567656e-11, 1.562598e-11, 1.568277e-11, 
    1.546966e-11, 1.558133e-11, 1.54064e-11, 1.545907e-11, 1.549568e-11, 
    1.547962e-11, 1.556303e-11, 1.558269e-11, 1.566257e-11, 1.562128e-11, 
    1.586716e-11, 1.575837e-11, 1.606029e-11, 1.59759e-11, 1.540697e-11, 
    1.543367e-11, 1.552662e-11, 1.548239e-11, 1.560888e-11, 1.564001e-11, 
    1.566532e-11, 1.569768e-11, 1.570117e-11, 1.572035e-11, 1.568893e-11, 
    1.57191e-11, 1.560496e-11, 1.565597e-11, 1.5516e-11, 1.555006e-11, 
    1.553439e-11, 1.55172e-11, 1.557026e-11, 1.562678e-11, 1.562799e-11, 
    1.564611e-11, 1.569718e-11, 1.560939e-11, 1.588119e-11, 1.571332e-11, 
    1.546279e-11, 1.551423e-11, 1.552158e-11, 1.550166e-11, 1.563689e-11, 
    1.558789e-11, 1.571988e-11, 1.568421e-11, 1.574266e-11, 1.571361e-11, 
    1.570934e-11, 1.567203e-11, 1.564881e-11, 1.559013e-11, 1.55424e-11, 
    1.550455e-11, 1.551335e-11, 1.555493e-11, 1.563024e-11, 1.570149e-11, 
    1.568588e-11, 1.573821e-11, 1.559971e-11, 1.565778e-11, 1.563533e-11, 
    1.569387e-11, 1.556562e-11, 1.567482e-11, 1.553771e-11, 1.554973e-11, 
    1.558692e-11, 1.566172e-11, 1.567827e-11, 1.569594e-11, 1.568504e-11, 
    1.563215e-11, 1.562349e-11, 1.558601e-11, 1.557566e-11, 1.554711e-11, 
    1.552347e-11, 1.554507e-11, 1.556775e-11, 1.563217e-11, 1.569023e-11, 
    1.575353e-11, 1.576903e-11, 1.584298e-11, 1.578277e-11, 1.588213e-11, 
    1.579765e-11, 1.594389e-11, 1.568115e-11, 1.579517e-11, 1.558861e-11, 
    1.561086e-11, 1.565111e-11, 1.574343e-11, 1.569359e-11, 1.575188e-11, 
    1.562315e-11, 1.555636e-11, 1.553908e-11, 1.550685e-11, 1.553982e-11, 
    1.553714e-11, 1.556869e-11, 1.555855e-11, 1.563431e-11, 1.559362e-11, 
    1.570923e-11, 1.575142e-11, 1.587058e-11, 1.594363e-11, 1.6018e-11, 
    1.605084e-11, 1.606083e-11, 1.606501e-11 ;

 SOIL2N_vr =
  1.818715, 1.818717, 1.818716, 1.818717, 1.818717, 1.818718, 1.818715, 
    1.818717, 1.818716, 1.818715, 1.81872, 1.818717, 1.818722, 1.818721, 
    1.818724, 1.818722, 1.818725, 1.818724, 1.818726, 1.818725, 1.818727, 
    1.818726, 1.818729, 1.818727, 1.818727, 1.818726, 1.818718, 1.81872, 
    1.818718, 1.818718, 1.818718, 1.818717, 1.818716, 1.818715, 1.818715, 
    1.818716, 1.818718, 1.818717, 1.818719, 1.818719, 1.818721, 1.81872, 
    1.818724, 1.818723, 1.818725, 1.818725, 1.818725, 1.818725, 1.818725, 
    1.818724, 1.818725, 1.818724, 1.81872, 1.818721, 1.818718, 1.818717, 
    1.818715, 1.818715, 1.818715, 1.818715, 1.818716, 1.818717, 1.818718, 
    1.818719, 1.818719, 1.818721, 1.818722, 1.818724, 1.818723, 1.818724, 
    1.818725, 1.818726, 1.818725, 1.818726, 1.818724, 1.818725, 1.818723, 
    1.818724, 1.818719, 1.818718, 1.818717, 1.818716, 1.818715, 1.818716, 
    1.818715, 1.818716, 1.818717, 1.818717, 1.818719, 1.818718, 1.818722, 
    1.81872, 1.818725, 1.818723, 1.818725, 1.818724, 1.818725, 1.818724, 
    1.818726, 1.818726, 1.818726, 1.818727, 1.818724, 1.818725, 1.818717, 
    1.818717, 1.818717, 1.818716, 1.818716, 1.818715, 1.818716, 1.818716, 
    1.818717, 1.818718, 1.818718, 1.818719, 1.818721, 1.818722, 1.818724, 
    1.818724, 1.818724, 1.818724, 1.818724, 1.818724, 1.818726, 1.818725, 
    1.818727, 1.818727, 1.818726, 1.818727, 1.818717, 1.818717, 1.818715, 
    1.818716, 1.818715, 1.818716, 1.818716, 1.818718, 1.818718, 1.818719, 
    1.818719, 1.81872, 1.818722, 1.818723, 1.818725, 1.818725, 1.818725, 
    1.818725, 1.818724, 1.818725, 1.818725, 1.818725, 1.818727, 1.818726, 
    1.818727, 1.818726, 1.818717, 1.818717, 1.818717, 1.818717, 1.818717, 
    1.818719, 1.818719, 1.818721, 1.81872, 1.818722, 1.81872, 1.818721, 
    1.818722, 1.81872, 1.818723, 1.818721, 1.818725, 1.818723, 1.818725, 
    1.818725, 1.818725, 1.818726, 1.818726, 1.818728, 1.818727, 1.818728, 
    1.818718, 1.818718, 1.818718, 1.818719, 1.81872, 1.818721, 1.818722, 
    1.818722, 1.818723, 1.818723, 1.818721, 1.818722, 1.818719, 1.81872, 
    1.818719, 1.818718, 1.818722, 1.81872, 1.818724, 1.818722, 1.818726, 
    1.818724, 1.818727, 1.818729, 1.81873, 1.818731, 1.818719, 1.818718, 
    1.818719, 1.81872, 1.818721, 1.818722, 1.818723, 1.818723, 1.818724, 
    1.818724, 1.818723, 1.818724, 1.81872, 1.818722, 1.818718, 1.818719, 
    1.81872, 1.81872, 1.818722, 1.818722, 1.818724, 1.818723, 1.818728, 
    1.818726, 1.818732, 1.818731, 1.818718, 1.818719, 1.818721, 1.81872, 
    1.818723, 1.818723, 1.818724, 1.818725, 1.818725, 1.818725, 1.818724, 
    1.818725, 1.818722, 1.818724, 1.818721, 1.818721, 1.818721, 1.818721, 
    1.818722, 1.818723, 1.818723, 1.818723, 1.818725, 1.818723, 1.818729, 
    1.818725, 1.81872, 1.818721, 1.818721, 1.81872, 1.818723, 1.818722, 
    1.818725, 1.818724, 1.818725, 1.818725, 1.818725, 1.818724, 1.818723, 
    1.818722, 1.818721, 1.81872, 1.818721, 1.818721, 1.818723, 1.818725, 
    1.818724, 1.818725, 1.818722, 1.818724, 1.818723, 1.818725, 1.818722, 
    1.818724, 1.818721, 1.818721, 1.818722, 1.818724, 1.818724, 1.818725, 
    1.818724, 1.818723, 1.818723, 1.818722, 1.818722, 1.818721, 1.818721, 
    1.818721, 1.818722, 1.818723, 1.818724, 1.818726, 1.818726, 1.818728, 
    1.818726, 1.818729, 1.818727, 1.81873, 1.818724, 1.818727, 1.818722, 
    1.818723, 1.818724, 1.818726, 1.818725, 1.818726, 1.818723, 1.818722, 
    1.818721, 1.81872, 1.818721, 1.818721, 1.818722, 1.818722, 1.818723, 
    1.818722, 1.818725, 1.818726, 1.818728, 1.81873, 1.818731, 1.818732, 
    1.818732, 1.818733,
  1.818667, 1.818669, 1.818668, 1.81867, 1.818669, 1.81867, 1.818667, 
    1.818669, 1.818668, 1.818667, 1.818673, 1.81867, 1.818676, 1.818674, 
    1.818678, 1.818676, 1.818679, 1.818678, 1.818681, 1.81868, 1.818683, 
    1.818681, 1.818684, 1.818682, 1.818682, 1.818681, 1.818671, 1.818673, 
    1.818671, 1.818671, 1.818671, 1.818669, 1.818668, 1.818667, 1.818667, 
    1.818668, 1.818671, 1.81867, 1.818672, 1.818672, 1.818675, 1.818674, 
    1.818678, 1.818676, 1.81868, 1.818679, 1.81868, 1.81868, 1.81868, 
    1.818679, 1.818679, 1.818678, 1.818674, 1.818675, 1.818671, 1.818669, 
    1.818668, 1.818666, 1.818667, 1.818667, 1.818668, 1.81867, 1.818671, 
    1.818671, 1.818672, 1.818674, 1.818675, 1.818678, 1.818677, 1.818678, 
    1.818679, 1.81868, 1.81868, 1.818681, 1.818678, 1.81868, 1.818677, 
    1.818678, 1.818672, 1.81867, 1.818669, 1.818669, 1.818667, 1.818668, 
    1.818668, 1.818669, 1.81867, 1.818669, 1.818671, 1.818671, 1.818676, 
    1.818673, 1.818679, 1.818678, 1.818679, 1.818678, 1.81868, 1.818678, 
    1.818681, 1.818681, 1.818681, 1.818682, 1.818678, 1.81868, 1.818669, 
    1.818669, 1.818669, 1.818668, 1.818668, 1.818667, 1.818668, 1.818668, 
    1.81867, 1.81867, 1.818671, 1.818672, 1.818674, 1.818676, 1.818678, 
    1.818679, 1.818678, 1.818679, 1.818678, 1.818678, 1.818681, 1.818679, 
    1.818682, 1.818682, 1.818681, 1.818682, 1.818669, 1.818669, 1.818668, 
    1.818669, 1.818667, 1.818668, 1.818668, 1.818671, 1.818671, 1.818672, 
    1.818672, 1.818674, 1.818676, 1.818677, 1.818679, 1.818679, 1.818679, 
    1.818679, 1.818678, 1.818679, 1.81868, 1.818679, 1.818682, 1.818681, 
    1.818682, 1.818681, 1.818669, 1.81867, 1.818669, 1.81867, 1.818669, 
    1.818671, 1.818672, 1.818675, 1.818674, 1.818675, 1.818674, 1.818674, 
    1.818675, 1.818674, 1.818677, 1.818675, 1.818679, 1.818677, 1.818679, 
    1.818679, 1.81868, 1.81868, 1.818681, 1.818683, 1.818682, 1.818684, 
    1.818671, 1.818671, 1.818671, 1.818672, 1.818673, 1.818674, 1.818676, 
    1.818675, 1.818677, 1.818677, 1.818675, 1.818676, 1.818672, 1.818673, 
    1.818672, 1.818671, 1.818676, 1.818673, 1.818678, 1.818676, 1.81868, 
    1.818678, 1.818682, 1.818684, 1.818686, 1.818687, 1.818672, 1.818671, 
    1.818672, 1.818673, 1.818675, 1.818676, 1.818677, 1.818677, 1.818678, 
    1.818678, 1.818677, 1.818678, 1.818673, 1.818676, 1.818671, 1.818672, 
    1.818673, 1.818673, 1.818675, 1.818676, 1.818678, 1.818677, 1.818684, 
    1.818681, 1.818689, 1.818686, 1.818671, 1.818672, 1.818674, 1.818673, 
    1.818676, 1.818677, 1.818678, 1.818679, 1.818679, 1.81868, 1.818679, 
    1.818679, 1.818676, 1.818678, 1.818674, 1.818675, 1.818674, 1.818674, 
    1.818675, 1.818677, 1.818677, 1.818678, 1.818679, 1.818676, 1.818684, 
    1.818679, 1.818673, 1.818674, 1.818674, 1.818674, 1.818677, 1.818676, 
    1.81868, 1.818678, 1.81868, 1.818679, 1.818679, 1.818678, 1.818678, 
    1.818676, 1.818675, 1.818674, 1.818674, 1.818675, 1.818677, 1.818679, 
    1.818679, 1.81868, 1.818676, 1.818678, 1.818677, 1.818679, 1.818675, 
    1.818678, 1.818675, 1.818675, 1.818676, 1.818678, 1.818678, 1.818679, 
    1.818679, 1.818677, 1.818677, 1.818676, 1.818676, 1.818675, 1.818674, 
    1.818675, 1.818675, 1.818677, 1.818679, 1.81868, 1.818681, 1.818683, 
    1.818681, 1.818684, 1.818682, 1.818686, 1.818678, 1.818682, 1.818676, 
    1.818677, 1.818678, 1.81868, 1.818679, 1.81868, 1.818677, 1.818675, 
    1.818675, 1.818674, 1.818675, 1.818675, 1.818675, 1.818675, 1.818677, 
    1.818676, 1.818679, 1.81868, 1.818684, 1.818686, 1.818688, 1.818689, 
    1.818689, 1.818689,
  1.818639, 1.818641, 1.818641, 1.818642, 1.818642, 1.818643, 1.81864, 
    1.818641, 1.81864, 1.818639, 1.818646, 1.818642, 1.818649, 1.818647, 
    1.818652, 1.818648, 1.818652, 1.818652, 1.818654, 1.818653, 1.818656, 
    1.818654, 1.818658, 1.818656, 1.818656, 1.818654, 1.818643, 1.818645, 
    1.818643, 1.818643, 1.818643, 1.818642, 1.818641, 1.818639, 1.818639, 
    1.818641, 1.818643, 1.818642, 1.818645, 1.818645, 1.818648, 1.818646, 
    1.818651, 1.81865, 1.818653, 1.818652, 1.818653, 1.818653, 1.818653, 
    1.818652, 1.818653, 1.818651, 1.818647, 1.818648, 1.818644, 1.818641, 
    1.81864, 1.818638, 1.818639, 1.818639, 1.818641, 1.818642, 1.818643, 
    1.818644, 1.818645, 1.818647, 1.818648, 1.818651, 1.818651, 1.818652, 
    1.818652, 1.818654, 1.818653, 1.818654, 1.818651, 1.818653, 1.81865, 
    1.818651, 1.818645, 1.818643, 1.818642, 1.818641, 1.818639, 1.81864, 
    1.81864, 1.818641, 1.818642, 1.818641, 1.818644, 1.818643, 1.818648, 
    1.818646, 1.818652, 1.818651, 1.818653, 1.818652, 1.818653, 1.818652, 
    1.818654, 1.818655, 1.818654, 1.818656, 1.818652, 1.818653, 1.818641, 
    1.818642, 1.818642, 1.81864, 1.81864, 1.818639, 1.81864, 1.818641, 
    1.818642, 1.818643, 1.818643, 1.818645, 1.818647, 1.818649, 1.818651, 
    1.818652, 1.818651, 1.818652, 1.818651, 1.818651, 1.818655, 1.818653, 
    1.818656, 1.818655, 1.818654, 1.818655, 1.818642, 1.818641, 1.81864, 
    1.818641, 1.818639, 1.81864, 1.818641, 1.818643, 1.818644, 1.818644, 
    1.818645, 1.818646, 1.818649, 1.818651, 1.818652, 1.818652, 1.818652, 
    1.818653, 1.818652, 1.818653, 1.818653, 1.818653, 1.818655, 1.818655, 
    1.818655, 1.818655, 1.818641, 1.818642, 1.818642, 1.818642, 1.818642, 
    1.818644, 1.818645, 1.818648, 1.818646, 1.818648, 1.818647, 1.818647, 
    1.818648, 1.818647, 1.81865, 1.818648, 1.818653, 1.81865, 1.818653, 
    1.818652, 1.818653, 1.818654, 1.818655, 1.818657, 1.818656, 1.818658, 
    1.818643, 1.818644, 1.818644, 1.818645, 1.818645, 1.818647, 1.818649, 
    1.818648, 1.81865, 1.81865, 1.818648, 1.818649, 1.818644, 1.818645, 
    1.818645, 1.818643, 1.818648, 1.818646, 1.818651, 1.818649, 1.818654, 
    1.818652, 1.818656, 1.818658, 1.81866, 1.818662, 1.818644, 1.818644, 
    1.818645, 1.818646, 1.818648, 1.818649, 1.81865, 1.81865, 1.818651, 
    1.818652, 1.81865, 1.818652, 1.818645, 1.818649, 1.818643, 1.818645, 
    1.818646, 1.818646, 1.818648, 1.818649, 1.818651, 1.81865, 1.818657, 
    1.818654, 1.818663, 1.818661, 1.818644, 1.818644, 1.818647, 1.818646, 
    1.81865, 1.81865, 1.818651, 1.818652, 1.818652, 1.818653, 1.818652, 
    1.818653, 1.818649, 1.818651, 1.818647, 1.818648, 1.818647, 1.818647, 
    1.818648, 1.81865, 1.81865, 1.818651, 1.818652, 1.81865, 1.818658, 
    1.818653, 1.818645, 1.818647, 1.818647, 1.818646, 1.81865, 1.818649, 
    1.818653, 1.818652, 1.818654, 1.818653, 1.818653, 1.818651, 1.818651, 
    1.818649, 1.818648, 1.818646, 1.818647, 1.818648, 1.81865, 1.818652, 
    1.818652, 1.818653, 1.818649, 1.818651, 1.81865, 1.818652, 1.818648, 
    1.818652, 1.818647, 1.818648, 1.818649, 1.818651, 1.818652, 1.818652, 
    1.818652, 1.81865, 1.81865, 1.818649, 1.818649, 1.818648, 1.818647, 
    1.818648, 1.818648, 1.81865, 1.818652, 1.818654, 1.818654, 1.818657, 
    1.818655, 1.818658, 1.818655, 1.81866, 1.818652, 1.818655, 1.818649, 
    1.81865, 1.818651, 1.818654, 1.818652, 1.818654, 1.81865, 1.818648, 
    1.818648, 1.818647, 1.818648, 1.818647, 1.818648, 1.818648, 1.81865, 
    1.818649, 1.818653, 1.818654, 1.818657, 1.81866, 1.818662, 1.818663, 
    1.818663, 1.818663,
  1.818617, 1.818619, 1.818619, 1.818621, 1.81862, 1.818621, 1.818618, 
    1.818619, 1.818618, 1.818618, 1.818624, 1.818621, 1.818627, 1.818625, 
    1.81863, 1.818627, 1.818631, 1.81863, 1.818632, 1.818632, 1.818635, 
    1.818633, 1.818636, 1.818634, 1.818635, 1.818633, 1.818621, 1.818624, 
    1.818621, 1.818622, 1.818622, 1.81862, 1.818619, 1.818617, 1.818618, 
    1.818619, 1.818622, 1.818621, 1.818623, 1.818623, 1.818626, 1.818625, 
    1.818629, 1.818628, 1.818632, 1.818631, 1.818632, 1.818632, 1.818632, 
    1.81863, 1.818631, 1.81863, 1.818625, 1.818626, 1.818622, 1.81862, 
    1.818618, 1.818617, 1.818617, 1.818617, 1.818619, 1.81862, 1.818622, 
    1.818622, 1.818623, 1.818626, 1.818627, 1.81863, 1.818629, 1.81863, 
    1.818631, 1.818632, 1.818632, 1.818633, 1.81863, 1.818632, 1.818629, 
    1.81863, 1.818623, 1.818621, 1.81862, 1.818619, 1.818617, 1.818618, 
    1.818618, 1.818619, 1.81862, 1.81862, 1.818622, 1.818621, 1.818627, 
    1.818624, 1.818631, 1.818629, 1.818631, 1.81863, 1.818632, 1.81863, 
    1.818633, 1.818633, 1.818633, 1.818634, 1.81863, 1.818632, 1.81862, 
    1.81862, 1.81862, 1.818619, 1.818619, 1.818617, 1.818618, 1.818619, 
    1.81862, 1.818621, 1.818622, 1.818623, 1.818625, 1.818628, 1.818629, 
    1.818631, 1.81863, 1.81863, 1.81863, 1.818629, 1.818633, 1.818631, 
    1.818634, 1.818634, 1.818633, 1.818634, 1.81862, 1.818619, 1.818618, 
    1.818619, 1.818617, 1.818618, 1.818619, 1.818621, 1.818622, 1.818622, 
    1.818623, 1.818625, 1.818627, 1.818629, 1.818631, 1.818631, 1.818631, 
    1.818631, 1.81863, 1.818631, 1.818632, 1.818631, 1.818634, 1.818633, 
    1.818634, 1.818633, 1.81862, 1.81862, 1.81862, 1.818621, 1.81862, 
    1.818622, 1.818623, 1.818626, 1.818625, 1.818627, 1.818625, 1.818625, 
    1.818627, 1.818625, 1.818629, 1.818626, 1.818631, 1.818629, 1.818631, 
    1.818631, 1.818632, 1.818632, 1.818633, 1.818635, 1.818635, 1.818636, 
    1.818621, 1.818622, 1.818622, 1.818623, 1.818624, 1.818625, 1.818628, 
    1.818627, 1.818628, 1.818629, 1.818626, 1.818628, 1.818623, 1.818624, 
    1.818623, 1.818621, 1.818627, 1.818624, 1.818629, 1.818628, 1.818632, 
    1.81863, 1.818635, 1.818636, 1.818638, 1.81864, 1.818623, 1.818622, 
    1.818623, 1.818625, 1.818626, 1.818628, 1.818628, 1.818628, 1.818629, 
    1.81863, 1.818629, 1.81863, 1.818624, 1.818627, 1.818622, 1.818623, 
    1.818625, 1.818624, 1.818627, 1.818627, 1.81863, 1.818628, 1.818636, 
    1.818633, 1.818642, 1.818639, 1.818622, 1.818623, 1.818625, 1.818624, 
    1.818628, 1.818629, 1.81863, 1.818631, 1.818631, 1.818631, 1.81863, 
    1.818631, 1.818628, 1.81863, 1.818625, 1.818626, 1.818626, 1.818625, 
    1.818627, 1.818629, 1.818629, 1.818629, 1.818631, 1.818628, 1.818636, 
    1.818631, 1.818624, 1.818625, 1.818625, 1.818625, 1.818629, 1.818627, 
    1.818631, 1.81863, 1.818632, 1.818631, 1.818631, 1.81863, 1.818629, 
    1.818627, 1.818626, 1.818625, 1.818625, 1.818626, 1.818629, 1.818631, 
    1.81863, 1.818632, 1.818628, 1.81863, 1.818629, 1.818631, 1.818627, 
    1.81863, 1.818626, 1.818626, 1.818627, 1.81863, 1.81863, 1.818631, 
    1.81863, 1.818629, 1.818628, 1.818627, 1.818627, 1.818626, 1.818625, 
    1.818626, 1.818627, 1.818629, 1.818631, 1.818632, 1.818633, 1.818635, 
    1.818633, 1.818636, 1.818634, 1.818638, 1.81863, 1.818634, 1.818627, 
    1.818628, 1.818629, 1.818632, 1.818631, 1.818632, 1.818628, 1.818626, 
    1.818626, 1.818625, 1.818626, 1.818626, 1.818627, 1.818627, 1.818629, 
    1.818628, 1.818631, 1.818632, 1.818636, 1.818638, 1.818641, 1.818642, 
    1.818642, 1.818642,
  1.818569, 1.81857, 1.81857, 1.818572, 1.818571, 1.818572, 1.818569, 
    1.81857, 1.81857, 1.818569, 1.818574, 1.818572, 1.818577, 1.818576, 
    1.81858, 1.818577, 1.818581, 1.81858, 1.818582, 1.818581, 1.818584, 
    1.818582, 1.818585, 1.818583, 1.818584, 1.818582, 1.818572, 1.818574, 
    1.818572, 1.818572, 1.818572, 1.818571, 1.81857, 1.818568, 1.818569, 
    1.81857, 1.818572, 1.818572, 1.818574, 1.818574, 1.818576, 1.818575, 
    1.818579, 1.818578, 1.818581, 1.818581, 1.818581, 1.818581, 1.818581, 
    1.81858, 1.818581, 1.818579, 1.818575, 1.818576, 1.818573, 1.818571, 
    1.818569, 1.818568, 1.818568, 1.818568, 1.81857, 1.818571, 1.818572, 
    1.818573, 1.818574, 1.818576, 1.818577, 1.818579, 1.818579, 1.81858, 
    1.81858, 1.818582, 1.818581, 1.818582, 1.81858, 1.818581, 1.818579, 
    1.818579, 1.818574, 1.818572, 1.818571, 1.81857, 1.818568, 1.81857, 
    1.818569, 1.81857, 1.818571, 1.818571, 1.818573, 1.818572, 1.818577, 
    1.818575, 1.81858, 1.818579, 1.818581, 1.81858, 1.818581, 1.81858, 
    1.818582, 1.818583, 1.818582, 1.818583, 1.81858, 1.818581, 1.818571, 
    1.818571, 1.818571, 1.81857, 1.81857, 1.818568, 1.81857, 1.81857, 
    1.818571, 1.818572, 1.818572, 1.818574, 1.818575, 1.818578, 1.818579, 
    1.81858, 1.818579, 1.81858, 1.818579, 1.818579, 1.818582, 1.818581, 
    1.818583, 1.818583, 1.818582, 1.818583, 1.818571, 1.81857, 1.818569, 
    1.81857, 1.818568, 1.818569, 1.81857, 1.818572, 1.818573, 1.818573, 
    1.818574, 1.818575, 1.818577, 1.818579, 1.81858, 1.81858, 1.81858, 
    1.818581, 1.81858, 1.818581, 1.818581, 1.818581, 1.818583, 1.818582, 
    1.818583, 1.818583, 1.81857, 1.818571, 1.818571, 1.818571, 1.818571, 
    1.818573, 1.818573, 1.818576, 1.818575, 1.818577, 1.818575, 1.818576, 
    1.818577, 1.818575, 1.818579, 1.818576, 1.818581, 1.818578, 1.818581, 
    1.81858, 1.818581, 1.818582, 1.818583, 1.818584, 1.818584, 1.818585, 
    1.818572, 1.818573, 1.818573, 1.818574, 1.818574, 1.818576, 1.818578, 
    1.818577, 1.818578, 1.818579, 1.818576, 1.818578, 1.818573, 1.818574, 
    1.818574, 1.818572, 1.818577, 1.818574, 1.818579, 1.818578, 1.818582, 
    1.81858, 1.818584, 1.818585, 1.818587, 1.818589, 1.818573, 1.818573, 
    1.818574, 1.818575, 1.818576, 1.818578, 1.818578, 1.818578, 1.818579, 
    1.81858, 1.818578, 1.81858, 1.818574, 1.818577, 1.818573, 1.818574, 
    1.818575, 1.818574, 1.818577, 1.818577, 1.818579, 1.818578, 1.818585, 
    1.818582, 1.81859, 1.818588, 1.818573, 1.818573, 1.818576, 1.818575, 
    1.818578, 1.818579, 1.818579, 1.81858, 1.81858, 1.818581, 1.81858, 
    1.818581, 1.818578, 1.818579, 1.818576, 1.818576, 1.818576, 1.818576, 
    1.818577, 1.818578, 1.818578, 1.818579, 1.81858, 1.818578, 1.818585, 
    1.818581, 1.818574, 1.818575, 1.818576, 1.818575, 1.818579, 1.818577, 
    1.818581, 1.81858, 1.818582, 1.818581, 1.818581, 1.81858, 1.818579, 
    1.818577, 1.818576, 1.818575, 1.818575, 1.818576, 1.818578, 1.81858, 
    1.81858, 1.818581, 1.818578, 1.818579, 1.818579, 1.81858, 1.818577, 
    1.81858, 1.818576, 1.818576, 1.818577, 1.818579, 1.81858, 1.81858, 
    1.81858, 1.818579, 1.818578, 1.818577, 1.818577, 1.818576, 1.818576, 
    1.818576, 1.818577, 1.818579, 1.81858, 1.818582, 1.818582, 1.818584, 
    1.818583, 1.818585, 1.818583, 1.818587, 1.81858, 1.818583, 1.818577, 
    1.818578, 1.818579, 1.818582, 1.81858, 1.818582, 1.818578, 1.818577, 
    1.818576, 1.818575, 1.818576, 1.818576, 1.818577, 1.818577, 1.818579, 
    1.818578, 1.818581, 1.818582, 1.818585, 1.818587, 1.818589, 1.81859, 
    1.81859, 1.81859,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL2_HR_S1 =
  1.292694e-09, 1.298399e-09, 1.29729e-09, 1.301891e-09, 1.299339e-09, 
    1.302352e-09, 1.293851e-09, 1.298625e-09, 1.295578e-09, 1.293208e-09, 
    1.310821e-09, 1.302097e-09, 1.319885e-09, 1.31432e-09, 1.328301e-09, 
    1.319019e-09, 1.330172e-09, 1.328033e-09, 1.334472e-09, 1.332628e-09, 
    1.340863e-09, 1.335324e-09, 1.345133e-09, 1.339541e-09, 1.340415e-09, 
    1.335141e-09, 1.303853e-09, 1.309735e-09, 1.303504e-09, 1.304343e-09, 
    1.303966e-09, 1.299392e-09, 1.297086e-09, 1.292259e-09, 1.293135e-09, 
    1.296681e-09, 1.30472e-09, 1.301991e-09, 1.308869e-09, 1.308714e-09, 
    1.316371e-09, 1.312919e-09, 1.32579e-09, 1.322132e-09, 1.332705e-09, 
    1.330046e-09, 1.33258e-09, 1.331811e-09, 1.33259e-09, 1.32869e-09, 
    1.330361e-09, 1.326929e-09, 1.313565e-09, 1.317493e-09, 1.30578e-09, 
    1.298737e-09, 1.29406e-09, 1.290742e-09, 1.291211e-09, 1.292105e-09, 
    1.296702e-09, 1.301024e-09, 1.304317e-09, 1.306521e-09, 1.308691e-09, 
    1.315262e-09, 1.318741e-09, 1.32653e-09, 1.325125e-09, 1.327506e-09, 
    1.329781e-09, 1.333601e-09, 1.332972e-09, 1.334655e-09, 1.327443e-09, 
    1.332236e-09, 1.324324e-09, 1.326488e-09, 1.309281e-09, 1.302727e-09, 
    1.299941e-09, 1.297503e-09, 1.291572e-09, 1.295668e-09, 1.294053e-09, 
    1.297895e-09, 1.300336e-09, 1.299129e-09, 1.306581e-09, 1.303683e-09, 
    1.318947e-09, 1.312372e-09, 1.329516e-09, 1.325413e-09, 1.330499e-09, 
    1.327904e-09, 1.33235e-09, 1.328349e-09, 1.335281e-09, 1.336791e-09, 
    1.335759e-09, 1.339722e-09, 1.328127e-09, 1.332579e-09, 1.299095e-09, 
    1.299292e-09, 1.300209e-09, 1.296176e-09, 1.29593e-09, 1.292234e-09, 
    1.295523e-09, 1.296923e-09, 1.300478e-09, 1.30258e-09, 1.304579e-09, 
    1.308974e-09, 1.313883e-09, 1.320747e-09, 1.325679e-09, 1.328985e-09, 
    1.326958e-09, 1.328748e-09, 1.326747e-09, 1.325809e-09, 1.336225e-09, 
    1.330376e-09, 1.339152e-09, 1.338667e-09, 1.334695e-09, 1.338721e-09, 
    1.29943e-09, 1.298297e-09, 1.294363e-09, 1.297442e-09, 1.291832e-09, 
    1.294972e-09, 1.296777e-09, 1.303744e-09, 1.305275e-09, 1.306694e-09, 
    1.309498e-09, 1.313095e-09, 1.319407e-09, 1.324899e-09, 1.329913e-09, 
    1.329546e-09, 1.329675e-09, 1.330795e-09, 1.328021e-09, 1.331251e-09, 
    1.331793e-09, 1.330376e-09, 1.338602e-09, 1.336251e-09, 1.338656e-09, 
    1.337126e-09, 1.298665e-09, 1.300572e-09, 1.299542e-09, 1.301479e-09, 
    1.300114e-09, 1.306183e-09, 1.308003e-09, 1.316519e-09, 1.313025e-09, 
    1.318587e-09, 1.31359e-09, 1.314475e-09, 1.318768e-09, 1.31386e-09, 
    1.324596e-09, 1.317317e-09, 1.330839e-09, 1.323569e-09, 1.331295e-09, 
    1.329892e-09, 1.332214e-09, 1.334295e-09, 1.336912e-09, 1.341741e-09, 
    1.340623e-09, 1.344661e-09, 1.303415e-09, 1.305888e-09, 1.30567e-09, 
    1.308259e-09, 1.310173e-09, 1.314322e-09, 1.320977e-09, 1.318474e-09, 
    1.323069e-09, 1.323991e-09, 1.317011e-09, 1.321297e-09, 1.307543e-09, 
    1.309765e-09, 1.308442e-09, 1.30361e-09, 1.319051e-09, 1.311126e-09, 
    1.325761e-09, 1.321467e-09, 1.333998e-09, 1.327766e-09, 1.340007e-09, 
    1.34524e-09, 1.350166e-09, 1.355922e-09, 1.307238e-09, 1.305557e-09, 
    1.308566e-09, 1.312729e-09, 1.316593e-09, 1.321729e-09, 1.322255e-09, 
    1.323217e-09, 1.325709e-09, 1.327805e-09, 1.323521e-09, 1.32833e-09, 
    1.31028e-09, 1.319739e-09, 1.304922e-09, 1.309383e-09, 1.312484e-09, 
    1.311124e-09, 1.318188e-09, 1.319854e-09, 1.32662e-09, 1.323122e-09, 
    1.343948e-09, 1.334734e-09, 1.360306e-09, 1.353159e-09, 1.30497e-09, 
    1.307232e-09, 1.315104e-09, 1.311359e-09, 1.322072e-09, 1.324709e-09, 
    1.326853e-09, 1.329593e-09, 1.329889e-09, 1.331513e-09, 1.328852e-09, 
    1.331408e-09, 1.32174e-09, 1.32606e-09, 1.314205e-09, 1.31709e-09, 
    1.315763e-09, 1.314307e-09, 1.318801e-09, 1.323588e-09, 1.323691e-09, 
    1.325226e-09, 1.329551e-09, 1.322115e-09, 1.345137e-09, 1.330918e-09, 
    1.309699e-09, 1.314055e-09, 1.314678e-09, 1.31299e-09, 1.324445e-09, 
    1.320294e-09, 1.331474e-09, 1.328452e-09, 1.333403e-09, 1.330943e-09, 
    1.330581e-09, 1.327421e-09, 1.325454e-09, 1.320484e-09, 1.316441e-09, 
    1.313235e-09, 1.31398e-09, 1.317502e-09, 1.323881e-09, 1.329916e-09, 
    1.328594e-09, 1.333027e-09, 1.321295e-09, 1.326214e-09, 1.324313e-09, 
    1.32927e-09, 1.318408e-09, 1.327657e-09, 1.316044e-09, 1.317062e-09, 
    1.320212e-09, 1.326547e-09, 1.32795e-09, 1.329446e-09, 1.328523e-09, 
    1.324043e-09, 1.323309e-09, 1.320135e-09, 1.319259e-09, 1.31684e-09, 
    1.314838e-09, 1.316667e-09, 1.318588e-09, 1.324045e-09, 1.328962e-09, 
    1.334324e-09, 1.335636e-09, 1.341901e-09, 1.336801e-09, 1.345216e-09, 
    1.338061e-09, 1.350448e-09, 1.328193e-09, 1.337851e-09, 1.320355e-09, 
    1.32224e-09, 1.325649e-09, 1.333468e-09, 1.329247e-09, 1.334184e-09, 
    1.32328e-09, 1.317624e-09, 1.31616e-09, 1.31343e-09, 1.316223e-09, 
    1.315996e-09, 1.318668e-09, 1.317809e-09, 1.324226e-09, 1.320779e-09, 
    1.330572e-09, 1.334145e-09, 1.344238e-09, 1.350426e-09, 1.356725e-09, 
    1.359506e-09, 1.360353e-09, 1.360706e-09 ;

 SOIL2_HR_S3 =
  9.233531e-11, 9.274279e-11, 9.266358e-11, 9.299224e-11, 9.280993e-11, 
    9.302513e-11, 9.241793e-11, 9.275895e-11, 9.254125e-11, 9.237201e-11, 
    9.363006e-11, 9.30069e-11, 9.427752e-11, 9.388003e-11, 9.487861e-11, 
    9.421566e-11, 9.50123e-11, 9.485952e-11, 9.531945e-11, 9.518768e-11, 
    9.577595e-11, 9.538027e-11, 9.608095e-11, 9.568147e-11, 9.574395e-11, 
    9.536721e-11, 9.313233e-11, 9.355247e-11, 9.310743e-11, 9.316734e-11, 
    9.314046e-11, 9.281369e-11, 9.2649e-11, 9.230418e-11, 9.236679e-11, 
    9.262006e-11, 9.319428e-11, 9.299937e-11, 9.349065e-11, 9.347956e-11, 
    9.402653e-11, 9.377991e-11, 9.469932e-11, 9.4438e-11, 9.519318e-11, 
    9.500326e-11, 9.518426e-11, 9.512938e-11, 9.518497e-11, 9.490642e-11, 
    9.502577e-11, 9.478067e-11, 9.382609e-11, 9.410661e-11, 9.326998e-11, 
    9.276693e-11, 9.243288e-11, 9.219583e-11, 9.222934e-11, 9.229322e-11, 
    9.262154e-11, 9.293025e-11, 9.316552e-11, 9.332289e-11, 9.347797e-11, 
    9.394731e-11, 9.419579e-11, 9.475215e-11, 9.465177e-11, 9.482184e-11, 
    9.498436e-11, 9.525719e-11, 9.521229e-11, 9.533248e-11, 9.481737e-11, 
    9.515971e-11, 9.459458e-11, 9.474914e-11, 9.352005e-11, 9.305196e-11, 
    9.285294e-11, 9.26788e-11, 9.225511e-11, 9.254769e-11, 9.243235e-11, 
    9.270678e-11, 9.288115e-11, 9.279491e-11, 9.33272e-11, 9.312025e-11, 
    9.421051e-11, 9.374088e-11, 9.49654e-11, 9.467237e-11, 9.503565e-11, 
    9.485027e-11, 9.516789e-11, 9.488204e-11, 9.537723e-11, 9.548505e-11, 
    9.541137e-11, 9.569445e-11, 9.486619e-11, 9.518425e-11, 9.279249e-11, 
    9.280655e-11, 9.287209e-11, 9.258402e-11, 9.256641e-11, 9.230246e-11, 
    9.253733e-11, 9.263734e-11, 9.289126e-11, 9.304145e-11, 9.318422e-11, 
    9.349815e-11, 9.384876e-11, 9.433907e-11, 9.469137e-11, 9.492751e-11, 
    9.478272e-11, 9.491055e-11, 9.476764e-11, 9.470066e-11, 9.544465e-11, 
    9.502688e-11, 9.565373e-11, 9.561904e-11, 9.533534e-11, 9.562295e-11, 
    9.281644e-11, 9.273549e-11, 9.245447e-11, 9.26744e-11, 9.227372e-11, 
    9.249799e-11, 9.262694e-11, 9.312456e-11, 9.323391e-11, 9.333529e-11, 
    9.353554e-11, 9.379253e-11, 9.424336e-11, 9.463566e-11, 9.499382e-11, 
    9.496758e-11, 9.497681e-11, 9.505682e-11, 9.485863e-11, 9.508935e-11, 
    9.512807e-11, 9.502683e-11, 9.56144e-11, 9.544653e-11, 9.56183e-11, 
    9.550901e-11, 9.276181e-11, 9.289799e-11, 9.28244e-11, 9.296279e-11, 
    9.286529e-11, 9.329882e-11, 9.342881e-11, 9.40371e-11, 9.378746e-11, 
    9.418478e-11, 9.382783e-11, 9.389108e-11, 9.419771e-11, 9.384712e-11, 
    9.461402e-11, 9.409405e-11, 9.505993e-11, 9.454063e-11, 9.509247e-11, 
    9.499227e-11, 9.515817e-11, 9.530676e-11, 9.54937e-11, 9.583864e-11, 
    9.575877e-11, 9.604725e-11, 9.310105e-11, 9.327769e-11, 9.326215e-11, 
    9.344703e-11, 9.358377e-11, 9.388014e-11, 9.43555e-11, 9.417675e-11, 
    9.450493e-11, 9.457082e-11, 9.407223e-11, 9.437833e-11, 9.339593e-11, 
    9.355463e-11, 9.346015e-11, 9.311497e-11, 9.421792e-11, 9.365186e-11, 
    9.469718e-11, 9.43905e-11, 9.528557e-11, 9.484041e-11, 9.57148e-11, 
    9.608858e-11, 9.644045e-11, 9.68516e-11, 9.337412e-11, 9.325409e-11, 
    9.346902e-11, 9.376638e-11, 9.404234e-11, 9.44092e-11, 9.444675e-11, 
    9.451548e-11, 9.469352e-11, 9.484321e-11, 9.45372e-11, 9.488074e-11, 
    9.359141e-11, 9.426706e-11, 9.32087e-11, 9.352735e-11, 9.374886e-11, 
    9.365171e-11, 9.415632e-11, 9.427525e-11, 9.475856e-11, 9.450873e-11, 
    9.599631e-11, 9.533813e-11, 9.716473e-11, 9.665421e-11, 9.321215e-11, 
    9.337371e-11, 9.393603e-11, 9.366848e-11, 9.44337e-11, 9.462207e-11, 
    9.477522e-11, 9.497095e-11, 9.49921e-11, 9.510808e-11, 9.491802e-11, 
    9.510058e-11, 9.440999e-11, 9.471859e-11, 9.387177e-11, 9.407786e-11, 
    9.398306e-11, 9.387906e-11, 9.420004e-11, 9.454201e-11, 9.454934e-11, 
    9.465899e-11, 9.496794e-11, 9.443681e-11, 9.608122e-11, 9.506559e-11, 
    9.35499e-11, 9.386109e-11, 9.390557e-11, 9.378501e-11, 9.460319e-11, 
    9.430672e-11, 9.510526e-11, 9.488944e-11, 9.524306e-11, 9.506734e-11, 
    9.504148e-11, 9.48158e-11, 9.467529e-11, 9.432031e-11, 9.40315e-11, 
    9.38025e-11, 9.385575e-11, 9.41073e-11, 9.456293e-11, 9.499401e-11, 
    9.489957e-11, 9.521619e-11, 9.437822e-11, 9.472957e-11, 9.459376e-11, 
    9.494789e-11, 9.4172e-11, 9.483263e-11, 9.400313e-11, 9.407586e-11, 
    9.430084e-11, 9.475339e-11, 9.485355e-11, 9.496046e-11, 9.48945e-11, 
    9.45745e-11, 9.452209e-11, 9.429537e-11, 9.423276e-11, 9.406002e-11, 
    9.391701e-11, 9.404767e-11, 9.418489e-11, 9.457465e-11, 9.492589e-11, 
    9.530887e-11, 9.540261e-11, 9.585005e-11, 9.548578e-11, 9.608687e-11, 
    9.557578e-11, 9.646056e-11, 9.487096e-11, 9.55608e-11, 9.431108e-11, 
    9.444571e-11, 9.46892e-11, 9.524774e-11, 9.494622e-11, 9.529886e-11, 
    9.452004e-11, 9.411597e-11, 9.401146e-11, 9.381642e-11, 9.401591e-11, 
    9.399969e-11, 9.419059e-11, 9.412925e-11, 9.458759e-11, 9.434138e-11, 
    9.504083e-11, 9.529608e-11, 9.601701e-11, 9.645897e-11, 9.690893e-11, 
    9.710758e-11, 9.716804e-11, 9.719332e-11 ;

 SOIL3C =
  5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.782611, 5.78261, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 5.782611, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 
    5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.78261, 5.78261, 5.78261, 5.78261, 
    5.78261, 5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.78261, 5.78261, 5.78261, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 
    5.782611, 5.782611, 5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 
    5.78261, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.78261, 5.78261, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 5.782611, 
    5.782611, 5.782611, 5.782611 ;

 SOIL3C_TO_SOIL1C =
  2.549161e-11, 2.560408e-11, 2.558222e-11, 2.567293e-11, 2.562261e-11, 
    2.568201e-11, 2.551441e-11, 2.560854e-11, 2.554845e-11, 2.550174e-11, 
    2.584898e-11, 2.567698e-11, 2.602769e-11, 2.591798e-11, 2.61936e-11, 
    2.601061e-11, 2.62305e-11, 2.618833e-11, 2.631528e-11, 2.627891e-11, 
    2.644128e-11, 2.633206e-11, 2.652546e-11, 2.64152e-11, 2.643244e-11, 
    2.632846e-11, 2.57116e-11, 2.582756e-11, 2.570473e-11, 2.572126e-11, 
    2.571384e-11, 2.562365e-11, 2.557819e-11, 2.548302e-11, 2.550029e-11, 
    2.55702e-11, 2.57287e-11, 2.56749e-11, 2.58105e-11, 2.580744e-11, 
    2.595841e-11, 2.589034e-11, 2.614411e-11, 2.607198e-11, 2.628043e-11, 
    2.6228e-11, 2.627796e-11, 2.626281e-11, 2.627816e-11, 2.620128e-11, 
    2.623422e-11, 2.616657e-11, 2.590309e-11, 2.598052e-11, 2.574959e-11, 
    2.561074e-11, 2.551854e-11, 2.545311e-11, 2.546236e-11, 2.547999e-11, 
    2.557061e-11, 2.565582e-11, 2.572076e-11, 2.57642e-11, 2.5807e-11, 
    2.593655e-11, 2.600513e-11, 2.61587e-11, 2.613099e-11, 2.617793e-11, 
    2.622279e-11, 2.629809e-11, 2.62857e-11, 2.631888e-11, 2.61767e-11, 
    2.627119e-11, 2.61152e-11, 2.615786e-11, 2.581861e-11, 2.568941e-11, 
    2.563448e-11, 2.558642e-11, 2.546947e-11, 2.555023e-11, 2.551839e-11, 
    2.559414e-11, 2.564227e-11, 2.561847e-11, 2.576539e-11, 2.570827e-11, 
    2.60092e-11, 2.587957e-11, 2.621756e-11, 2.613667e-11, 2.623694e-11, 
    2.618578e-11, 2.627345e-11, 2.619455e-11, 2.633123e-11, 2.636099e-11, 
    2.634065e-11, 2.641878e-11, 2.619017e-11, 2.627796e-11, 2.56178e-11, 
    2.562168e-11, 2.563977e-11, 2.556026e-11, 2.555539e-11, 2.548254e-11, 
    2.554737e-11, 2.557497e-11, 2.564506e-11, 2.568651e-11, 2.572592e-11, 
    2.581257e-11, 2.590934e-11, 2.604468e-11, 2.614192e-11, 2.62071e-11, 
    2.616713e-11, 2.620242e-11, 2.616297e-11, 2.614448e-11, 2.634983e-11, 
    2.623452e-11, 2.640754e-11, 2.639797e-11, 2.631967e-11, 2.639905e-11, 
    2.562441e-11, 2.560207e-11, 2.55245e-11, 2.55852e-11, 2.547461e-11, 
    2.553651e-11, 2.55721e-11, 2.570945e-11, 2.573964e-11, 2.576762e-11, 
    2.582289e-11, 2.589383e-11, 2.601826e-11, 2.612654e-11, 2.62254e-11, 
    2.621816e-11, 2.622071e-11, 2.624279e-11, 2.618809e-11, 2.625177e-11, 
    2.626245e-11, 2.623451e-11, 2.639669e-11, 2.635035e-11, 2.639777e-11, 
    2.63676e-11, 2.560933e-11, 2.564692e-11, 2.562661e-11, 2.56648e-11, 
    2.563789e-11, 2.575755e-11, 2.579343e-11, 2.596133e-11, 2.589243e-11, 
    2.600209e-11, 2.590357e-11, 2.592102e-11, 2.600566e-11, 2.590889e-11, 
    2.612057e-11, 2.597705e-11, 2.624364e-11, 2.610031e-11, 2.625263e-11, 
    2.622497e-11, 2.627076e-11, 2.631178e-11, 2.636338e-11, 2.645858e-11, 
    2.643654e-11, 2.651616e-11, 2.570296e-11, 2.575172e-11, 2.574743e-11, 
    2.579846e-11, 2.58362e-11, 2.591801e-11, 2.604921e-11, 2.599988e-11, 
    2.609046e-11, 2.610864e-11, 2.597103e-11, 2.605552e-11, 2.578436e-11, 
    2.582816e-11, 2.580208e-11, 2.570681e-11, 2.601124e-11, 2.5855e-11, 
    2.614352e-11, 2.605888e-11, 2.630593e-11, 2.618306e-11, 2.64244e-11, 
    2.652757e-11, 2.662469e-11, 2.673817e-11, 2.577834e-11, 2.574521e-11, 
    2.580453e-11, 2.588661e-11, 2.596278e-11, 2.606404e-11, 2.60744e-11, 
    2.609337e-11, 2.614251e-11, 2.618383e-11, 2.609936e-11, 2.619419e-11, 
    2.583831e-11, 2.60248e-11, 2.573268e-11, 2.582063e-11, 2.588177e-11, 
    2.585496e-11, 2.599424e-11, 2.602706e-11, 2.616046e-11, 2.609151e-11, 
    2.65021e-11, 2.632043e-11, 2.68246e-11, 2.668369e-11, 2.573363e-11, 
    2.577823e-11, 2.593343e-11, 2.585959e-11, 2.60708e-11, 2.612279e-11, 
    2.616506e-11, 2.621909e-11, 2.622493e-11, 2.625694e-11, 2.620448e-11, 
    2.625487e-11, 2.606425e-11, 2.614943e-11, 2.59157e-11, 2.597258e-11, 
    2.594642e-11, 2.591771e-11, 2.600631e-11, 2.610069e-11, 2.610272e-11, 
    2.613298e-11, 2.621826e-11, 2.607166e-11, 2.652554e-11, 2.624521e-11, 
    2.582685e-11, 2.591275e-11, 2.592503e-11, 2.589175e-11, 2.611758e-11, 
    2.603575e-11, 2.625616e-11, 2.619659e-11, 2.629419e-11, 2.624569e-11, 
    2.623855e-11, 2.617626e-11, 2.613748e-11, 2.60395e-11, 2.595978e-11, 
    2.589658e-11, 2.591127e-11, 2.598071e-11, 2.610647e-11, 2.622545e-11, 
    2.619939e-11, 2.628678e-11, 2.605548e-11, 2.615246e-11, 2.611498e-11, 
    2.621272e-11, 2.599856e-11, 2.618091e-11, 2.595195e-11, 2.597203e-11, 
    2.603412e-11, 2.615904e-11, 2.618668e-11, 2.621619e-11, 2.619798e-11, 
    2.610966e-11, 2.60952e-11, 2.603262e-11, 2.601534e-11, 2.596766e-11, 
    2.592818e-11, 2.596425e-11, 2.600212e-11, 2.61097e-11, 2.620665e-11, 
    2.631236e-11, 2.633823e-11, 2.646173e-11, 2.636119e-11, 2.65271e-11, 
    2.638603e-11, 2.663024e-11, 2.619149e-11, 2.638189e-11, 2.603695e-11, 
    2.607411e-11, 2.614132e-11, 2.629548e-11, 2.621226e-11, 2.63096e-11, 
    2.609463e-11, 2.59831e-11, 2.595425e-11, 2.590042e-11, 2.595548e-11, 
    2.595101e-11, 2.60037e-11, 2.598676e-11, 2.611327e-11, 2.604532e-11, 
    2.623837e-11, 2.630883e-11, 2.650781e-11, 2.66298e-11, 2.6754e-11, 
    2.680882e-11, 2.682551e-11, 2.683249e-11 ;

 SOIL3C_vr =
  20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 20.00008, 
    20.00008, 20.00008,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 20.00007, 20.00007, 
    20.00006, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00007, 20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00006, 
    20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 
    20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00007, 20.00006, 20.00007, 20.00007, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00007, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007, 20.00007, 20.00007, 20.00006, 20.00007, 20.00006, 
    20.00006, 20.00006, 20.00007, 20.00006, 20.00007, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 20.00007, 
    20.00007, 20.00007,
  20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 20.00006, 
    20.00006, 20.00006,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N =
  0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 0.5256919, 
    0.5256919, 0.5256919 ;

 SOIL3N_TNDNCY_VERT_TRANS =
  1.28498e-20, -1.28498e-20, -1.027984e-20, -1.541976e-20, 1.798972e-20, 
    -5.139921e-21, -1.027984e-20, -2.569961e-21, 2.569961e-21, -1.003089e-36, 
    -1.027984e-20, 2.569961e-21, 2.569961e-21, -2.055969e-20, -5.139921e-21, 
    2.569961e-21, 5.139921e-21, 2.569961e-21, -5.139921e-21, 2.569961e-21, 
    1.027984e-20, 1.28498e-20, 1.798972e-20, 1.027984e-20, 5.139921e-21, 
    -5.139921e-21, 2.569961e-21, -7.709882e-21, -1.798972e-20, 1.027984e-20, 
    1.28498e-20, 1.027984e-20, 5.139921e-21, -1.027984e-20, 5.139921e-21, 
    -5.139921e-21, -7.709882e-21, 1.28498e-20, -5.139921e-21, -7.709882e-21, 
    -1.027984e-20, -1.28498e-20, 2.569961e-21, -5.139921e-21, 1.798972e-20, 
    5.139921e-21, 5.139921e-21, -7.709882e-21, 0, -2.569961e-21, 
    -7.709882e-21, 1.28498e-20, 1.28498e-20, -2.569961e-21, -1.798972e-20, 
    2.569961e-21, 1.28498e-20, 1.798972e-20, -1.003089e-36, -7.709882e-21, 
    1.003089e-36, -1.027984e-20, -5.139921e-21, -2.569961e-21, 7.709882e-21, 
    -5.139921e-21, 1.28498e-20, 7.709882e-21, -1.28498e-20, 1.027984e-20, 0, 
    -5.139921e-21, -2.569961e-21, 2.569961e-21, -1.003089e-36, 5.139921e-21, 
    7.709882e-21, 2.569961e-21, -1.027984e-20, 2.312965e-20, 0, 2.312965e-20, 
    1.541976e-20, -2.569961e-21, -1.541976e-20, 2.569961e-21, -7.709882e-21, 
    -5.139921e-21, 2.569961e-21, -2.569961e-21, 7.709882e-21, -1.003089e-36, 
    0, -1.798972e-20, 1.027984e-20, 7.709882e-21, -1.798972e-20, 
    1.003089e-36, 2.569961e-21, 1.541976e-20, -1.28498e-20, -2.569961e-21, 
    -5.139921e-21, -2.569961e-21, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    1.003089e-36, 0, -1.003089e-36, 7.709882e-21, 1.541976e-20, 
    -2.569961e-21, 5.139921e-21, -5.139921e-21, -2.569961e-21, 5.139921e-21, 
    -1.28498e-20, -1.003089e-36, -5.139921e-21, -7.709882e-21, -5.139921e-21, 
    -1.027984e-20, -1.027984e-20, -7.709882e-21, 0, 7.709882e-21, 
    1.027984e-20, -5.139921e-21, 1.28498e-20, 1.541976e-20, 5.139921e-21, 
    -1.541976e-20, 7.709882e-21, -1.027984e-20, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 7.709882e-21, 2.055969e-20, -2.569961e-21, 
    0, -5.139921e-21, -2.569961e-21, -1.28498e-20, 5.139921e-21, 
    -5.139921e-21, 1.28498e-20, 2.055969e-20, 1.28498e-20, -1.28498e-20, 
    1.027984e-20, -1.003089e-36, -2.569961e-21, -5.139921e-21, 5.139921e-21, 
    -1.027984e-20, 2.569961e-21, -1.027984e-20, -1.28498e-20, 1.027984e-20, 
    2.055969e-20, 0, 7.709882e-21, 1.003089e-36, -5.139921e-21, 1.798972e-20, 
    1.28498e-20, -2.055969e-20, 5.139921e-21, -2.055969e-20, 5.139921e-21, 
    -1.027984e-20, 2.569961e-21, 2.569961e-21, 1.28498e-20, -1.28498e-20, 
    -5.139921e-21, -5.139921e-21, -7.709882e-21, -1.003089e-36, 5.139921e-21, 
    5.139921e-21, -1.027984e-20, 1.027984e-20, -1.027984e-20, 5.139921e-21, 
    2.055969e-20, -5.139921e-21, 5.139921e-21, 5.139921e-21, -2.569961e-20, 
    0, -1.027984e-20, 2.569961e-21, 1.28498e-20, -1.28498e-20, -1.003089e-36, 
    -1.027984e-20, 7.709882e-21, -2.569961e-21, -7.709882e-21, 2.569961e-21, 
    5.139921e-21, 1.798972e-20, 1.28498e-20, 2.569961e-21, -1.798972e-20, 
    -1.003089e-36, 1.027984e-20, -1.003089e-36, 2.569961e-21, 2.569961e-21, 
    7.709882e-21, 5.139921e-21, 2.569961e-21, 7.709882e-21, -1.027984e-20, 
    -1.027984e-20, 2.055969e-20, -2.569961e-21, 2.569961e-21, -1.28498e-20, 
    2.569961e-21, -2.569961e-21, 1.28498e-20, -1.027984e-20, -2.569961e-21, 
    -1.003089e-36, 1.027984e-20, -2.569961e-21, 2.569961e-21, 1.28498e-20, 
    -2.569961e-21, 2.569961e-21, 1.027984e-20, 1.541976e-20, -5.139921e-21, 
    -5.139921e-21, 2.569961e-21, 0, -2.569961e-21, 7.709882e-21, 
    1.003089e-36, -1.027984e-20, -1.28498e-20, -7.709882e-21, 7.709882e-21, 
    2.569961e-21, 7.709882e-21, -5.139921e-21, -7.709882e-21, -1.541976e-20, 
    2.569961e-21, 0, 1.28498e-20, -1.541976e-20, 1.003089e-36, -2.569961e-21, 
    1.541976e-20, -1.541976e-20, 1.027984e-20, 0, -1.027984e-20, 
    1.003089e-36, -5.139921e-21, 2.569961e-21, 1.28498e-20, -7.709882e-21, 
    5.139921e-21, -5.139921e-21, -1.027984e-20, -5.139921e-21, -5.139921e-21, 
    1.027984e-20, 1.003089e-36, -1.798972e-20, 5.139921e-21, 5.139921e-21, 
    -1.027984e-20, -7.709882e-21, -1.027984e-20, -1.003089e-36, 1.027984e-20, 
    -2.569961e-21, -1.027984e-20, 1.027984e-20, 1.027984e-20, 7.709882e-21, 
    5.139921e-21, 5.139921e-21, 1.28498e-20, -5.139921e-21, 1.798972e-20, 
    -1.798972e-20, -5.015443e-37, 5.139921e-21, -2.569961e-21, 5.139921e-21, 
    -2.569961e-21, 5.139921e-21, -2.569961e-21, -1.003089e-36, 2.569961e-21, 
    -1.541976e-20, 5.139921e-21, -7.709882e-21, 1.027984e-20, 1.28498e-20, 
    1.798972e-20, -5.139921e-21, 5.139921e-21, -1.003089e-36, -5.139921e-21, 
    -2.569961e-21, -2.055969e-20, 5.139921e-21, -1.003089e-36, -5.139921e-21, 
    -1.541976e-20, 0, -1.027984e-20, -7.709882e-21, 2.569961e-21, 
    1.28498e-20, -2.569961e-21, 7.709882e-21, -5.139921e-21, 1.798972e-20, 
    1.003089e-36, 5.139921e-21, -2.569961e-21, 7.709882e-21, -7.709882e-21, 
    -1.027984e-20, 5.139921e-21, -1.28498e-20,
  -2.569961e-21, -2.569961e-21, 2.569961e-21, 1.027984e-20, -1.28498e-20, 
    -2.569961e-21, 2.569961e-21, 2.569961e-21, -7.709882e-21, 5.139921e-21, 
    0, 7.709882e-21, -2.569961e-21, 0, -1.027984e-20, 0, -5.139921e-21, 
    -2.055969e-20, -2.569961e-21, 2.569961e-21, 7.709882e-21, -7.709882e-21, 
    2.569961e-21, 0, -2.569961e-21, 1.027984e-20, -2.569961e-21, 
    -2.569961e-21, 5.139921e-21, -2.569961e-21, 5.139921e-21, 7.709882e-21, 
    0, 7.709882e-21, -2.569961e-21, -5.139921e-21, -5.139921e-21, 
    2.569961e-21, -5.139921e-21, 2.569961e-21, 2.569961e-21, 7.709882e-21, 
    -7.709882e-21, -5.139921e-21, 5.139921e-21, -2.569961e-21, 1.027984e-20, 
    1.027984e-20, -2.569961e-21, 7.709882e-21, 5.139921e-21, 0, 0, 
    -1.027984e-20, 1.003089e-36, 2.569961e-21, 1.027984e-20, 2.569961e-21, 
    5.139921e-21, 2.569961e-21, -1.28498e-20, 2.569961e-21, 2.569961e-21, 
    -1.003089e-36, -7.709882e-21, 5.139921e-21, -2.569961e-21, -1.28498e-20, 
    7.709882e-21, -5.139921e-21, -1.027984e-20, -2.569961e-21, 1.027984e-20, 
    0, -1.027984e-20, 2.569961e-21, -5.139921e-21, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, 5.139921e-21, -7.709882e-21, 5.139921e-21, 
    2.569961e-21, -5.139921e-21, 2.569961e-21, -5.139921e-21, 1.003089e-36, 
    5.139921e-21, -1.027984e-20, 2.569961e-21, -2.569961e-21, 1.541976e-20, 
    5.139921e-21, -2.569961e-21, 2.569961e-21, -2.569961e-21, 5.139921e-21, 
    5.139921e-21, -2.569961e-21, -1.027984e-20, 7.709882e-21, 5.139921e-21, 
    -1.003089e-36, 2.569961e-21, 5.139921e-21, -1.28498e-20, -1.541976e-20, 
    2.569961e-21, -5.139921e-21, -5.139921e-21, 5.139921e-21, 1.027984e-20, 
    -1.027984e-20, -1.798972e-20, 1.541976e-20, -5.139921e-21, -5.139921e-21, 
    -2.569961e-21, -2.569961e-21, 1.027984e-20, 1.28498e-20, 0, 
    -2.569961e-21, -7.709882e-21, -5.139921e-21, -5.139921e-21, 
    -2.569961e-21, -5.139921e-21, 2.569961e-21, -1.003089e-36, -2.569961e-21, 
    -2.569961e-21, 1.28498e-20, 1.003089e-36, 7.709882e-21, 2.569961e-21, 
    2.569961e-21, -1.28498e-20, 7.709882e-21, 5.139921e-21, 7.709882e-21, 
    2.569961e-21, -2.569961e-21, -1.28498e-20, -5.139921e-21, 1.541976e-20, 
    -1.003089e-36, 5.139921e-21, 5.139921e-21, 2.569961e-21, -1.027984e-20, 
    0, -5.139921e-21, -5.139921e-21, 5.139921e-21, 5.139921e-21, 
    2.569961e-21, 7.709882e-21, -1.003089e-36, -7.709882e-21, -7.709882e-21, 
    1.027984e-20, -5.139921e-21, 5.139921e-21, 7.709882e-21, 2.569961e-21, 
    -1.003089e-36, -1.798972e-20, 2.569961e-21, 0, -7.709882e-21, 
    -1.027984e-20, 5.139921e-21, -7.709882e-21, -2.569961e-21, 2.569961e-21, 
    -2.569961e-21, 2.569961e-21, -1.28498e-20, -2.569961e-21, 0, 0, 
    -1.027984e-20, 5.139921e-21, 5.139921e-21, -1.28498e-20, -5.139921e-21, 
    -7.709882e-21, -2.569961e-21, -7.709882e-21, 7.709882e-21, -1.003089e-36, 
    -5.139921e-21, -5.139921e-21, -1.28498e-20, 1.027984e-20, 5.139921e-21, 
    -1.027984e-20, -5.139921e-21, -5.139921e-21, 5.139921e-21, -7.709882e-21, 
    -1.541976e-20, -2.569961e-21, 5.139921e-21, -7.709882e-21, 5.139921e-21, 
    0, -2.569961e-21, 1.28498e-20, 5.139921e-21, -1.003089e-36, 5.139921e-21, 
    2.569961e-21, 2.569961e-21, -5.139921e-21, -7.709882e-21, 2.569961e-21, 
    7.709882e-21, 2.569961e-21, -2.569961e-21, -2.569961e-21, 1.003089e-36, 
    5.139921e-21, 1.003089e-36, -1.28498e-20, -1.541976e-20, 1.003089e-36, 
    5.139921e-21, 7.709882e-21, 0, -5.139921e-21, 2.569961e-21, 2.569961e-21, 
    7.709882e-21, 0, -1.541976e-20, -7.709882e-21, -2.569961e-21, 
    -7.709882e-21, -2.569961e-21, 2.569961e-21, -1.027984e-20, -2.569961e-21, 
    -2.569961e-21, -2.055969e-20, 5.139921e-21, -5.139921e-21, 0, 
    1.027984e-20, 2.569961e-21, -2.569961e-21, 1.798972e-20, -5.139921e-21, 
    -5.139921e-21, -5.139921e-21, 1.027984e-20, 0, 0, -2.569961e-21, 
    -2.569961e-21, 7.709882e-21, 1.003089e-36, 1.28498e-20, -5.139921e-21, 
    5.139921e-21, -7.709882e-21, -1.003089e-36, 5.139921e-21, 2.569961e-21, 
    0, 7.709882e-21, 2.569961e-21, 2.569961e-21, 2.569961e-21, -5.139921e-21, 
    7.709882e-21, 1.027984e-20, -7.709882e-21, 0, 2.569961e-21, 2.569961e-21, 
    -2.569961e-21, 5.139921e-21, 2.569961e-21, -1.003089e-36, 7.709882e-21, 
    -2.569961e-21, -1.541976e-20, -2.569961e-21, 5.139921e-21, -2.569961e-21, 
    -1.027984e-20, -2.569961e-21, -1.027984e-20, 1.027984e-20, 1.027984e-20, 
    1.027984e-20, 1.027984e-20, -5.139921e-21, -2.569961e-21, 7.709882e-21, 
    1.28498e-20, -2.569961e-21, -7.709882e-21, -7.709882e-21, -2.569961e-21, 
    7.709882e-21, 1.027984e-20, -5.139921e-21, -1.003089e-36, 5.139921e-21, 
    -2.569961e-21, -2.569961e-21, -5.139921e-21, -7.709882e-21, 5.139921e-21, 
    1.027984e-20, -1.28498e-20, -2.569961e-21, 1.003089e-36, -2.569961e-21, 
    2.569961e-21, 5.139921e-21, -1.003089e-36, 1.027984e-20, 5.139921e-21, 
    2.569961e-21, -7.709882e-21, -1.027984e-20, 7.709882e-21, -1.003089e-36, 
    0, -7.709882e-21, 0, -2.569961e-21, 2.055969e-20,
  -1.027984e-20, 1.003089e-36, 1.003089e-36, -2.569961e-21, 1.798972e-20, 
    -7.709882e-21, 1.28498e-20, -1.541976e-20, 0, 0, 1.003089e-36, 0, 
    -1.541976e-20, 2.569961e-21, 2.569961e-21, 2.569961e-21, 0, 
    -2.569961e-21, 1.027984e-20, 1.027984e-20, -5.139921e-21, -2.569961e-21, 
    1.027984e-20, -1.28498e-20, 5.139921e-21, 2.569961e-21, 1.027984e-20, 
    1.003089e-36, 7.709882e-21, -1.003089e-36, -1.798972e-20, -2.569961e-21, 
    -1.28498e-20, 2.569961e-21, 1.28498e-20, 5.139921e-21, 7.709882e-21, 
    1.027984e-20, 7.709882e-21, -1.003089e-36, -5.139921e-21, -7.709882e-21, 
    7.709882e-21, 7.709882e-21, 1.003089e-36, -1.28498e-20, 7.709882e-21, 
    -5.139921e-21, 5.139921e-21, -1.027984e-20, -5.139921e-21, -1.541976e-20, 
    0, 1.003089e-36, -5.139921e-21, 5.139921e-21, -7.709882e-21, 
    7.709882e-21, 2.569961e-21, -5.139921e-21, 5.139921e-21, 1.027984e-20, 
    1.798972e-20, 1.798972e-20, -2.569961e-21, 1.541976e-20, 5.139921e-21, 
    -7.709882e-21, -2.569961e-21, 2.569961e-21, -1.003089e-36, -2.569961e-21, 
    -1.003089e-36, -1.541976e-20, 0, -5.139921e-21, 2.569961e-21, 
    7.709882e-21, 2.569961e-21, 1.027984e-20, 7.709882e-21, 1.28498e-20, 
    -2.569961e-21, -5.139921e-21, 1.003089e-36, 2.569961e-21, 2.569961e-21, 
    2.055969e-20, 2.569961e-21, 1.027984e-20, -2.055969e-20, 5.139921e-21, 0, 
    0, -1.027984e-20, -5.139921e-21, -1.798972e-20, 2.569961e-21, 
    -1.28498e-20, 5.139921e-21, -7.709882e-21, -1.027984e-20, -2.569961e-21, 
    -2.569961e-21, -5.139921e-21, 5.139921e-21, -7.709882e-21, -1.027984e-20, 
    -5.139921e-21, -5.139921e-21, -5.139921e-21, 2.569961e-21, -1.027984e-20, 
    1.28498e-20, -5.139921e-21, 0, 2.569961e-21, 2.569961e-21, 1.027984e-20, 
    7.709882e-21, 1.003089e-36, -7.709882e-21, -7.709882e-21, 5.139921e-21, 
    1.027984e-20, 5.139921e-21, -5.139921e-21, -1.027984e-20, 1.027984e-20, 
    0, -2.569961e-21, 7.709882e-21, -1.027984e-20, 5.139921e-21, 
    5.139921e-21, 1.003089e-36, -2.569961e-21, -2.569961e-21, -5.139921e-21, 
    7.709882e-21, -5.139921e-21, -5.139921e-21, 2.569961e-21, -5.139921e-21, 
    -2.569961e-21, -5.139921e-21, 1.027984e-20, 0, -7.709882e-21, 
    1.003089e-36, -2.569961e-21, -2.569961e-21, 2.569961e-21, -2.569961e-21, 
    1.027984e-20, 7.709882e-21, -2.569961e-21, 5.139921e-21, 5.139921e-21, 
    1.28498e-20, -2.569961e-21, 7.709882e-21, -5.139921e-21, 5.139921e-21, 
    5.139921e-21, -1.003089e-36, -7.709882e-21, -1.027984e-20, -5.139921e-21, 
    5.139921e-21, -1.28498e-20, 2.569961e-21, 7.709882e-21, -1.798972e-20, 
    1.28498e-20, 5.139921e-21, 7.709882e-21, -1.027984e-20, -2.569961e-21, 
    -2.569961e-21, -1.541976e-20, -1.541976e-20, -2.569961e-21, 5.139921e-21, 
    7.709882e-21, 2.569961e-21, 0, 5.139921e-21, 7.709882e-21, 1.027984e-20, 
    -1.28498e-20, -1.28498e-20, 1.28498e-20, -2.569961e-21, 1.027984e-20, 
    5.139921e-21, 7.709882e-21, 7.709882e-21, 2.569961e-21, 2.569961e-21, 
    -5.139921e-21, -1.003089e-36, 5.139921e-21, 2.569961e-21, -5.139921e-21, 
    -7.709882e-21, 5.139921e-21, -5.139921e-21, -5.139921e-21, 5.139921e-21, 
    5.139921e-21, 1.541976e-20, 5.139921e-21, -5.139921e-21, -7.709882e-21, 
    0, 1.28498e-20, -7.709882e-21, 5.139921e-21, 7.709882e-21, -7.709882e-21, 
    0, -2.569961e-21, 1.541976e-20, 0, 7.709882e-21, 5.139921e-21, 
    -2.569961e-21, -1.027984e-20, -1.027984e-20, -1.28498e-20, -2.569961e-21, 
    -2.569961e-21, -7.709882e-21, -1.798972e-20, -5.139921e-21, 
    -1.541976e-20, -7.709882e-21, -1.003089e-36, -2.569961e-21, 
    -2.569961e-21, -7.709882e-21, 0, -2.569961e-21, 2.312965e-20, 
    -1.027984e-20, 0, 2.569961e-21, 2.569961e-21, 0, 0, -1.003089e-36, 
    5.139921e-21, 5.139921e-21, 1.027984e-20, 0, 2.569961e-21, 0, 
    -5.139921e-21, 1.003089e-36, 7.709882e-21, 5.139921e-21, -1.027984e-20, 
    0, -2.569961e-21, -2.569961e-21, 0, -5.139921e-21, -1.28498e-20, 
    -2.569961e-21, -5.139921e-21, -1.027984e-20, 1.28498e-20, -2.055969e-20, 
    1.027984e-20, 2.569961e-21, -2.569961e-21, 7.709882e-21, -2.569961e-21, 
    -1.027984e-20, 5.139921e-21, -5.139921e-21, -1.027984e-20, 1.027984e-20, 
    -2.569961e-21, 2.055969e-20, 1.28498e-20, -2.055969e-20, -5.139921e-21, 
    1.027984e-20, 1.027984e-20, 2.569961e-21, -7.709882e-21, -7.709882e-21, 
    -1.027984e-20, 2.569961e-21, 1.027984e-20, 5.139921e-21, -1.28498e-20, 0, 
    1.027984e-20, 2.569961e-21, -1.541976e-20, -1.027984e-20, -2.569961e-21, 
    -7.709882e-21, -7.709882e-21, -5.139921e-21, -5.139921e-21, 
    -5.139921e-21, -1.027984e-20, -5.139921e-21, -5.139921e-21, 0, 
    -1.003089e-36, 1.027984e-20, 7.709882e-21, -2.569961e-21, -1.027984e-20, 
    2.569961e-21, 7.709882e-21, -1.003089e-36, 0, -2.569961e-21, 
    -5.139921e-21, 5.139921e-21, -2.569961e-21, 1.003089e-36, 5.139921e-21, 
    1.027984e-20, 2.569961e-21, 0, 0, 1.28498e-20, -7.709882e-21, 
    2.569961e-21, 7.709882e-21, 1.28498e-20,
  2.569961e-21, -5.139921e-21, 2.569961e-21, 5.139921e-21, 2.569961e-21, 
    -1.027984e-20, 5.139921e-21, -1.798972e-20, 5.139921e-21, 2.569961e-21, 
    5.139921e-21, 1.798972e-20, 7.709882e-21, -1.28498e-20, 1.027984e-20, 
    2.055969e-20, 1.027984e-20, -7.709882e-21, 2.569961e-21, 1.027984e-20, 
    -1.027984e-20, 2.055969e-20, -7.709882e-21, 7.709882e-21, -5.139921e-21, 
    1.541976e-20, -1.027984e-20, 5.139921e-21, -1.003089e-36, 1.798972e-20, 
    0, 5.139921e-21, 2.569961e-21, -1.798972e-20, -1.798972e-20, 
    1.027984e-20, -5.139921e-21, 1.027984e-20, -1.28498e-20, -5.139921e-21, 
    -5.139921e-21, -2.569961e-21, 0, 2.569961e-21, -7.709882e-21, 
    -2.569961e-21, 5.139921e-21, -1.027984e-20, -2.569961e-21, -5.139921e-21, 
    2.569961e-21, 1.027984e-20, 2.569961e-21, 7.709882e-21, 1.003089e-36, 
    -1.28498e-20, 2.569961e-21, -2.569961e-21, -1.28498e-20, -2.569961e-21, 
    1.003089e-36, -5.139921e-21, -5.139921e-21, -1.027984e-20, -5.139921e-21, 
    -5.139921e-21, -7.709882e-21, -7.709882e-21, 5.139921e-21, 2.569961e-21, 
    -1.28498e-20, 5.139921e-21, 1.027984e-20, 7.709882e-21, -1.28498e-20, 
    1.027984e-20, -7.709882e-21, 1.003089e-36, 1.798972e-20, 1.027984e-20, 
    2.569961e-21, 7.709882e-21, -2.569961e-21, 5.139921e-21, 1.28498e-20, 
    2.312965e-20, 7.709882e-21, 1.28498e-20, 5.139921e-21, -1.28498e-20, 
    -7.709882e-21, -5.139921e-21, 2.569961e-21, 1.28498e-20, 0, 2.569961e-21, 
    -5.139921e-21, -5.139921e-21, -5.139921e-21, 7.709882e-21, 1.003089e-36, 
    -1.28498e-20, 1.003089e-36, -1.541976e-20, 2.569961e-21, 0, 0, 
    -2.569961e-21, -2.569961e-21, 1.003089e-36, 1.003089e-36, -2.569961e-21, 
    -1.027984e-20, 1.027984e-20, -5.139921e-21, 2.569961e-21, 1.003089e-36, 
    1.28498e-20, 7.709882e-21, 0, -2.569961e-21, -2.569961e-21, 
    -2.312965e-20, -1.28498e-20, 1.28498e-20, 0, 1.798972e-20, 2.569961e-21, 
    1.541976e-20, 1.798972e-20, -7.709882e-21, 2.569961e-21, 1.541976e-20, 
    -5.139921e-21, 1.28498e-20, -5.139921e-21, 1.027984e-20, 2.569961e-21, 
    -1.28498e-20, -5.139921e-21, -2.569961e-21, -2.569961e-21, 5.139921e-21, 
    2.569961e-21, -2.055969e-20, -5.139921e-21, 7.709882e-21, 1.027984e-20, 
    -1.798972e-20, 0, -1.027984e-20, -1.003089e-36, -5.139921e-21, 
    -2.569961e-21, -7.709882e-21, 7.709882e-21, -7.709882e-21, 1.798972e-20, 
    -1.541976e-20, 1.541976e-20, -2.569961e-20, 1.027984e-20, 7.709882e-21, 
    2.569961e-21, -5.139921e-21, 0, -2.569961e-21, 2.569961e-21, 
    1.003089e-36, -2.826957e-20, -2.569961e-21, -2.569961e-21, -2.569961e-21, 
    1.541976e-20, 1.28498e-20, 7.709882e-21, 2.055969e-20, -1.541976e-20, 
    -7.709882e-21, -5.139921e-21, -2.569961e-21, -2.569961e-21, 7.709882e-21, 
    1.28498e-20, -5.139921e-21, 1.027984e-20, 1.027984e-20, -5.139921e-21, 
    -1.798972e-20, 1.798972e-20, -2.569961e-21, 2.569961e-21, -2.312965e-20, 
    -1.003089e-36, -7.709882e-21, -7.709882e-21, -7.709882e-21, 
    -2.569961e-21, 1.003089e-36, 5.139921e-21, -5.139921e-21, -1.541976e-20, 
    -5.139921e-21, 1.28498e-20, -2.569961e-21, -5.139921e-21, 1.027984e-20, 
    2.569961e-21, -1.027984e-20, -1.027984e-20, -5.139921e-21, -1.027984e-20, 
    -2.569961e-21, -5.139921e-21, 1.027984e-20, -2.569961e-21, 2.569961e-20, 
    2.569961e-21, 1.027984e-20, -2.569961e-21, 5.139921e-21, 1.798972e-20, 
    -1.28498e-20, 0, -1.003089e-36, -2.569961e-21, -1.541976e-20, 
    1.541976e-20, -5.139921e-21, 7.709882e-21, 2.569961e-21, 1.28498e-20, 
    -7.709882e-21, 2.569961e-21, -1.798972e-20, 1.541976e-20, -5.139921e-21, 
    5.139921e-21, -1.798972e-20, -5.139921e-21, -1.28498e-20, 1.027984e-20, 
    -5.139921e-21, 1.541976e-20, -2.569961e-21, -5.139921e-21, 7.709882e-21, 
    -5.139921e-21, -2.569961e-21, 5.139921e-21, 5.139921e-21, 1.027984e-20, 
    -7.709882e-21, 2.569961e-21, 2.569961e-21, -7.709882e-21, -1.003089e-36, 
    -1.28498e-20, -7.709882e-21, 0, 2.055969e-20, -2.569961e-21, 1.28498e-20, 
    -1.027984e-20, 1.798972e-20, 1.003089e-36, -5.139921e-21, 5.139921e-21, 
    5.139921e-21, -5.139921e-21, -5.139921e-21, 1.798972e-20, -7.709882e-21, 
    1.027984e-20, -7.709882e-21, 5.139921e-21, -2.569961e-21, 1.541976e-20, 
    1.28498e-20, 2.055969e-20, -7.709882e-21, -5.139921e-21, 5.139921e-21, 
    1.027984e-20, 1.541976e-20, 7.709882e-21, 1.541976e-20, -7.709882e-21, 
    -1.027984e-20, 7.709882e-21, 5.139921e-21, 1.003089e-36, -1.027984e-20, 
    -2.569961e-21, 1.027984e-20, -5.139921e-21, 1.541976e-20, -5.139921e-21, 
    -1.28498e-20, -2.569961e-21, -1.027984e-20, -1.798972e-20, 2.569961e-21, 
    1.541976e-20, -1.027984e-20, 7.709882e-21, 0, -7.709882e-21, 
    7.709882e-21, -5.139921e-21, -1.027984e-20, -2.569961e-21, 2.569961e-21, 
    -2.569961e-21, -7.709882e-21, -7.709882e-21, 1.28498e-20, -1.027984e-20, 
    7.709882e-21, 1.28498e-20, -7.709882e-21, -1.003089e-36, -7.709882e-21, 
    -1.027984e-20, -7.709882e-21, 5.139921e-21, -7.709882e-21, -5.139921e-21, 
    -5.139921e-21, -1.28498e-20, -1.798972e-20, -5.139921e-21, -1.798972e-20, 
    5.139921e-21, 2.569961e-21, -1.541976e-20, 5.139921e-21, 7.709882e-21,
  5.139921e-21, -7.709882e-21, 1.027984e-20, -5.139921e-21, -2.569961e-21, 
    -1.027984e-20, -7.709882e-21, 1.28498e-20, 1.027984e-20, 2.569961e-21, 
    -1.027984e-20, 1.027984e-20, 7.709882e-21, -7.709882e-21, 5.139921e-21, 
    1.798972e-20, 2.569961e-21, 2.569961e-21, -1.541976e-20, 7.709882e-21, 
    5.139921e-21, -7.709882e-21, -2.569961e-21, -2.569961e-21, -1.003089e-36, 
    1.027984e-20, 2.569961e-21, -5.139921e-21, -2.569961e-21, 1.798972e-20, 
    1.003089e-36, 1.003089e-36, 1.003089e-36, -7.709882e-21, 5.139921e-21, 
    5.139921e-21, 7.709882e-21, -2.569961e-21, -5.139921e-21, 7.709882e-21, 
    5.139921e-21, -7.709882e-21, -7.709882e-21, -2.055969e-20, 1.28498e-20, 
    -1.28498e-20, 1.027984e-20, 5.139921e-21, 2.569961e-21, -1.027984e-20, 
    -2.055969e-20, 5.139921e-21, 2.569961e-20, -1.798972e-20, 1.28498e-20, 
    1.28498e-20, 2.569961e-21, 7.709882e-21, 1.798972e-20, -1.027984e-20, 
    7.709882e-21, -5.139921e-21, 1.28498e-20, 1.027984e-20, 5.139921e-21, 
    -7.709882e-21, -2.569961e-21, 1.541976e-20, -5.139921e-21, -5.139921e-21, 
    2.569961e-21, 2.569961e-21, -5.139921e-21, 2.569961e-21, -2.055969e-20, 
    2.569961e-21, 2.569961e-21, 7.709882e-21, -7.709882e-21, 5.139921e-21, 
    7.709882e-21, 5.139921e-21, -1.28498e-20, 5.139921e-21, -2.055969e-20, 0, 
    1.798972e-20, -7.709882e-21, -7.709882e-21, -1.027984e-20, 1.541976e-20, 
    -2.569961e-21, 1.027984e-20, 2.569961e-21, 2.569961e-21, -1.28498e-20, 0, 
    7.709882e-21, -1.28498e-20, 7.709882e-21, 1.28498e-20, 1.027984e-20, 
    5.139921e-21, 7.709882e-21, 0, -1.28498e-20, -1.027984e-20, 1.28498e-20, 
    1.798972e-20, -1.28498e-20, 5.139921e-21, 1.28498e-20, -5.139921e-21, 
    2.569961e-21, 5.139921e-21, 1.003089e-36, 7.709882e-21, -1.003089e-36, 
    1.541976e-20, -5.139921e-21, -1.003089e-36, -2.569961e-21, -2.569961e-21, 
    -2.569961e-21, -1.541976e-20, 2.569961e-21, 1.28498e-20, 2.055969e-20, 
    -1.28498e-20, -2.569961e-21, 1.003089e-36, 5.139921e-21, -2.569961e-21, 
    -7.709882e-21, 7.709882e-21, 7.709882e-21, -7.709882e-21, -5.139921e-21, 
    2.569961e-21, 2.569961e-21, -2.312965e-20, 1.541976e-20, 1.027984e-20, 
    1.027984e-20, 5.139921e-21, -2.569961e-21, -2.569961e-21, -1.027984e-20, 
    -2.569961e-21, 1.541976e-20, -7.709882e-21, -1.798972e-20, 7.709882e-21, 
    -5.139921e-21, -5.139921e-21, 5.139921e-21, 2.569961e-21, -7.709882e-21, 
    5.139921e-21, -7.709882e-21, 1.027984e-20, -1.541976e-20, 1.28498e-20, 
    2.312965e-20, -2.312965e-20, 1.28498e-20, -5.139921e-21, -5.139921e-21, 
    -1.541976e-20, 0, -1.541976e-20, 2.312965e-20, -2.569961e-21, 
    -1.003089e-36, -2.055969e-20, 2.569961e-20, -1.28498e-20, -2.569961e-21, 
    -2.569961e-20, -1.027984e-20, -7.709882e-21, 2.055969e-20, 2.569961e-21, 
    1.027984e-20, 1.027984e-20, 1.027984e-20, -7.709882e-21, 1.027984e-20, 
    7.709882e-21, -2.569961e-21, -5.139921e-21, -2.569961e-21, -1.541976e-20, 
    2.055969e-20, 5.139921e-21, -7.709882e-21, 0, 5.139921e-21, -1.28498e-20, 
    -1.027984e-20, -1.003089e-36, 0, -7.709882e-21, 0, -2.569961e-21, 
    -2.569961e-21, -1.28498e-20, -1.027984e-20, 7.709882e-21, -1.541976e-20, 
    5.139921e-21, 5.139921e-21, 0, -2.569961e-21, 1.027984e-20, 
    -1.003089e-36, -1.798972e-20, 2.055969e-20, -1.027984e-20, 5.139921e-21, 
    2.569961e-21, 1.28498e-20, 7.709882e-21, 7.709882e-21, 5.139921e-21, 
    1.003089e-36, 1.28498e-20, 1.027984e-20, 2.569961e-21, 2.569961e-21, 
    -7.709882e-21, -1.027984e-20, -1.003089e-36, 5.139921e-21, 0, 
    2.569961e-21, 5.139921e-21, 0, -2.569961e-21, -5.139921e-21, 
    1.541976e-20, 1.027984e-20, 1.027984e-20, -1.28498e-20, 2.055969e-20, 
    1.003089e-36, 1.003089e-36, 1.027984e-20, 1.027984e-20, 1.28498e-20, 
    1.28498e-20, 1.003089e-36, 2.569961e-21, 1.541976e-20, 1.003089e-36, 
    -2.055969e-20, 2.569961e-21, 1.28498e-20, -5.139921e-21, -1.027984e-20, 
    -2.569961e-21, 5.139921e-21, -1.28498e-20, 2.569961e-21, 2.569961e-21, 
    1.28498e-20, 5.139921e-21, 1.027984e-20, -2.569961e-21, -2.569961e-21, 
    1.541976e-20, -1.003089e-36, -2.569961e-21, -2.569961e-21, 5.139921e-21, 
    -5.139921e-21, -2.826957e-20, -2.055969e-20, -1.003089e-36, 
    -7.709882e-21, 5.139921e-21, 5.139921e-21, -1.28498e-20, -2.569961e-21, 
    1.027984e-20, 1.027984e-20, 1.027984e-20, 2.055969e-20, -2.569961e-21, 
    2.569961e-21, 1.027984e-20, 0, 2.569961e-21, -1.003089e-36, 
    -5.139921e-21, -5.139921e-21, 7.709882e-21, -1.027984e-20, 2.055969e-20, 
    1.28498e-20, 1.003089e-36, -7.709882e-21, 5.139921e-21, -2.055969e-20, 
    2.569961e-21, 1.28498e-20, -2.569961e-21, -2.569961e-21, -5.139921e-21, 
    2.569961e-21, -5.139921e-21, -1.027984e-20, -2.569961e-21, 1.003089e-36, 
    -2.569961e-21, -2.569961e-21, -7.709882e-21, -2.312965e-20, 
    -2.569961e-21, -7.709882e-21, -2.569961e-21, -1.541976e-20, 
    -2.569961e-21, 1.027984e-20, 1.027984e-20, -7.709882e-21, 1.28498e-20, 
    -1.28498e-20, -7.709882e-21, -7.709882e-21, 2.569961e-21, 5.139921e-21, 
    -5.139921e-21, -1.003089e-36, -2.569961e-21, -1.027984e-20, 1.027984e-20, 
    -1.003089e-36,
  6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 
    6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 
    6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258065e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258065e-29, 
    6.258065e-29, 6.258065e-29, 6.258065e-29, 6.258066e-29, 6.258065e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 6.258066e-29, 
    6.258066e-29, 6.258066e-29, 6.258066e-29,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3N_TO_SOIL1N =
  5.14982e-12, 5.172541e-12, 5.168124e-12, 5.186451e-12, 5.176285e-12, 
    5.188285e-12, 5.154427e-12, 5.173443e-12, 5.161304e-12, 5.151866e-12, 
    5.222016e-12, 5.187269e-12, 5.258119e-12, 5.235955e-12, 5.291636e-12, 
    5.25467e-12, 5.299091e-12, 5.290571e-12, 5.316218e-12, 5.308871e-12, 
    5.341672e-12, 5.319609e-12, 5.358679e-12, 5.336404e-12, 5.339888e-12, 
    5.318881e-12, 5.194262e-12, 5.21769e-12, 5.192874e-12, 5.196215e-12, 
    5.194716e-12, 5.176495e-12, 5.167311e-12, 5.148084e-12, 5.151575e-12, 
    5.165697e-12, 5.197717e-12, 5.186848e-12, 5.214243e-12, 5.213624e-12, 
    5.244124e-12, 5.230372e-12, 5.281639e-12, 5.267068e-12, 5.309177e-12, 
    5.298587e-12, 5.308679e-12, 5.305619e-12, 5.308719e-12, 5.293187e-12, 
    5.299842e-12, 5.286175e-12, 5.232947e-12, 5.248589e-12, 5.201938e-12, 
    5.173888e-12, 5.15526e-12, 5.142042e-12, 5.14391e-12, 5.147473e-12, 
    5.16578e-12, 5.182994e-12, 5.196113e-12, 5.204889e-12, 5.213535e-12, 
    5.239707e-12, 5.253562e-12, 5.284585e-12, 5.278987e-12, 5.288471e-12, 
    5.297533e-12, 5.312746e-12, 5.310242e-12, 5.316945e-12, 5.288222e-12, 
    5.307311e-12, 5.275798e-12, 5.284417e-12, 5.215882e-12, 5.18978e-12, 
    5.178683e-12, 5.168973e-12, 5.145347e-12, 5.161662e-12, 5.155231e-12, 
    5.170533e-12, 5.180256e-12, 5.175448e-12, 5.205128e-12, 5.193589e-12, 
    5.254383e-12, 5.228196e-12, 5.296476e-12, 5.280136e-12, 5.300393e-12, 
    5.290057e-12, 5.307767e-12, 5.291828e-12, 5.319439e-12, 5.325452e-12, 
    5.321343e-12, 5.337127e-12, 5.290944e-12, 5.308679e-12, 5.175313e-12, 
    5.176097e-12, 5.179751e-12, 5.163688e-12, 5.162706e-12, 5.147988e-12, 
    5.161085e-12, 5.166661e-12, 5.18082e-12, 5.189195e-12, 5.197156e-12, 
    5.214661e-12, 5.234211e-12, 5.261551e-12, 5.281195e-12, 5.294363e-12, 
    5.286289e-12, 5.293418e-12, 5.285449e-12, 5.281714e-12, 5.323198e-12, 
    5.299904e-12, 5.334857e-12, 5.332923e-12, 5.317104e-12, 5.333141e-12, 
    5.176648e-12, 5.172134e-12, 5.156464e-12, 5.168727e-12, 5.146385e-12, 
    5.158891e-12, 5.166081e-12, 5.193829e-12, 5.199927e-12, 5.20558e-12, 
    5.216746e-12, 5.231076e-12, 5.256215e-12, 5.27809e-12, 5.29806e-12, 
    5.296597e-12, 5.297112e-12, 5.301573e-12, 5.290523e-12, 5.303388e-12, 
    5.305546e-12, 5.299901e-12, 5.332664e-12, 5.323304e-12, 5.332882e-12, 
    5.326788e-12, 5.173602e-12, 5.181196e-12, 5.177092e-12, 5.184809e-12, 
    5.179372e-12, 5.203546e-12, 5.210794e-12, 5.244713e-12, 5.230793e-12, 
    5.252948e-12, 5.233044e-12, 5.236571e-12, 5.253669e-12, 5.23412e-12, 
    5.276883e-12, 5.247889e-12, 5.301746e-12, 5.27279e-12, 5.303561e-12, 
    5.297974e-12, 5.307225e-12, 5.31551e-12, 5.325935e-12, 5.345168e-12, 
    5.340714e-12, 5.3568e-12, 5.192518e-12, 5.202368e-12, 5.201502e-12, 
    5.211811e-12, 5.219435e-12, 5.235961e-12, 5.262468e-12, 5.2525e-12, 
    5.2708e-12, 5.274474e-12, 5.246672e-12, 5.263741e-12, 5.208961e-12, 
    5.21781e-12, 5.212542e-12, 5.193295e-12, 5.254796e-12, 5.223232e-12, 
    5.28152e-12, 5.264419e-12, 5.314329e-12, 5.289506e-12, 5.338262e-12, 
    5.359105e-12, 5.378725e-12, 5.401651e-12, 5.207745e-12, 5.201052e-12, 
    5.213037e-12, 5.229618e-12, 5.245005e-12, 5.265462e-12, 5.267555e-12, 
    5.271388e-12, 5.281316e-12, 5.289662e-12, 5.272599e-12, 5.291755e-12, 
    5.219861e-12, 5.257536e-12, 5.19852e-12, 5.21629e-12, 5.228641e-12, 
    5.223223e-12, 5.251361e-12, 5.257993e-12, 5.284942e-12, 5.271011e-12, 
    5.35396e-12, 5.317259e-12, 5.41911e-12, 5.390645e-12, 5.198713e-12, 
    5.207722e-12, 5.239078e-12, 5.224159e-12, 5.266828e-12, 5.277332e-12, 
    5.285871e-12, 5.296786e-12, 5.297965e-12, 5.304432e-12, 5.293834e-12, 
    5.304014e-12, 5.265505e-12, 5.282714e-12, 5.235494e-12, 5.246986e-12, 
    5.2417e-12, 5.235901e-12, 5.253799e-12, 5.272867e-12, 5.273276e-12, 
    5.27939e-12, 5.296618e-12, 5.267001e-12, 5.358694e-12, 5.302063e-12, 
    5.217546e-12, 5.234899e-12, 5.237379e-12, 5.230657e-12, 5.276279e-12, 
    5.259747e-12, 5.304274e-12, 5.29224e-12, 5.311959e-12, 5.30216e-12, 
    5.300718e-12, 5.288134e-12, 5.280299e-12, 5.260505e-12, 5.244401e-12, 
    5.231632e-12, 5.234601e-12, 5.248627e-12, 5.274034e-12, 5.298071e-12, 
    5.292805e-12, 5.31046e-12, 5.263734e-12, 5.283326e-12, 5.275753e-12, 
    5.295499e-12, 5.252235e-12, 5.289073e-12, 5.242819e-12, 5.246875e-12, 
    5.259419e-12, 5.284654e-12, 5.290239e-12, 5.2962e-12, 5.292522e-12, 
    5.274679e-12, 5.271757e-12, 5.259115e-12, 5.255624e-12, 5.245992e-12, 
    5.238017e-12, 5.245302e-12, 5.252954e-12, 5.274687e-12, 5.294273e-12, 
    5.315628e-12, 5.320855e-12, 5.345804e-12, 5.325493e-12, 5.35901e-12, 
    5.330511e-12, 5.379846e-12, 5.29121e-12, 5.329675e-12, 5.25999e-12, 
    5.267497e-12, 5.281075e-12, 5.312219e-12, 5.295406e-12, 5.31507e-12, 
    5.271642e-12, 5.249111e-12, 5.243283e-12, 5.232408e-12, 5.243532e-12, 
    5.242627e-12, 5.253272e-12, 5.249851e-12, 5.275409e-12, 5.26168e-12, 
    5.300682e-12, 5.314915e-12, 5.355114e-12, 5.379758e-12, 5.404848e-12, 
    5.415924e-12, 5.419296e-12, 5.420705e-12 ;

 SOIL3N_vr =
  1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 1.818188, 1.818189, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818188, 1.818189, 1.818189, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818189, 
    1.818188, 1.818189, 1.818188, 1.818189, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818189, 1.818189, 1.818189, 1.818189, 
    1.818189, 1.818189,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 1.818188, 
    1.818188, 1.818188,
  1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 1.818187, 
    1.818187, 1.818187,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOIL3_HR =
  3.115641e-11, 3.129387e-11, 3.126715e-11, 3.137803e-11, 3.131653e-11, 
    3.138912e-11, 3.118428e-11, 3.129933e-11, 3.122589e-11, 3.116879e-11, 
    3.15932e-11, 3.138298e-11, 3.181162e-11, 3.167753e-11, 3.20144e-11, 
    3.179075e-11, 3.20595e-11, 3.200796e-11, 3.216312e-11, 3.211867e-11, 
    3.231712e-11, 3.218363e-11, 3.242001e-11, 3.228524e-11, 3.230632e-11, 
    3.217923e-11, 3.142529e-11, 3.156702e-11, 3.141689e-11, 3.14371e-11, 
    3.142803e-11, 3.131779e-11, 3.126224e-11, 3.114591e-11, 3.116703e-11, 
    3.125247e-11, 3.144619e-11, 3.138043e-11, 3.154617e-11, 3.154243e-11, 
    3.172695e-11, 3.164375e-11, 3.195392e-11, 3.186576e-11, 3.212052e-11, 
    3.205645e-11, 3.211751e-11, 3.2099e-11, 3.211775e-11, 3.202378e-11, 
    3.206404e-11, 3.198136e-11, 3.165933e-11, 3.175396e-11, 3.147172e-11, 
    3.130202e-11, 3.118933e-11, 3.110935e-11, 3.112066e-11, 3.114221e-11, 
    3.125297e-11, 3.135711e-11, 3.143649e-11, 3.148957e-11, 3.154189e-11, 
    3.170023e-11, 3.178405e-11, 3.197174e-11, 3.193787e-11, 3.199525e-11, 
    3.205007e-11, 3.214212e-11, 3.212697e-11, 3.216752e-11, 3.199374e-11, 
    3.210923e-11, 3.191858e-11, 3.197072e-11, 3.155608e-11, 3.139817e-11, 
    3.133103e-11, 3.127229e-11, 3.112935e-11, 3.122806e-11, 3.118915e-11, 
    3.128173e-11, 3.134055e-11, 3.131146e-11, 3.149103e-11, 3.142121e-11, 
    3.178902e-11, 3.163059e-11, 3.204368e-11, 3.194483e-11, 3.206738e-11, 
    3.200484e-11, 3.211199e-11, 3.201556e-11, 3.218261e-11, 3.221898e-11, 
    3.219413e-11, 3.228962e-11, 3.201021e-11, 3.211751e-11, 3.131064e-11, 
    3.131539e-11, 3.13375e-11, 3.124032e-11, 3.123437e-11, 3.114533e-11, 
    3.122456e-11, 3.12583e-11, 3.134396e-11, 3.139463e-11, 3.14428e-11, 
    3.15487e-11, 3.166698e-11, 3.183238e-11, 3.195123e-11, 3.20309e-11, 
    3.198205e-11, 3.202517e-11, 3.197696e-11, 3.195437e-11, 3.220535e-11, 
    3.206442e-11, 3.227589e-11, 3.226418e-11, 3.216848e-11, 3.22655e-11, 
    3.131872e-11, 3.129141e-11, 3.119661e-11, 3.12708e-11, 3.113563e-11, 
    3.121129e-11, 3.125479e-11, 3.142267e-11, 3.145956e-11, 3.149376e-11, 
    3.156131e-11, 3.164801e-11, 3.18001e-11, 3.193244e-11, 3.205327e-11, 
    3.204441e-11, 3.204753e-11, 3.207452e-11, 3.200766e-11, 3.208549e-11, 
    3.209856e-11, 3.20644e-11, 3.226262e-11, 3.220599e-11, 3.226394e-11, 
    3.222706e-11, 3.130029e-11, 3.134623e-11, 3.132141e-11, 3.136809e-11, 
    3.13352e-11, 3.148145e-11, 3.152531e-11, 3.173051e-11, 3.16463e-11, 
    3.178034e-11, 3.165992e-11, 3.168125e-11, 3.17847e-11, 3.166643e-11, 
    3.192514e-11, 3.174973e-11, 3.207557e-11, 3.190038e-11, 3.208655e-11, 
    3.205274e-11, 3.210871e-11, 3.215884e-11, 3.22219e-11, 3.233826e-11, 
    3.231132e-11, 3.240864e-11, 3.141473e-11, 3.147433e-11, 3.146908e-11, 
    3.153145e-11, 3.157758e-11, 3.167756e-11, 3.183793e-11, 3.177763e-11, 
    3.188834e-11, 3.191056e-11, 3.174237e-11, 3.184563e-11, 3.151421e-11, 
    3.156775e-11, 3.153588e-11, 3.141943e-11, 3.179151e-11, 3.160055e-11, 
    3.195319e-11, 3.184974e-11, 3.215169e-11, 3.200151e-11, 3.229649e-11, 
    3.242258e-11, 3.254129e-11, 3.267999e-11, 3.150686e-11, 3.146636e-11, 
    3.153887e-11, 3.163919e-11, 3.173228e-11, 3.185605e-11, 3.186871e-11, 
    3.18919e-11, 3.195196e-11, 3.200246e-11, 3.189922e-11, 3.201512e-11, 
    3.158016e-11, 3.180809e-11, 3.145105e-11, 3.155855e-11, 3.163328e-11, 
    3.16005e-11, 3.177074e-11, 3.181086e-11, 3.19739e-11, 3.188962e-11, 
    3.239146e-11, 3.216942e-11, 3.278562e-11, 3.26134e-11, 3.145221e-11, 
    3.150672e-11, 3.169642e-11, 3.160616e-11, 3.186431e-11, 3.192786e-11, 
    3.197952e-11, 3.204555e-11, 3.205269e-11, 3.209181e-11, 3.20277e-11, 
    3.208928e-11, 3.185631e-11, 3.196042e-11, 3.167474e-11, 3.174427e-11, 
    3.171229e-11, 3.16772e-11, 3.178548e-11, 3.190085e-11, 3.190332e-11, 
    3.194031e-11, 3.204454e-11, 3.186536e-11, 3.24201e-11, 3.207748e-11, 
    3.156616e-11, 3.167114e-11, 3.168614e-11, 3.164547e-11, 3.192148e-11, 
    3.182147e-11, 3.209086e-11, 3.201805e-11, 3.213735e-11, 3.207807e-11, 
    3.206935e-11, 3.199321e-11, 3.194581e-11, 3.182606e-11, 3.172863e-11, 
    3.165137e-11, 3.166934e-11, 3.17542e-11, 3.190791e-11, 3.205333e-11, 
    3.202147e-11, 3.212828e-11, 3.184559e-11, 3.196412e-11, 3.191831e-11, 
    3.203777e-11, 3.177602e-11, 3.199889e-11, 3.171905e-11, 3.174359e-11, 
    3.181949e-11, 3.197216e-11, 3.200595e-11, 3.204201e-11, 3.201976e-11, 
    3.191181e-11, 3.189413e-11, 3.181764e-11, 3.179652e-11, 3.173825e-11, 
    3.169e-11, 3.173408e-11, 3.178037e-11, 3.191186e-11, 3.203035e-11, 
    3.215955e-11, 3.219117e-11, 3.234212e-11, 3.221923e-11, 3.242201e-11, 
    3.224959e-11, 3.254807e-11, 3.201182e-11, 3.224453e-11, 3.182294e-11, 
    3.186836e-11, 3.19505e-11, 3.213893e-11, 3.203721e-11, 3.215617e-11, 
    3.189344e-11, 3.175712e-11, 3.172186e-11, 3.165607e-11, 3.172337e-11, 
    3.17179e-11, 3.17823e-11, 3.17616e-11, 3.191622e-11, 3.183316e-11, 
    3.206913e-11, 3.215523e-11, 3.239844e-11, 3.254753e-11, 3.269933e-11, 
    3.276634e-11, 3.278674e-11, 3.279527e-11 ;

 SOILC =
  17.34481, 17.3448, 17.3448, 17.34479, 17.34479, 17.34479, 17.34481, 
    17.3448, 17.3448, 17.34481, 17.34477, 17.34479, 17.34475, 17.34476, 
    17.34473, 17.34475, 17.34472, 17.34473, 17.34471, 17.34472, 17.3447, 
    17.34471, 17.34469, 17.3447, 17.3447, 17.34471, 17.34478, 17.34477, 
    17.34478, 17.34478, 17.34478, 17.34479, 17.3448, 17.34481, 17.34481, 
    17.3448, 17.34478, 17.34479, 17.34477, 17.34477, 17.34476, 17.34476, 
    17.34473, 17.34474, 17.34472, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34473, 17.34472, 17.34473, 17.34476, 17.34475, 17.34478, 17.3448, 
    17.34481, 17.34481, 17.34481, 17.34481, 17.3448, 17.34479, 17.34478, 
    17.34478, 17.34477, 17.34476, 17.34475, 17.34473, 17.34473, 17.34473, 
    17.34472, 17.34472, 17.34472, 17.34471, 17.34473, 17.34472, 17.34474, 
    17.34473, 17.34477, 17.34479, 17.34479, 17.3448, 17.34481, 17.3448, 
    17.34481, 17.3448, 17.34479, 17.3448, 17.34478, 17.34478, 17.34475, 
    17.34476, 17.34472, 17.34473, 17.34472, 17.34473, 17.34472, 17.34473, 
    17.34471, 17.34471, 17.34471, 17.3447, 17.34473, 17.34472, 17.3448, 
    17.34479, 17.34479, 17.3448, 17.3448, 17.34481, 17.3448, 17.3448, 
    17.34479, 17.34479, 17.34478, 17.34477, 17.34476, 17.34475, 17.34473, 
    17.34473, 17.34473, 17.34473, 17.34473, 17.34473, 17.34471, 17.34472, 
    17.3447, 17.3447, 17.34471, 17.3447, 17.34479, 17.3448, 17.3448, 17.3448, 
    17.34481, 17.3448, 17.3448, 17.34478, 17.34478, 17.34478, 17.34477, 
    17.34476, 17.34475, 17.34474, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34473, 17.34472, 17.34472, 17.34472, 17.3447, 17.34471, 17.3447, 
    17.34471, 17.3448, 17.34479, 17.34479, 17.34479, 17.34479, 17.34478, 
    17.34477, 17.34476, 17.34476, 17.34475, 17.34476, 17.34476, 17.34475, 
    17.34476, 17.34474, 17.34475, 17.34472, 17.34474, 17.34472, 17.34472, 
    17.34472, 17.34471, 17.34471, 17.3447, 17.3447, 17.34469, 17.34478, 
    17.34478, 17.34478, 17.34477, 17.34477, 17.34476, 17.34474, 17.34475, 
    17.34474, 17.34474, 17.34475, 17.34474, 17.34477, 17.34477, 17.34477, 
    17.34478, 17.34475, 17.34477, 17.34473, 17.34474, 17.34472, 17.34473, 
    17.3447, 17.34469, 17.34468, 17.34466, 17.34478, 17.34478, 17.34477, 
    17.34476, 17.34476, 17.34474, 17.34474, 17.34474, 17.34473, 17.34473, 
    17.34474, 17.34473, 17.34477, 17.34475, 17.34478, 17.34477, 17.34476, 
    17.34477, 17.34475, 17.34475, 17.34473, 17.34474, 17.34469, 17.34471, 
    17.34465, 17.34467, 17.34478, 17.34478, 17.34476, 17.34477, 17.34474, 
    17.34474, 17.34473, 17.34472, 17.34472, 17.34472, 17.34473, 17.34472, 
    17.34474, 17.34473, 17.34476, 17.34475, 17.34476, 17.34476, 17.34475, 
    17.34474, 17.34474, 17.34473, 17.34472, 17.34474, 17.34469, 17.34472, 
    17.34477, 17.34476, 17.34476, 17.34476, 17.34474, 17.34475, 17.34472, 
    17.34473, 17.34472, 17.34472, 17.34472, 17.34473, 17.34473, 17.34475, 
    17.34476, 17.34476, 17.34476, 17.34475, 17.34474, 17.34472, 17.34473, 
    17.34472, 17.34474, 17.34473, 17.34474, 17.34472, 17.34475, 17.34473, 
    17.34476, 17.34475, 17.34475, 17.34473, 17.34473, 17.34472, 17.34473, 
    17.34474, 17.34474, 17.34475, 17.34475, 17.34475, 17.34476, 17.34475, 
    17.34475, 17.34474, 17.34473, 17.34471, 17.34471, 17.3447, 17.34471, 
    17.34469, 17.34471, 17.34468, 17.34473, 17.34471, 17.34475, 17.34474, 
    17.34473, 17.34472, 17.34472, 17.34471, 17.34474, 17.34475, 17.34476, 
    17.34476, 17.34476, 17.34476, 17.34475, 17.34475, 17.34474, 17.34475, 
    17.34472, 17.34471, 17.34469, 17.34468, 17.34466, 17.34466, 17.34465, 
    17.34465 ;

 SOILC_HR =
  6.191113e-08, 6.218415e-08, 6.213108e-08, 6.235129e-08, 6.222914e-08, 
    6.237333e-08, 6.196649e-08, 6.219499e-08, 6.204912e-08, 6.193572e-08, 
    6.277865e-08, 6.236112e-08, 6.321246e-08, 6.294614e-08, 6.361521e-08, 
    6.317101e-08, 6.370478e-08, 6.360241e-08, 6.391058e-08, 6.382229e-08, 
    6.421644e-08, 6.395133e-08, 6.44208e-08, 6.415313e-08, 6.4195e-08, 
    6.394257e-08, 6.244515e-08, 6.272666e-08, 6.242847e-08, 6.246862e-08, 
    6.24506e-08, 6.223166e-08, 6.212131e-08, 6.189027e-08, 6.193222e-08, 
    6.210192e-08, 6.248666e-08, 6.235607e-08, 6.268525e-08, 6.267781e-08, 
    6.304429e-08, 6.287905e-08, 6.349508e-08, 6.331999e-08, 6.382597e-08, 
    6.369872e-08, 6.382e-08, 6.378323e-08, 6.382047e-08, 6.363384e-08, 
    6.37138e-08, 6.354958e-08, 6.290999e-08, 6.309795e-08, 6.253738e-08, 
    6.220033e-08, 6.197651e-08, 6.181767e-08, 6.184013e-08, 6.188293e-08, 
    6.210291e-08, 6.230976e-08, 6.246739e-08, 6.257284e-08, 6.267674e-08, 
    6.299121e-08, 6.31577e-08, 6.353047e-08, 6.346321e-08, 6.357717e-08, 
    6.368606e-08, 6.386886e-08, 6.383878e-08, 6.391931e-08, 6.357418e-08, 
    6.380355e-08, 6.34249e-08, 6.352845e-08, 6.270493e-08, 6.23913e-08, 
    6.225795e-08, 6.214128e-08, 6.185739e-08, 6.205343e-08, 6.197615e-08, 
    6.216003e-08, 6.227686e-08, 6.221908e-08, 6.257572e-08, 6.243706e-08, 
    6.316757e-08, 6.285291e-08, 6.367335e-08, 6.347702e-08, 6.372042e-08, 
    6.359622e-08, 6.380903e-08, 6.361751e-08, 6.394929e-08, 6.402153e-08, 
    6.397217e-08, 6.416183e-08, 6.360688e-08, 6.381999e-08, 6.221745e-08, 
    6.222687e-08, 6.227079e-08, 6.207778e-08, 6.206597e-08, 6.188912e-08, 
    6.204649e-08, 6.21135e-08, 6.228363e-08, 6.238426e-08, 6.247993e-08, 
    6.269027e-08, 6.292518e-08, 6.32537e-08, 6.348974e-08, 6.364797e-08, 
    6.355095e-08, 6.363661e-08, 6.354085e-08, 6.349597e-08, 6.399446e-08, 
    6.371454e-08, 6.413455e-08, 6.411131e-08, 6.392123e-08, 6.411393e-08, 
    6.22335e-08, 6.217927e-08, 6.199097e-08, 6.213833e-08, 6.186986e-08, 
    6.202013e-08, 6.210653e-08, 6.243995e-08, 6.251322e-08, 6.258114e-08, 
    6.271532e-08, 6.288751e-08, 6.318957e-08, 6.345243e-08, 6.36924e-08, 
    6.367481e-08, 6.3681e-08, 6.373461e-08, 6.360182e-08, 6.375641e-08, 
    6.378234e-08, 6.371452e-08, 6.410819e-08, 6.399572e-08, 6.411081e-08, 
    6.403759e-08, 6.21969e-08, 6.228814e-08, 6.223884e-08, 6.233156e-08, 
    6.226623e-08, 6.255671e-08, 6.264381e-08, 6.305137e-08, 6.288411e-08, 
    6.315032e-08, 6.291116e-08, 6.295353e-08, 6.315899e-08, 6.292409e-08, 
    6.343792e-08, 6.308954e-08, 6.373669e-08, 6.338875e-08, 6.375849e-08, 
    6.369136e-08, 6.380252e-08, 6.390207e-08, 6.402733e-08, 6.425844e-08, 
    6.420493e-08, 6.439821e-08, 6.242419e-08, 6.254255e-08, 6.253214e-08, 
    6.265601e-08, 6.274763e-08, 6.294621e-08, 6.326471e-08, 6.314495e-08, 
    6.336484e-08, 6.340898e-08, 6.307491e-08, 6.328001e-08, 6.262177e-08, 
    6.272811e-08, 6.26648e-08, 6.243353e-08, 6.317253e-08, 6.279325e-08, 
    6.349364e-08, 6.328816e-08, 6.388787e-08, 6.358961e-08, 6.417547e-08, 
    6.44259e-08, 6.466167e-08, 6.493715e-08, 6.260716e-08, 6.252674e-08, 
    6.267075e-08, 6.286999e-08, 6.305489e-08, 6.33007e-08, 6.332585e-08, 
    6.33719e-08, 6.349119e-08, 6.359149e-08, 6.338645e-08, 6.361663e-08, 
    6.275275e-08, 6.320546e-08, 6.249633e-08, 6.270984e-08, 6.285825e-08, 
    6.279316e-08, 6.313125e-08, 6.321094e-08, 6.353477e-08, 6.336737e-08, 
    6.436409e-08, 6.392309e-08, 6.514694e-08, 6.480489e-08, 6.249864e-08, 
    6.260689e-08, 6.298366e-08, 6.280439e-08, 6.331711e-08, 6.344332e-08, 
    6.354593e-08, 6.367708e-08, 6.369125e-08, 6.376896e-08, 6.364161e-08, 
    6.376393e-08, 6.330121e-08, 6.350799e-08, 6.29406e-08, 6.307869e-08, 
    6.301516e-08, 6.294548e-08, 6.316055e-08, 6.338968e-08, 6.339459e-08, 
    6.346806e-08, 6.367506e-08, 6.331919e-08, 6.442097e-08, 6.374049e-08, 
    6.272494e-08, 6.293345e-08, 6.296325e-08, 6.288247e-08, 6.343066e-08, 
    6.323202e-08, 6.376707e-08, 6.362246e-08, 6.38594e-08, 6.374166e-08, 
    6.372434e-08, 6.357312e-08, 6.347897e-08, 6.324113e-08, 6.304762e-08, 
    6.289419e-08, 6.292986e-08, 6.309841e-08, 6.34037e-08, 6.369253e-08, 
    6.362925e-08, 6.384139e-08, 6.327993e-08, 6.351534e-08, 6.342435e-08, 
    6.366162e-08, 6.314175e-08, 6.35844e-08, 6.302862e-08, 6.307734e-08, 
    6.322809e-08, 6.35313e-08, 6.359841e-08, 6.367004e-08, 6.362585e-08, 
    6.341145e-08, 6.337633e-08, 6.322442e-08, 6.318248e-08, 6.306674e-08, 
    6.297091e-08, 6.305846e-08, 6.31504e-08, 6.341154e-08, 6.364689e-08, 
    6.390349e-08, 6.39663e-08, 6.426609e-08, 6.402202e-08, 6.442477e-08, 
    6.408233e-08, 6.467514e-08, 6.361008e-08, 6.407228e-08, 6.323495e-08, 
    6.332515e-08, 6.34883e-08, 6.386253e-08, 6.366051e-08, 6.389678e-08, 
    6.337496e-08, 6.310422e-08, 6.303419e-08, 6.290352e-08, 6.303718e-08, 
    6.302631e-08, 6.315422e-08, 6.311311e-08, 6.342022e-08, 6.325525e-08, 
    6.37239e-08, 6.389492e-08, 6.437795e-08, 6.467408e-08, 6.497555e-08, 
    6.510865e-08, 6.514917e-08, 6.51661e-08 ;

 SOILC_LOSS =
  6.191113e-08, 6.218415e-08, 6.213108e-08, 6.235129e-08, 6.222914e-08, 
    6.237333e-08, 6.196649e-08, 6.219499e-08, 6.204912e-08, 6.193572e-08, 
    6.277865e-08, 6.236112e-08, 6.321246e-08, 6.294614e-08, 6.361521e-08, 
    6.317101e-08, 6.370478e-08, 6.360241e-08, 6.391058e-08, 6.382229e-08, 
    6.421644e-08, 6.395133e-08, 6.44208e-08, 6.415313e-08, 6.4195e-08, 
    6.394257e-08, 6.244515e-08, 6.272666e-08, 6.242847e-08, 6.246862e-08, 
    6.24506e-08, 6.223166e-08, 6.212131e-08, 6.189027e-08, 6.193222e-08, 
    6.210192e-08, 6.248666e-08, 6.235607e-08, 6.268525e-08, 6.267781e-08, 
    6.304429e-08, 6.287905e-08, 6.349508e-08, 6.331999e-08, 6.382597e-08, 
    6.369872e-08, 6.382e-08, 6.378323e-08, 6.382047e-08, 6.363384e-08, 
    6.37138e-08, 6.354958e-08, 6.290999e-08, 6.309795e-08, 6.253738e-08, 
    6.220033e-08, 6.197651e-08, 6.181767e-08, 6.184013e-08, 6.188293e-08, 
    6.210291e-08, 6.230976e-08, 6.246739e-08, 6.257284e-08, 6.267674e-08, 
    6.299121e-08, 6.31577e-08, 6.353047e-08, 6.346321e-08, 6.357717e-08, 
    6.368606e-08, 6.386886e-08, 6.383878e-08, 6.391931e-08, 6.357418e-08, 
    6.380355e-08, 6.34249e-08, 6.352845e-08, 6.270493e-08, 6.23913e-08, 
    6.225795e-08, 6.214128e-08, 6.185739e-08, 6.205343e-08, 6.197615e-08, 
    6.216003e-08, 6.227686e-08, 6.221908e-08, 6.257572e-08, 6.243706e-08, 
    6.316757e-08, 6.285291e-08, 6.367335e-08, 6.347702e-08, 6.372042e-08, 
    6.359622e-08, 6.380903e-08, 6.361751e-08, 6.394929e-08, 6.402153e-08, 
    6.397217e-08, 6.416183e-08, 6.360688e-08, 6.381999e-08, 6.221745e-08, 
    6.222687e-08, 6.227079e-08, 6.207778e-08, 6.206597e-08, 6.188912e-08, 
    6.204649e-08, 6.21135e-08, 6.228363e-08, 6.238426e-08, 6.247993e-08, 
    6.269027e-08, 6.292518e-08, 6.32537e-08, 6.348974e-08, 6.364797e-08, 
    6.355095e-08, 6.363661e-08, 6.354085e-08, 6.349597e-08, 6.399446e-08, 
    6.371454e-08, 6.413455e-08, 6.411131e-08, 6.392123e-08, 6.411393e-08, 
    6.22335e-08, 6.217927e-08, 6.199097e-08, 6.213833e-08, 6.186986e-08, 
    6.202013e-08, 6.210653e-08, 6.243995e-08, 6.251322e-08, 6.258114e-08, 
    6.271532e-08, 6.288751e-08, 6.318957e-08, 6.345243e-08, 6.36924e-08, 
    6.367481e-08, 6.3681e-08, 6.373461e-08, 6.360182e-08, 6.375641e-08, 
    6.378234e-08, 6.371452e-08, 6.410819e-08, 6.399572e-08, 6.411081e-08, 
    6.403759e-08, 6.21969e-08, 6.228814e-08, 6.223884e-08, 6.233156e-08, 
    6.226623e-08, 6.255671e-08, 6.264381e-08, 6.305137e-08, 6.288411e-08, 
    6.315032e-08, 6.291116e-08, 6.295353e-08, 6.315899e-08, 6.292409e-08, 
    6.343792e-08, 6.308954e-08, 6.373669e-08, 6.338875e-08, 6.375849e-08, 
    6.369136e-08, 6.380252e-08, 6.390207e-08, 6.402733e-08, 6.425844e-08, 
    6.420493e-08, 6.439821e-08, 6.242419e-08, 6.254255e-08, 6.253214e-08, 
    6.265601e-08, 6.274763e-08, 6.294621e-08, 6.326471e-08, 6.314495e-08, 
    6.336484e-08, 6.340898e-08, 6.307491e-08, 6.328001e-08, 6.262177e-08, 
    6.272811e-08, 6.26648e-08, 6.243353e-08, 6.317253e-08, 6.279325e-08, 
    6.349364e-08, 6.328816e-08, 6.388787e-08, 6.358961e-08, 6.417547e-08, 
    6.44259e-08, 6.466167e-08, 6.493715e-08, 6.260716e-08, 6.252674e-08, 
    6.267075e-08, 6.286999e-08, 6.305489e-08, 6.33007e-08, 6.332585e-08, 
    6.33719e-08, 6.349119e-08, 6.359149e-08, 6.338645e-08, 6.361663e-08, 
    6.275275e-08, 6.320546e-08, 6.249633e-08, 6.270984e-08, 6.285825e-08, 
    6.279316e-08, 6.313125e-08, 6.321094e-08, 6.353477e-08, 6.336737e-08, 
    6.436409e-08, 6.392309e-08, 6.514694e-08, 6.480489e-08, 6.249864e-08, 
    6.260689e-08, 6.298366e-08, 6.280439e-08, 6.331711e-08, 6.344332e-08, 
    6.354593e-08, 6.367708e-08, 6.369125e-08, 6.376896e-08, 6.364161e-08, 
    6.376393e-08, 6.330121e-08, 6.350799e-08, 6.29406e-08, 6.307869e-08, 
    6.301516e-08, 6.294548e-08, 6.316055e-08, 6.338968e-08, 6.339459e-08, 
    6.346806e-08, 6.367506e-08, 6.331919e-08, 6.442097e-08, 6.374049e-08, 
    6.272494e-08, 6.293345e-08, 6.296325e-08, 6.288247e-08, 6.343066e-08, 
    6.323202e-08, 6.376707e-08, 6.362246e-08, 6.38594e-08, 6.374166e-08, 
    6.372434e-08, 6.357312e-08, 6.347897e-08, 6.324113e-08, 6.304762e-08, 
    6.289419e-08, 6.292986e-08, 6.309841e-08, 6.34037e-08, 6.369253e-08, 
    6.362925e-08, 6.384139e-08, 6.327993e-08, 6.351534e-08, 6.342435e-08, 
    6.366162e-08, 6.314175e-08, 6.35844e-08, 6.302862e-08, 6.307734e-08, 
    6.322809e-08, 6.35313e-08, 6.359841e-08, 6.367004e-08, 6.362585e-08, 
    6.341145e-08, 6.337633e-08, 6.322442e-08, 6.318248e-08, 6.306674e-08, 
    6.297091e-08, 6.305846e-08, 6.31504e-08, 6.341154e-08, 6.364689e-08, 
    6.390349e-08, 6.39663e-08, 6.426609e-08, 6.402202e-08, 6.442477e-08, 
    6.408233e-08, 6.467514e-08, 6.361008e-08, 6.407228e-08, 6.323495e-08, 
    6.332515e-08, 6.34883e-08, 6.386253e-08, 6.366051e-08, 6.389678e-08, 
    6.337496e-08, 6.310422e-08, 6.303419e-08, 6.290352e-08, 6.303718e-08, 
    6.302631e-08, 6.315422e-08, 6.311311e-08, 6.342022e-08, 6.325525e-08, 
    6.37239e-08, 6.389492e-08, 6.437795e-08, 6.467408e-08, 6.497555e-08, 
    6.510865e-08, 6.514917e-08, 6.51661e-08 ;

 SOILICE =
  95.00039, 95.4491, 95.36176, 95.7245, 95.52316, 95.76085, 95.09124, 
    95.46696, 95.22699, 95.04072, 96.4311, 95.7407, 97.15166, 96.70879, 
    97.82378, 97.08266, 97.97365, 97.80232, 98.31852, 98.17046, 98.83266, 
    98.3869, 99.17702, 98.72607, 98.79654, 98.37222, 95.87936, 96.34497, 
    95.85182, 95.91811, 95.88836, 95.52732, 95.34573, 94.96614, 95.03497, 
    95.31381, 95.94793, 95.73235, 96.27625, 96.26395, 96.87184, 96.59744, 
    97.62294, 97.33075, 98.17664, 97.96346, 98.16662, 98.10498, 98.16742, 
    97.8549, 97.98872, 97.714, 96.6488, 96.96107, 96.03172, 95.47579, 
    95.1077, 94.84708, 94.8839, 94.95411, 95.31544, 95.65599, 95.91607, 
    96.0903, 96.26218, 96.78374, 97.06049, 97.6821, 97.56971, 97.76014, 
    97.94227, 98.24856, 98.1981, 98.33319, 97.7551, 98.13906, 97.50574, 
    97.6787, 96.30901, 95.79047, 95.57069, 95.37855, 94.91222, 95.23409, 
    95.10712, 95.40937, 95.60177, 95.50658, 96.09507, 95.866, 97.07691, 
    96.5541, 97.92101, 97.59277, 97.99979, 97.79196, 98.14825, 97.82755, 
    98.3835, 98.50484, 98.42191, 98.74068, 97.8098, 98.16662, 95.50391, 
    95.51943, 95.59176, 95.27412, 95.2547, 94.96426, 95.22266, 95.33285, 
    95.61292, 95.77886, 95.93678, 96.28458, 96.67403, 97.22032, 97.61403, 
    97.87852, 97.71628, 97.85951, 97.69941, 97.62442, 98.45937, 97.98997, 
    98.69479, 98.6557, 98.33641, 98.6601, 95.53033, 95.44103, 95.13145, 
    95.37367, 94.93266, 95.17935, 95.3214, 95.87079, 95.99177, 96.10405, 
    96.32606, 96.61148, 97.11353, 97.55173, 97.95287, 97.92344, 97.9338, 
    98.02355, 97.80133, 98.06007, 98.10354, 97.98991, 98.65047, 98.46146, 
    98.65487, 98.53177, 95.47005, 95.62037, 95.53913, 95.69195, 95.58427, 
    96.06368, 96.20773, 96.88365, 96.60586, 97.04819, 96.65073, 96.72108, 
    97.06268, 96.67217, 97.52754, 96.94711, 98.02704, 97.4455, 98.06356, 
    97.95113, 98.13731, 98.30427, 98.51455, 98.90334, 98.81322, 99.1389, 
    95.84475, 96.04027, 96.02303, 96.22789, 96.37959, 96.7089, 97.23864, 
    97.03921, 97.40553, 97.47918, 96.92273, 97.26414, 96.17126, 96.34728, 
    96.24244, 95.86017, 97.08516, 96.45521, 97.62054, 97.27771, 98.28046, 
    97.78095, 98.76363, 99.18568, 99.58389, 100.0506, 96.14707, 96.0141, 
    96.25227, 96.58245, 96.88945, 97.29861, 97.34052, 97.41733, 97.61643, 
    97.78404, 97.44163, 97.8261, 96.38816, 97.13996, 95.96387, 96.31703, 
    96.56297, 96.45502, 97.01643, 97.14906, 97.68927, 97.40977, 99.08142, 
    98.33957, 100.4068, 99.82637, 95.96767, 96.14661, 96.77112, 96.47364, 
    97.32595, 97.53651, 97.70788, 97.92725, 97.95095, 98.08109, 97.86788, 
    98.07266, 97.29948, 97.6445, 96.69958, 96.92902, 96.82343, 96.70769, 
    97.06518, 97.44701, 97.45516, 97.57782, 97.92403, 97.32941, 99.17747, 
    98.03354, 96.34198, 96.68776, 96.7372, 96.60311, 97.51538, 97.18419, 
    98.07792, 97.83585, 98.23267, 98.03535, 98.00635, 97.75334, 97.59604, 
    97.19936, 96.87738, 96.62255, 96.68176, 96.96183, 97.4704, 97.9531, 
    97.84724, 98.20248, 97.26398, 97.65681, 97.50487, 97.90137, 97.03392, 
    97.77235, 96.84576, 96.92677, 97.17762, 97.68351, 97.79563, 97.91547, 
    97.84151, 97.48333, 97.42472, 97.17152, 97.10169, 96.90913, 96.74991, 
    96.89538, 97.04831, 97.48347, 97.87673, 98.30665, 98.41203, 98.91629, 
    98.50571, 99.18387, 98.60715, 99.6068, 97.81522, 98.59019, 97.18904, 
    97.33936, 97.61165, 98.23799, 97.89951, 98.29543, 97.42242, 96.97151, 
    96.85504, 96.63803, 96.86001, 96.84194, 97.05463, 96.98625, 97.49794, 
    97.22286, 98.00562, 98.29229, 99.10474, 99.60493, 100.1157, 100.3417, 
    100.4106, 100.4394,
  95.09608, 95.56266, 95.47182, 95.84899, 95.63962, 95.88678, 95.19051, 
    95.58125, 95.33168, 95.13796, 96.58361, 95.86583, 97.33221, 96.872, 
    98.0304, 97.26057, 98.18604, 98.00804, 98.54411, 98.39036, 99.07811, 
    98.61513, 99.43556, 98.96737, 99.04057, 98.59989, 96.00993, 96.4941, 
    95.98131, 96.05025, 96.01929, 95.64397, 95.45524, 95.06041, 95.132, 
    95.42199, 96.08125, 95.85709, 96.42245, 96.40965, 97.04141, 96.75626, 
    97.82172, 97.51817, 98.39677, 98.17539, 98.38638, 98.32236, 98.38721, 
    98.06265, 98.20164, 97.91629, 96.80965, 97.13414, 96.16832, 95.59051, 
    95.20765, 94.9366, 94.97489, 95.04794, 95.42369, 95.77771, 96.04807, 
    96.22918, 96.40781, 96.95, 97.2375, 97.88321, 97.76641, 97.96426, 
    98.15338, 98.47148, 98.41907, 98.55939, 97.95898, 98.3578, 97.69994, 
    97.87962, 96.45674, 95.91752, 95.68916, 95.48929, 95.00435, 95.3391, 
    95.20705, 95.5213, 95.72134, 95.62236, 96.23413, 95.99603, 97.25455, 
    96.71126, 98.13131, 97.79037, 98.21312, 97.99725, 98.36732, 98.03423, 
    98.61161, 98.73764, 98.65151, 98.98248, 98.01579, 98.38641, 95.61961, 
    95.63574, 95.71093, 95.38071, 95.36052, 95.05846, 95.32718, 95.44177, 
    95.73293, 95.90545, 96.06961, 96.43113, 96.8359, 97.4035, 97.81245, 
    98.08716, 97.91864, 98.06741, 97.90112, 97.82323, 98.69043, 98.20296, 
    98.93484, 98.89425, 98.56274, 98.89882, 95.64707, 95.55421, 95.23234, 
    95.48418, 95.0256, 95.28217, 95.4299, 96.00107, 96.12675, 96.24349, 
    96.47422, 96.77085, 97.29254, 97.74776, 98.16438, 98.1338, 98.14457, 
    98.23781, 98.007, 98.27573, 98.3209, 98.20286, 98.88881, 98.69255, 
    98.89339, 98.76556, 95.58439, 95.74068, 95.65621, 95.81511, 95.70317, 
    96.20159, 96.35133, 97.05375, 96.76502, 97.22469, 96.81163, 96.88477, 
    97.23984, 96.8339, 97.72269, 97.11972, 98.24143, 97.63754, 98.27935, 
    98.16257, 98.35593, 98.52934, 98.74769, 99.15141, 99.05782, 99.39595, 
    95.97394, 96.17722, 96.15925, 96.37218, 96.52986, 96.87207, 97.42251, 
    97.21529, 97.59585, 97.67238, 97.09425, 97.44903, 96.31335, 96.49637, 
    96.38733, 95.99, 97.2631, 96.60852, 97.81924, 97.46309, 98.50462, 
    97.98589, 99.00634, 99.44463, 99.84852, 100.3182, 96.2882, 96.14996, 
    96.39751, 96.74075, 97.05971, 97.4848, 97.52832, 97.60812, 97.81493, 
    97.98904, 97.63342, 98.03271, 96.53896, 97.32001, 96.09779, 96.46494, 
    96.72047, 96.60826, 97.1916, 97.32941, 97.89065, 97.60025, 99.33641, 
    98.56608, 100.6764, 100.0926, 96.1017, 96.2877, 96.93678, 96.62761, 
    97.51318, 97.73193, 97.90991, 98.13781, 98.16239, 98.29758, 98.07611, 
    98.2888, 97.48571, 97.8441, 96.86238, 97.10082, 96.99107, 96.8708, 
    97.24226, 97.63903, 97.64742, 97.77487, 98.13472, 97.51678, 99.43627, 
    98.24842, 96.49076, 96.8502, 96.90149, 96.76213, 97.70999, 97.36593, 
    98.29427, 98.04284, 98.45497, 98.25005, 98.21993, 97.95714, 97.79376, 
    97.38171, 97.04716, 96.78233, 96.84386, 97.13492, 97.66331, 98.16466, 
    98.05472, 98.42361, 97.44881, 97.85693, 97.6991, 98.11091, 97.2098, 
    97.97714, 97.01427, 97.09845, 97.3591, 97.8847, 98.00107, 98.12558, 
    98.04872, 97.67673, 97.61581, 97.35274, 97.28023, 97.08012, 96.91467, 
    97.06585, 97.22478, 97.67684, 98.08534, 98.53183, 98.64124, 99.165, 
    98.73865, 99.44293, 98.84418, 99.87183, 98.02157, 98.8264, 97.37094, 
    97.52711, 97.81004, 98.4606, 98.10897, 98.52023, 97.61342, 97.14502, 
    97.02392, 96.79843, 97.02908, 97.01031, 97.2313, 97.16024, 97.69187, 
    97.40608, 98.2192, 98.51695, 99.36052, 99.86979, 100.3835, 100.6109, 
    100.6801, 100.7091,
  129.4504, 130.1381, 130.0042, 130.5603, 130.2516, 130.616, 129.5896, 
    130.1655, 129.7976, 129.5121, 131.6441, 130.5851, 132.7492, 132.0697, 
    133.7806, 132.6434, 134.0107, 133.7476, 134.54, 134.3127, 135.3298, 
    134.645, 135.8586, 135.166, 135.2742, 134.6225, 130.7977, 131.512, 
    130.7555, 130.8571, 130.8115, 130.258, 129.9798, 129.3978, 129.5033, 
    129.9307, 130.9029, 130.5723, 131.4062, 131.3874, 132.3198, 131.8989, 
    133.4723, 133.0238, 134.3222, 133.9949, 134.3068, 134.2122, 134.308, 
    133.8283, 134.0337, 133.612, 131.9777, 132.4567, 131.0313, 130.1792, 
    129.6148, 129.2154, 129.2718, 129.3794, 129.9332, 130.4552, 130.8539, 
    131.1211, 131.3846, 132.1848, 132.6093, 133.5631, 133.3906, 133.6829, 
    133.9624, 134.4326, 134.3551, 134.5626, 133.6751, 134.2646, 133.2924, 
    133.5578, 131.4568, 130.6614, 130.3246, 130.03, 129.3152, 129.8086, 
    129.6139, 130.0771, 130.3721, 130.2261, 131.1284, 130.7772, 132.6345, 
    131.8324, 133.9298, 133.426, 134.0507, 133.7317, 134.2787, 133.7863, 
    134.6398, 134.8262, 134.6988, 135.1883, 133.759, 134.3069, 130.2221, 
    130.2459, 130.3567, 129.8699, 129.8401, 129.395, 129.791, 129.9599, 
    130.3892, 130.6436, 130.8857, 131.419, 132.0164, 132.8545, 133.4586, 
    133.8645, 133.6155, 133.8354, 133.5896, 133.4745, 134.7564, 134.0357, 
    135.1178, 135.0578, 134.5676, 135.0646, 130.2626, 130.1257, 129.6512, 
    130.0224, 129.3465, 129.7246, 129.9424, 130.7846, 130.97, 131.1422, 
    131.4826, 131.9204, 132.6906, 133.363, 133.9787, 133.9335, 133.9494, 
    134.0872, 133.7461, 134.1432, 134.21, 134.0355, 135.0498, 134.7595, 
    135.0565, 134.8675, 130.1702, 130.4006, 130.276, 130.5103, 130.3453, 
    131.0804, 131.3013, 132.338, 131.9118, 132.5904, 131.9806, 132.0885, 
    132.6128, 132.0135, 133.326, 132.4354, 134.0925, 133.2002, 134.1486, 
    133.976, 134.2618, 134.5182, 134.841, 135.4382, 135.2998, 135.8, 
    130.7446, 131.0444, 131.0179, 131.3321, 131.5647, 132.0698, 132.8826, 
    132.5765, 133.1386, 133.2516, 132.3978, 132.9217, 131.2453, 131.5153, 
    131.3544, 130.7683, 132.6471, 131.6808, 133.4686, 132.9425, 134.4816, 
    133.7149, 135.2236, 135.8721, 136.4837, 137.2012, 131.2082, 131.0042, 
    131.3694, 131.876, 132.3468, 132.9746, 133.0388, 133.1567, 133.4622, 
    133.7195, 133.1941, 133.7841, 131.5782, 132.7312, 130.9273, 131.4689, 
    131.846, 131.6804, 132.5416, 132.7451, 133.5741, 133.1451, 135.7119, 
    134.5725, 137.7487, 136.8565, 130.933, 131.2074, 132.1653, 131.709, 
    133.0165, 133.3396, 133.6026, 133.9394, 133.9757, 134.1755, 133.8482, 
    134.1626, 132.9759, 133.5054, 132.0555, 132.4075, 132.2455, 132.0679, 
    132.6164, 133.2024, 133.2148, 133.4031, 133.9348, 133.0218, 135.8597, 
    134.1029, 131.507, 132.0375, 132.1132, 131.9075, 133.3072, 132.799, 
    134.1706, 133.799, 134.4082, 134.1053, 134.0608, 133.6724, 133.431, 
    132.8223, 132.3283, 131.9373, 132.0282, 132.4579, 133.2383, 133.9791, 
    133.8166, 134.3619, 132.9214, 133.5243, 133.2911, 133.8996, 132.5684, 
    133.7019, 132.2797, 132.404, 132.7889, 133.5654, 133.7373, 133.9213, 
    133.8077, 133.2581, 133.1681, 132.7795, 132.6724, 132.3769, 132.1327, 
    132.3559, 132.5906, 133.2582, 133.8618, 134.5219, 134.6836, 135.4583, 
    134.8277, 135.8696, 134.9837, 136.5193, 133.7676, 134.9575, 132.8064, 
    133.037, 133.455, 134.4165, 133.8968, 134.5047, 133.1646, 132.4728, 
    132.294, 131.9611, 132.3016, 132.2739, 132.6002, 132.4953, 133.2804, 
    132.8583, 134.0597, 134.4998, 135.7476, 136.5162, 137.3011, 137.6486, 
    137.7544, 137.7987,
  194.4182, 195.5316, 195.3148, 196.1981, 195.7148, 196.2854, 194.6435, 
    195.576, 194.9803, 194.5181, 197.8958, 196.237, 199.6292, 198.5633, 
    201.2486, 199.4631, 201.61, 201.1967, 202.442, 202.0846, 203.6839, 
    202.607, 204.5163, 203.4263, 203.5966, 202.5716, 196.5698, 197.6888, 
    196.5037, 196.663, 196.5915, 195.7249, 195.2751, 194.3331, 194.5039, 
    195.1958, 196.7346, 196.2169, 197.5232, 197.4937, 198.9555, 198.2954, 
    200.7643, 200.0603, 202.0995, 201.5853, 202.0754, 201.9267, 202.0773, 
    201.3235, 201.6462, 200.9838, 198.419, 199.1703, 196.9358, 195.5981, 
    194.6843, 194.0379, 194.1292, 194.3034, 195.1999, 196.0336, 196.6579, 
    197.0764, 197.4894, 198.7438, 199.4097, 200.907, 200.636, 201.0951, 
    201.5342, 202.2731, 202.1513, 202.4774, 201.0828, 202.009, 200.4818, 
    200.8987, 197.6024, 196.3564, 195.8291, 195.3565, 194.1994, 194.998, 
    194.6829, 195.4329, 195.9035, 195.6743, 197.0879, 196.5377, 199.4492, 
    198.1913, 201.4829, 200.6916, 201.6729, 201.1717, 202.0311, 201.2575, 
    202.5989, 202.8919, 202.6916, 203.4615, 201.2147, 202.0754, 195.6677, 
    195.7059, 195.8794, 195.0973, 195.0491, 194.3285, 194.9696, 195.243, 
    195.9302, 196.3285, 196.7077, 197.5433, 198.4797, 199.7944, 200.7428, 
    201.3804, 200.9892, 201.3346, 200.9486, 200.7678, 202.7821, 201.6493, 
    203.3506, 203.2562, 202.4852, 203.2668, 195.732, 195.5115, 194.7433, 
    195.3443, 194.2501, 194.8621, 195.2147, 196.5493, 196.8398, 197.1095, 
    197.643, 198.3292, 199.5373, 200.5927, 201.5597, 201.4887, 201.5137, 
    201.7302, 201.1943, 201.8183, 201.9232, 201.6491, 203.2435, 202.787, 
    203.2542, 202.9568, 195.5836, 195.9481, 195.7531, 196.1199, 195.8615, 
    197.0126, 197.3587, 198.9841, 198.3157, 199.38, 198.4236, 198.5928, 
    199.4151, 198.4751, 200.5345, 199.1368, 201.7386, 200.337, 201.8267, 
    201.5555, 202.0047, 202.4076, 202.9153, 203.8546, 203.6368, 204.4241, 
    196.4867, 196.9563, 196.9148, 197.407, 197.7716, 198.5635, 199.8385, 
    199.3583, 200.2404, 200.4179, 199.0779, 199.8999, 197.271, 197.6941, 
    197.442, 196.5238, 199.469, 197.9536, 200.7585, 199.9326, 202.3501, 
    201.1453, 203.517, 204.5374, 205.5007, 206.6313, 197.2129, 196.8934, 
    197.4656, 198.2595, 198.9979, 199.9829, 200.0838, 200.2688, 200.7486, 
    201.1526, 200.3275, 201.254, 197.7926, 199.6009, 196.7728, 197.6214, 
    198.2126, 197.953, 199.3034, 199.6227, 200.9242, 200.2506, 204.2853, 
    202.493, 207.4948, 206.088, 196.7819, 197.2117, 198.7132, 197.9977, 
    200.0487, 200.556, 200.969, 201.498, 201.5551, 201.8691, 201.3548, 
    201.8487, 199.985, 200.8163, 198.541, 199.0931, 198.839, 198.5605, 
    199.4208, 200.3405, 200.36, 200.6556, 201.4907, 200.0571, 204.5179, 
    201.7547, 197.6812, 198.5128, 198.6316, 198.309, 200.5051, 199.7074, 
    201.8614, 201.2775, 202.2348, 201.7587, 201.6887, 201.0786, 200.6994, 
    199.7439, 198.9689, 198.3558, 198.4982, 199.1721, 200.3968, 201.5603, 
    201.3051, 202.1619, 199.8995, 200.846, 200.4798, 201.4355, 199.3456, 
    201.1248, 198.8927, 199.0876, 199.6915, 200.9104, 201.1805, 201.4696, 
    201.2912, 200.4279, 200.2867, 199.6768, 199.5087, 199.0452, 198.6621, 
    199.0121, 199.3803, 200.4282, 201.3762, 202.4134, 202.6677, 203.8862, 
    202.8941, 204.5334, 203.1395, 205.5566, 201.228, 203.0982, 199.719, 
    200.081, 200.7372, 202.2478, 201.431, 202.3864, 200.2811, 199.1955, 
    198.9151, 198.393, 198.927, 198.8835, 199.3954, 199.2308, 200.4631, 
    199.8004, 201.687, 202.3788, 204.3415, 205.5518, 206.7889, 207.3368, 
    207.5038, 207.5737,
  318.5583, 320.3577, 320.0071, 321.464, 320.655, 321.6101, 318.9223, 
    320.4294, 319.4665, 318.7198, 324.3092, 321.5291, 327.1899, 325.4295, 
    329.8228, 326.9202, 330.4111, 329.7385, 331.7664, 331.1842, 333.7917, 
    332.0354, 335.1509, 333.3713, 333.6492, 331.9777, 322.0866, 323.9619, 
    321.9758, 322.2426, 322.1228, 320.6718, 319.943, 318.4211, 318.6968, 
    319.8148, 322.3625, 321.4954, 323.6845, 323.6349, 326.0882, 324.9799, 
    329.035, 327.8904, 331.2085, 330.371, 331.1691, 330.9269, 331.1723, 
    329.9448, 330.4702, 329.3921, 325.1873, 326.4448, 322.6997, 320.4651, 
    318.9883, 317.9443, 318.0917, 318.3729, 319.8214, 321.1886, 322.2342, 
    322.9355, 323.6278, 325.7325, 326.8334, 329.2671, 328.8264, 329.5731, 
    330.2878, 331.4913, 331.2928, 331.8242, 329.5533, 331.0609, 328.5757, 
    329.2536, 323.817, 321.7291, 320.8461, 320.0745, 318.2051, 319.4951, 
    318.986, 320.1982, 320.9707, 320.5884, 322.9547, 322.0328, 326.8976, 
    324.8051, 330.2043, 328.9168, 330.5136, 329.6978, 331.097, 329.8375, 
    332.0221, 332.4997, 332.1733, 333.4288, 329.7678, 331.1692, 320.5777, 
    320.64, 320.9305, 319.6555, 319.5777, 318.4135, 319.4491, 319.8911, 
    321.0155, 321.6824, 322.3176, 323.7181, 325.2892, 327.4584, 329.0001, 
    330.0375, 329.4009, 329.9629, 329.3348, 329.0408, 332.3207, 330.4752, 
    333.2479, 333.0939, 331.8369, 333.1112, 320.6838, 320.3252, 319.0835, 
    320.0549, 318.287, 319.2755, 319.8453, 322.0522, 322.5388, 322.9909, 
    323.8853, 325.0366, 327.0407, 328.756, 330.3294, 330.2138, 330.2545, 
    330.607, 329.7346, 330.7504, 330.9213, 330.4749, 333.0733, 332.3289, 
    333.0906, 332.6057, 320.4417, 321.0454, 320.7191, 321.3331, 320.9005, 
    322.8285, 323.4086, 326.1361, 325.0139, 326.7853, 325.195, 325.4792, 
    326.8421, 325.2816, 328.6613, 326.3904, 330.6207, 328.3401, 330.7641, 
    330.3225, 331.0539, 331.7104, 332.5379, 334.0704, 333.7149, 335.0003, 
    321.9474, 322.7341, 322.6646, 323.4896, 324.1011, 325.4299, 327.53, 
    326.7501, 328.1832, 328.4717, 326.2939, 327.6299, 323.2615, 323.971, 
    323.5483, 322.0094, 326.9298, 324.4062, 329.0257, 327.6829, 331.6167, 
    329.6548, 333.5193, 335.1853, 336.76, 338.6103, 323.1641, 322.6287, 
    323.5878, 324.9196, 326.1594, 327.7647, 327.9287, 328.2294, 329.0095, 
    329.6668, 328.3247, 329.8318, 324.136, 327.1441, 322.4266, 323.8491, 
    324.8409, 324.4053, 326.661, 327.1796, 329.2952, 328.1998, 334.7735, 
    331.8494, 340.0253, 337.7209, 322.4418, 323.1622, 325.6813, 324.4804, 
    327.8716, 328.6963, 329.368, 330.2289, 330.3218, 330.8331, 329.9958, 
    330.7999, 327.7681, 329.1195, 325.3922, 326.3194, 325.8925, 325.425, 
    326.8516, 328.3458, 328.3776, 328.8582, 330.2167, 327.8852, 335.1532, 
    330.6467, 323.9494, 325.3447, 325.5442, 325.0028, 328.6135, 327.317, 
    330.8206, 329.87, 331.4288, 330.6533, 330.5394, 329.5463, 328.9296, 
    327.3764, 326.1106, 325.0812, 325.3203, 326.4477, 328.4374, 330.3304, 
    329.9148, 331.3101, 327.6292, 329.1679, 328.5724, 330.1272, 326.7294, 
    329.6214, 325.9828, 326.3102, 327.2913, 329.2726, 329.7122, 330.1826, 
    329.8922, 328.488, 328.2584, 327.2674, 326.9944, 326.2389, 325.5955, 
    326.1833, 326.7857, 328.4885, 330.0305, 331.7198, 332.1344, 334.1218, 
    332.5034, 335.1785, 332.9033, 336.8512, 329.7894, 332.8362, 327.3359, 
    327.9241, 328.9909, 331.4499, 330.1199, 331.6758, 328.2494, 326.4856, 
    326.0203, 325.1438, 326.0403, 325.9673, 326.8103, 326.543, 328.5452, 
    327.4682, 330.5366, 331.6634, 334.8654, 336.8435, 338.8685, 339.7664, 
    340.0402, 340.1547,
  524.3475, 527.6201, 526.9819, 529.6358, 528.1615, 529.9022, 525.0089, 
    527.7507, 525.9983, 524.6409, 534.8331, 529.7545, 540.1705, 536.8851, 
    545.1851, 539.6578, 546.308, 545.0242, 548.8986, 547.7851, 552.779, 
    549.4134, 555.3896, 551.9727, 552.5056, 549.3029, 530.7715, 534.1978, 
    530.5694, 531.0561, 530.8376, 528.192, 526.8651, 524.0982, 524.5991, 
    526.6319, 531.2751, 529.6931, 533.6904, 533.5998, 538.0928, 536.0613, 
    543.6827, 541.5029, 547.8315, 546.2314, 547.7563, 547.2933, 547.7623, 
    545.4179, 546.4208, 544.3634, 536.4411, 538.7546, 531.8907, 527.8155, 
    525.1288, 523.2264, 523.5002, 524.0108, 526.6438, 529.1337, 531.0409, 
    532.3214, 533.5867, 537.4403, 539.493, 544.1251, 543.2852, 544.7087, 
    546.0725, 548.3723, 547.9929, 549.0091, 544.6708, 547.5494, 542.8076, 
    544.0994, 533.9326, 530.1193, 528.5096, 527.1046, 523.7061, 526.0502, 
    525.1246, 527.3296, 528.7367, 528.0402, 532.3564, 530.6733, 539.615, 
    535.741, 545.9132, 543.4574, 546.5038, 544.9466, 547.6183, 545.2131, 
    549.3878, 550.3023, 549.6772, 552.0829, 545.0801, 547.7564, 528.0207, 
    528.1342, 528.6634, 526.3422, 526.2005, 524.0845, 525.9667, 526.7708, 
    528.8183, 530.0342, 531.1931, 533.752, 536.6279, 540.681, 543.6161, 
    545.5948, 544.3804, 545.4523, 544.2542, 543.6937, 549.9595, 546.4303, 
    551.7361, 551.4408, 549.0333, 551.4741, 528.2139, 527.561, 525.3018, 
    527.0688, 523.8547, 525.651, 526.6874, 530.7087, 531.597, 532.4226, 
    534.0576, 536.165, 539.8868, 543.1509, 546.1519, 545.9313, 546.009, 
    546.6821, 545.0168, 546.9561, 547.2825, 546.4297, 551.4012, 549.9752, 
    551.4345, 550.5053, 527.7731, 528.8729, 528.2783, 529.3971, 528.6086, 
    532.1259, 533.186, 538.1805, 536.1235, 539.4016, 536.4553, 536.976, 
    539.5094, 536.6139, 542.9706, 538.6514, 546.7083, 542.3587, 546.9823, 
    546.1389, 547.5361, 548.7914, 550.3755, 553.3138, 552.6316, 555.1, 
    530.5175, 531.9536, 531.8267, 533.3342, 534.4524, 536.8857, 540.8173, 
    539.3346, 542.0602, 542.6095, 538.47, 541.0072, 532.9172, 534.2144, 
    533.4414, 530.6307, 539.6761, 535.0107, 543.6649, 541.1081, 548.6122, 
    544.8644, 552.2566, 555.4557, 558.4688, 561.9195, 532.7391, 531.761, 
    533.5137, 535.9507, 538.2234, 541.2636, 541.5757, 542.1482, 543.634, 
    544.8874, 542.3295, 545.2021, 534.5162, 540.0834, 531.392, 533.9913, 
    535.8065, 535.0091, 539.1654, 540.1509, 544.1786, 542.0917, 554.6642, 
    549.0573, 564.5649, 560.2596, 531.4199, 532.7357, 537.3465, 535.1465, 
    541.4672, 543.0373, 544.3176, 545.96, 546.1376, 547.114, 545.5151, 
    547.0506, 541.2701, 543.8439, 536.8167, 538.5168, 537.7338, 536.8767, 
    539.5275, 542.3698, 542.4303, 543.3458, 545.9366, 541.493, 555.3938, 
    546.7578, 534.175, 536.7296, 537.0952, 536.1031, 542.8796, 540.4122, 
    547.0901, 545.2751, 548.2527, 546.7706, 546.553, 544.6576, 543.4818, 
    540.525, 538.1339, 536.2468, 536.6849, 538.7603, 542.5441, 546.1538, 
    545.3606, 548.0258, 541.0059, 543.936, 542.8013, 545.766, 539.2953, 
    544.8006, 537.8994, 538.5001, 540.3633, 544.1357, 544.9741, 545.8718, 
    545.3176, 542.6406, 542.2034, 540.3178, 539.7988, 538.3692, 537.1893, 
    538.2673, 539.4023, 542.6415, 545.5815, 548.8093, 549.6027, 553.4124, 
    550.3092, 555.4424, 551.0753, 558.6385, 545.1212, 550.9467, 540.4481, 
    541.5671, 543.5986, 548.2931, 545.752, 548.725, 542.1862, 538.8322, 
    537.9682, 536.3614, 538.005, 537.871, 539.4492, 538.9414, 542.7495, 
    540.6998, 546.5477, 548.7014, 554.8409, 558.6242, 562.4019, 564.0806, 
    564.5928, 564.8071,
  947.2584, 954.1312, 952.7881, 958.3819, 955.2715, 958.9448, 948.6444, 
    954.4061, 950.7208, 947.8731, 969.2601, 958.6327, 980.2999, 973.493, 
    990.7612, 979.2353, 993.116, 990.4244, 998.5654, 996.2202, 1006.774, 
    999.6512, 1012.327, 1005.063, 1006.194, 999.418, 960.7828, 967.9522, 
    960.3553, 961.3853, 960.9227, 955.3358, 952.5424, 946.7361, 947.7855, 
    952.0521, 961.8489, 958.5031, 966.9091, 966.7227, 975.9911, 971.7919, 
    987.618, 983.0712, 996.3179, 992.9552, 996.1596, 995.1858, 996.1723, 
    991.2491, 993.3528, 989.0411, 972.576, 977.3621, 963.1533, 954.5426, 
    948.896, 944.9249, 945.4845, 946.5532, 952.0771, 957.3218, 961.3531, 
    964.0666, 966.6959, 974.6408, 978.8933, 988.5425, 986.7874, 989.7637, 
    992.6218, 997.4564, 996.6575, 998.7985, 989.6844, 995.7243, 985.7904, 
    988.489, 967.4069, 959.4036, 956.0052, 953.0461, 945.9153, 950.8298, 
    948.8872, 953.5197, 956.4842, 955.0159, 964.141, 960.5753, 979.1464, 
    971.1312, 992.2876, 987.1471, 993.5271, 990.2618, 995.8694, 990.8199, 
    999.5973, 1001.528, 1000.208, 1005.297, 990.5414, 996.1598, 954.9749, 
    955.2141, 956.3296, 951.4432, 951.1456, 946.7075, 950.6545, 952.3442, 
    956.6563, 959.2236, 961.6752, 967.0354, 972.9616, 981.3611, 987.4789, 
    991.6199, 989.0767, 991.3214, 988.8127, 987.6409, 1000.804, 993.3727, 
    1004.562, 1003.937, 998.8496, 1004.007, 955.3821, 954.0067, 949.2589, 
    952.9709, 946.2264, 949.9916, 952.1687, 960.6501, 962.5308, 964.2812, 
    967.6639, 972.0061, 979.7109, 986.5072, 992.7885, 992.3256, 992.4885, 
    993.9015, 990.4088, 994.4771, 995.1631, 993.3715, 1003.853, 1000.837, 
    1003.923, 1001.957, 954.4533, 956.7714, 955.5176, 957.8779, 956.2142, 
    963.6519, 965.8724, 976.1727, 971.9204, 978.7036, 972.6053, 973.6808, 
    978.9274, 972.9329, 986.1307, 977.1479, 993.9564, 984.8542, 994.5322, 
    992.7611, 995.6964, 998.3395, 1001.683, 1007.909, 1006.461, 1011.71, 
    960.2454, 963.2866, 963.0177, 966.1768, 968.4763, 973.4944, 981.6444, 
    978.5647, 984.232, 985.3773, 976.7723, 982.0394, 965.3205, 967.9865, 
    966.3972, 960.485, 979.2734, 969.6259, 987.5806, 982.2493, 997.9619, 
    990.0897, 1005.665, 1012.468, 1018.949, 1026.627, 964.953, 962.8785, 
    966.5457, 971.5637, 976.2614, 982.5731, 983.2228, 984.4153, 987.5162, 
    990.1378, 984.7934, 990.797, 968.6076, 980.119, 962.0967, 967.5276, 
    971.2664, 969.6226, 978.2137, 980.2593, 988.6545, 984.2977, 1010.781, 
    998.9001, 1032.433, 1022.927, 962.1556, 964.9456, 974.4469, 969.9058, 
    982.9968, 986.2699, 988.9453, 992.3859, 992.7583, 994.8088, 991.4529, 
    994.6757, 982.5865, 987.9547, 973.3518, 976.8693, 975.248, 973.4758, 
    978.9649, 984.8773, 985.0035, 986.9141, 992.3367, 983.0505, 1012.336, 
    994.0604, 967.9055, 973.1718, 973.9273, 971.8783, 985.9409, 980.8021, 
    994.7587, 990.95, 997.2047, 994.0874, 993.6304, 989.6567, 987.1981, 
    981.0368, 976.076, 972.1749, 973.0794, 977.3737, 985.2409, 992.7924, 
    991.129, 996.7267, 982.0366, 988.1472, 985.7773, 991.9789, 978.4833, 
    989.9561, 975.5906, 976.8345, 980.7006, 988.5648, 990.3193, 992.2007, 
    991.0389, 985.442, 984.5303, 980.6061, 979.5281, 976.5634, 974.1217, 
    976.3523, 978.7052, 985.444, 991.592, 998.3773, 1000.051, 1008.119, 
    1001.543, 1012.44, 1003.163, 1019.325, 990.6274, 1002.891, 980.877, 
    983.2047, 987.4421, 997.2896, 991.9496, 998.1996, 984.4946, 977.5229, 
    975.733, 972.4114, 975.8092, 975.532, 978.8023, 977.7491, 985.6693, 
    981.4001, 993.6191, 998.1498, 1011.158, 1019.293, 1027.704, 1031.382, 
    1032.494, 1032.959,
  1829.891, 1849.353, 1845.525, 1861.55, 1852.613, 1863.175, 1833.791, 
    1850.138, 1839.657, 1831.62, 1893.772, 1862.273, 1928.095, 1906.814, 
    1960.691, 1924.741, 1968.121, 1959.632, 1985.507, 1977.992, 2012.212, 
    1989.003, 2030.648, 2006.596, 2010.304, 1988.252, 1868.494, 1889.771, 
    1867.255, 1870.243, 1868.9, 1852.797, 1844.827, 1828.425, 1831.373, 
    1843.433, 1871.591, 1861.899, 1886.589, 1886.022, 1914.579, 1901.556, 
    1950.848, 1936.759, 1978.304, 1967.612, 1977.798, 1974.693, 1977.839, 
    1962.226, 1968.871, 1955.293, 1903.977, 1918.863, 1875.39, 1850.529, 
    1834.5, 1823.354, 1824.919, 1827.912, 1843.504, 1858.497, 1870.15, 
    1878.058, 1885.94, 1910.376, 1923.666, 1953.734, 1948.261, 1957.557, 
    1966.558, 1981.947, 1979.389, 1986.256, 1957.309, 1976.409, 1945.164, 
    1953.567, 1888.107, 1864.5, 1854.715, 1846.26, 1826.124, 1839.966, 
    1834.475, 1847.609, 1856.09, 1851.882, 1878.275, 1867.892, 1924.461, 
    1899.519, 1965.502, 1949.38, 1969.423, 1959.121, 1976.872, 1960.875, 
    1988.829, 1995.074, 1990.801, 2007.361, 1960, 1977.799, 1851.764, 
    1852.449, 1855.646, 1841.704, 1840.86, 1828.345, 1839.469, 1844.263, 
    1856.584, 1863.98, 1871.086, 1886.974, 1905.169, 1931.447, 1950.414, 
    1963.395, 1955.405, 1962.454, 1954.579, 1950.919, 1992.728, 1968.934, 
    2004.954, 2002.91, 1986.421, 2003.14, 1852.93, 1848.998, 1835.524, 
    1846.046, 1826.996, 1837.594, 1843.764, 1868.109, 1873.575, 1878.686, 
    1888.891, 1902.216, 1926.238, 1947.389, 1967.085, 1965.622, 1966.136, 
    1970.611, 1959.583, 1972.438, 1974.621, 1968.93, 2002.637, 1992.835, 
    2002.867, 1996.466, 1850.273, 1856.914, 1853.318, 1860.097, 1855.315, 
    1876.846, 1883.436, 1915.146, 1901.952, 1923.069, 1904.067, 1907.396, 
    1923.773, 1905.08, 1946.22, 1918.193, 1970.785, 1942.263, 1972.614, 
    1966.998, 1976.32, 1984.781, 1995.575, 2015.958, 2011.183, 2028.584, 
    1866.936, 1875.779, 1874.995, 1884.361, 1891.372, 1906.819, 1932.344, 
    1922.633, 1940.339, 1943.882, 1917.018, 1933.586, 1881.761, 1889.876, 
    1885.031, 1867.631, 1924.861, 1894.893, 1950.731, 1934.231, 1983.568, 
    1958.581, 2008.569, 2031.119, 2053.034, 2079.24, 1880.652, 1874.589, 
    1885.483, 1900.852, 1915.423, 1935.226, 1937.226, 1940.906, 1950.53, 
    1958.732, 1942.075, 1960.803, 1891.774, 1927.524, 1872.311, 1888.475, 
    1899.936, 1894.883, 1921.532, 1927.967, 1954.084, 1940.542, 2025.485, 
    1986.584, 2099.509, 2066.705, 1872.483, 1880.631, 1909.773, 1895.752, 
    1936.53, 1946.652, 1954.993, 1965.812, 1966.989, 1973.493, 1962.868, 
    1973.07, 1935.267, 1951.898, 1906.377, 1917.321, 1912.264, 1906.761, 
    1923.891, 1942.334, 1942.725, 1948.655, 1965.657, 1936.695, 2030.677, 
    1971.115, 1889.628, 1905.819, 1908.161, 1901.822, 1945.63, 1929.68, 
    1973.334, 1961.285, 1981.141, 1971.201, 1969.751, 1957.222, 1949.539, 
    1930.422, 1914.845, 1902.738, 1905.534, 1918.899, 1943.46, 1967.097, 
    1961.848, 1979.611, 1933.577, 1952.499, 1945.123, 1964.527, 1922.378, 
    1958.161, 1913.331, 1917.213, 1929.359, 1953.803, 1959.302, 1965.227, 
    1961.564, 1944.083, 1941.261, 1929.061, 1925.662, 1916.366, 1908.764, 
    1915.707, 1923.074, 1944.089, 1963.307, 1984.902, 1990.293, 2016.649, 
    1995.121, 2031.025, 2000.386, 2054.321, 1960.27, 1999.5, 1929.916, 
    1937.17, 1950.299, 1981.412, 1964.434, 1984.332, 1941.151, 1919.366, 
    1913.775, 1903.468, 1914.012, 1913.149, 1923.38, 1920.075, 1944.788, 
    1931.57, 1969.715, 1984.171, 2026.74, 2054.213, 2082.9, 2095.761, 
    2099.724, 2101.388,
  5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 5434.597, 
    5434.597, 5434.597,
  8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 8960.136, 
    8960.136, 8960.136,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILLIQ =
  4.483961, 4.502318, 4.498744, 4.513585, 4.505348, 4.515072, 4.487678, 
    4.503048, 4.493231, 4.48561, 4.542492, 4.514247, 4.571972, 4.553854, 
    4.599471, 4.56915, 4.605603, 4.598594, 4.619713, 4.613656, 4.640749, 
    4.622511, 4.654838, 4.636388, 4.639271, 4.621911, 4.51992, 4.538969, 
    4.518794, 4.521506, 4.520288, 4.505518, 4.498089, 4.48256, 4.485376, 
    4.496783, 4.522726, 4.513906, 4.536158, 4.535655, 4.560525, 4.549299, 
    4.591255, 4.5793, 4.613908, 4.605186, 4.613498, 4.610977, 4.613531, 
    4.600745, 4.60622, 4.59498, 4.5514, 4.564175, 4.526154, 4.50341, 
    4.488351, 4.477689, 4.479195, 4.482068, 4.49685, 4.510782, 4.521422, 
    4.528551, 4.535582, 4.55692, 4.568243, 4.593675, 4.589077, 4.596868, 
    4.60432, 4.616851, 4.614787, 4.620314, 4.596662, 4.612371, 4.58646, 
    4.593536, 4.537497, 4.516284, 4.507292, 4.499432, 4.480353, 4.493522, 
    4.488327, 4.500693, 4.508564, 4.50467, 4.528746, 4.519373, 4.568915, 
    4.547525, 4.60345, 4.59002, 4.606673, 4.59817, 4.612747, 4.599626, 
    4.622372, 4.627336, 4.623943, 4.636985, 4.5989, 4.613499, 4.50456, 
    4.505196, 4.508154, 4.495159, 4.494365, 4.482482, 4.493054, 4.497562, 
    4.50902, 4.515809, 4.522269, 4.536499, 4.552432, 4.574782, 4.59089, 
    4.601711, 4.595074, 4.600934, 4.594383, 4.591315, 4.625476, 4.606271, 
    4.635108, 4.633509, 4.620445, 4.633689, 4.505641, 4.501988, 4.489323, 
    4.499232, 4.48119, 4.491282, 4.497094, 4.51957, 4.524519, 4.529113, 
    4.538196, 4.549873, 4.570413, 4.588341, 4.604753, 4.603549, 4.603973, 
    4.607645, 4.598553, 4.609139, 4.610918, 4.606268, 4.633295, 4.625561, 
    4.633475, 4.628438, 4.503175, 4.509325, 4.506001, 4.512253, 4.507848, 
    4.527461, 4.533354, 4.561008, 4.549643, 4.56774, 4.551478, 4.554357, 
    4.568332, 4.552356, 4.587351, 4.563604, 4.607788, 4.583995, 4.609282, 
    4.604682, 4.612299, 4.61913, 4.627734, 4.643641, 4.639953, 4.653278, 
    4.518505, 4.526503, 4.525798, 4.534179, 4.540385, 4.553859, 4.575532, 
    4.567372, 4.58236, 4.585373, 4.562607, 4.576575, 4.531862, 4.539064, 
    4.534775, 4.519135, 4.569252, 4.543479, 4.591156, 4.57713, 4.618156, 
    4.597719, 4.637925, 4.655192, 4.671485, 4.690579, 4.530873, 4.525433, 
    4.535177, 4.548685, 4.561245, 4.577985, 4.5797, 4.582842, 4.590988, 
    4.597846, 4.583837, 4.599566, 4.540736, 4.571494, 4.523377, 4.537826, 
    4.547888, 4.543472, 4.566441, 4.571867, 4.593968, 4.582533, 4.650927, 
    4.620574, 4.705154, 4.681406, 4.523533, 4.530854, 4.556404, 4.544233, 
    4.579104, 4.587718, 4.59473, 4.603705, 4.604675, 4.609999, 4.601276, 
    4.609654, 4.578021, 4.592137, 4.553477, 4.562864, 4.558544, 4.553809, 
    4.568435, 4.584057, 4.584391, 4.589408, 4.603572, 4.579246, 4.654856, 
    4.608053, 4.538847, 4.552994, 4.555016, 4.549531, 4.586854, 4.573304, 
    4.609869, 4.599966, 4.616201, 4.608128, 4.606941, 4.59659, 4.590154, 
    4.573925, 4.560751, 4.550326, 4.552748, 4.564207, 4.585013, 4.604763, 
    4.600431, 4.614966, 4.576569, 4.59264, 4.586424, 4.602646, 4.567156, 
    4.597367, 4.559458, 4.562772, 4.573035, 4.593732, 4.59832, 4.603223, 
    4.600197, 4.585543, 4.583145, 4.572785, 4.569929, 4.56205, 4.555536, 
    4.561488, 4.567745, 4.585548, 4.601638, 4.619227, 4.623539, 4.64417, 
    4.627372, 4.655118, 4.631522, 4.672422, 4.599121, 4.630828, 4.573503, 
    4.579652, 4.590793, 4.616418, 4.60257, 4.618768, 4.583051, 4.564602, 
    4.559838, 4.550959, 4.560041, 4.559302, 4.568004, 4.565206, 4.586141, 
    4.574886, 4.606912, 4.61864, 4.651881, 4.672346, 4.693244, 4.702491, 
    4.705308, 4.706486,
  5.614914, 5.637934, 5.633453, 5.65206, 5.641732, 5.653924, 5.619575, 
    5.63885, 5.626539, 5.616982, 5.6883, 5.652891, 5.725242, 5.702536, 
    5.759693, 5.721705, 5.767375, 5.758593, 5.785047, 5.777459, 5.811394, 
    5.788551, 5.829036, 5.805932, 5.809543, 5.787799, 5.660002, 5.683884, 
    5.65859, 5.66199, 5.660464, 5.641946, 5.632632, 5.613156, 5.616688, 
    5.630993, 5.66352, 5.652462, 5.680356, 5.679725, 5.710896, 5.696826, 
    5.749398, 5.734421, 5.777776, 5.766851, 5.777263, 5.774104, 5.777304, 
    5.761287, 5.768146, 5.754066, 5.69946, 5.71547, 5.667816, 5.639305, 
    5.62042, 5.607048, 5.608937, 5.61254, 5.631077, 5.648545, 5.661884, 
    5.67082, 5.679635, 5.70638, 5.720568, 5.752431, 5.74667, 5.756431, 
    5.765765, 5.781462, 5.778876, 5.7858, 5.756172, 5.775851, 5.74339, 
    5.752256, 5.68204, 5.655443, 5.644172, 5.634315, 5.61039, 5.626904, 
    5.62039, 5.635895, 5.645764, 5.640881, 5.671065, 5.659317, 5.72141, 
    5.694604, 5.764676, 5.747852, 5.768713, 5.758061, 5.776321, 5.759885, 
    5.788377, 5.794595, 5.790346, 5.806679, 5.758976, 5.777263, 5.640745, 
    5.641541, 5.645251, 5.628957, 5.627961, 5.61306, 5.626317, 5.63197, 
    5.646336, 5.654848, 5.662947, 5.680784, 5.700754, 5.728761, 5.748941, 
    5.762497, 5.754182, 5.761523, 5.753317, 5.749474, 5.792265, 5.76821, 
    5.804328, 5.802325, 5.785964, 5.80255, 5.6421, 5.637519, 5.621638, 
    5.634064, 5.611439, 5.624096, 5.631383, 5.659564, 5.665767, 5.671525, 
    5.68291, 5.697546, 5.723286, 5.745749, 5.766308, 5.7648, 5.76533, 
    5.769931, 5.758542, 5.771802, 5.77403, 5.768207, 5.802057, 5.792371, 
    5.802282, 5.795975, 5.639008, 5.646719, 5.642551, 5.65039, 5.644867, 
    5.669456, 5.676844, 5.711502, 5.697258, 5.719937, 5.699558, 5.703166, 
    5.720681, 5.700657, 5.74451, 5.714756, 5.77011, 5.740306, 5.771981, 
    5.766219, 5.775761, 5.784317, 5.795092, 5.815014, 5.810396, 5.827083, 
    5.658227, 5.668255, 5.66737, 5.677876, 5.685655, 5.702541, 5.7297, 
    5.719475, 5.738254, 5.74203, 5.713503, 5.731008, 5.674972, 5.684, 
    5.678623, 5.659018, 5.721832, 5.689534, 5.749276, 5.731702, 5.783097, 
    5.757498, 5.807856, 5.829482, 5.849879, 5.873788, 5.673732, 5.666912, 
    5.679126, 5.696059, 5.711798, 5.732773, 5.734922, 5.738859, 5.749064, 
    5.757656, 5.740106, 5.75981, 5.686098, 5.724641, 5.664336, 5.682449, 
    5.695059, 5.689523, 5.718307, 5.725107, 5.752799, 5.738471, 5.82414, 
    5.786127, 5.892033, 5.862302, 5.664531, 5.673707, 5.705731, 5.690478, 
    5.734175, 5.744968, 5.753751, 5.764996, 5.76621, 5.77288, 5.761952, 
    5.772448, 5.732818, 5.750504, 5.702063, 5.713827, 5.708412, 5.702478, 
    5.720807, 5.740382, 5.740798, 5.747086, 5.764835, 5.734352, 5.829063, 
    5.770447, 5.683727, 5.701458, 5.703992, 5.697116, 5.743886, 5.726908, 
    5.772717, 5.76031, 5.780648, 5.770535, 5.769049, 5.756082, 5.748019, 
    5.727686, 5.711179, 5.698113, 5.701149, 5.715509, 5.74158, 5.766321, 
    5.760895, 5.7791, 5.730999, 5.751135, 5.743347, 5.763669, 5.719204, 
    5.75706, 5.709558, 5.713711, 5.726571, 5.752504, 5.758249, 5.764392, 
    5.760601, 5.742243, 5.739238, 5.726258, 5.722679, 5.712806, 5.704643, 
    5.712101, 5.719943, 5.742249, 5.762406, 5.784439, 5.789839, 5.815681, 
    5.794641, 5.829391, 5.799843, 5.851058, 5.759256, 5.798971, 5.727156, 
    5.734862, 5.748821, 5.780922, 5.763573, 5.783865, 5.73912, 5.716006, 
    5.710033, 5.698907, 5.710288, 5.709362, 5.720266, 5.71676, 5.742991, 
    5.72889, 5.769012, 5.783704, 5.825334, 5.850959, 5.87712, 5.888698, 
    5.892224, 5.893699,
  8.093365, 8.12752, 8.12087, 8.148486, 8.133156, 8.151254, 8.100279, 
    8.12888, 8.110611, 8.096433, 8.2023, 8.149719, 8.257191, 8.223448, 
    8.308416, 8.251934, 8.319841, 8.306779, 8.346133, 8.334844, 8.385349, 
    8.351348, 8.411619, 8.377217, 8.382593, 8.350229, 8.160275, 8.195741, 
    8.158179, 8.163228, 8.160961, 8.133473, 8.119653, 8.090757, 8.095996, 
    8.117221, 8.165499, 8.149082, 8.190499, 8.189562, 8.235868, 8.214964, 
    8.293105, 8.270835, 8.335315, 8.319062, 8.334552, 8.329852, 8.334613, 
    8.310786, 8.320989, 8.300045, 8.218877, 8.242667, 8.171878, 8.129555, 
    8.101532, 8.081697, 8.084498, 8.089843, 8.117345, 8.143269, 8.163071, 
    8.176338, 8.189427, 8.22916, 8.250244, 8.297616, 8.289047, 8.303564, 
    8.317447, 8.340799, 8.336951, 8.347254, 8.303179, 8.332452, 8.284171, 
    8.297355, 8.193002, 8.153507, 8.136778, 8.122149, 8.086654, 8.111153, 
    8.101488, 8.124494, 8.139141, 8.131893, 8.176702, 8.159258, 8.251495, 
    8.211663, 8.315826, 8.290805, 8.321832, 8.305987, 8.333152, 8.308702, 
    8.351089, 8.360344, 8.354019, 8.37833, 8.307347, 8.334553, 8.131691, 
    8.132873, 8.138378, 8.1142, 8.112721, 8.090614, 8.110282, 8.11867, 
    8.13999, 8.152623, 8.164648, 8.191134, 8.220799, 8.262422, 8.292425, 
    8.312587, 8.300219, 8.311137, 8.298933, 8.293217, 8.356876, 8.321084, 
    8.37483, 8.371848, 8.347499, 8.372184, 8.133702, 8.126904, 8.103339, 
    8.121776, 8.088209, 8.106986, 8.117799, 8.159625, 8.168835, 8.177385, 
    8.194293, 8.216033, 8.254284, 8.287678, 8.318254, 8.31601, 8.3168, 
    8.323644, 8.306703, 8.326427, 8.329742, 8.321078, 8.371449, 8.357034, 
    8.371785, 8.362396, 8.129113, 8.140556, 8.134372, 8.146007, 8.137809, 
    8.174314, 8.185284, 8.236771, 8.215606, 8.249307, 8.219023, 8.224383, 
    8.250413, 8.220656, 8.285836, 8.241606, 8.32391, 8.279586, 8.326694, 
    8.318122, 8.332316, 8.345048, 8.361083, 8.390738, 8.383863, 8.40871, 
    8.15764, 8.172529, 8.171215, 8.186816, 8.19837, 8.223454, 8.263817, 
    8.24862, 8.276534, 8.282147, 8.239744, 8.265761, 8.182504, 8.195912, 
    8.187925, 8.158815, 8.252123, 8.204132, 8.292923, 8.266794, 8.343232, 
    8.305151, 8.380081, 8.412282, 8.442664, 8.478292, 8.180662, 8.170535, 
    8.188672, 8.213824, 8.23721, 8.268386, 8.27158, 8.277433, 8.292608, 
    8.305385, 8.279287, 8.30859, 8.199029, 8.256298, 8.166711, 8.193608, 
    8.212339, 8.204116, 8.246883, 8.25699, 8.298162, 8.276856, 8.404328, 
    8.347742, 8.505489, 8.461175, 8.167, 8.180626, 8.228196, 8.205534, 
    8.27047, 8.286517, 8.299579, 8.316302, 8.318108, 8.328032, 8.311775, 
    8.327388, 8.268453, 8.294748, 8.222744, 8.240225, 8.232179, 8.223362, 
    8.250598, 8.279698, 8.280317, 8.289666, 8.316065, 8.270733, 8.41166, 
    8.324412, 8.195505, 8.221847, 8.225611, 8.215395, 8.284907, 8.259667, 
    8.327788, 8.309333, 8.339588, 8.324543, 8.322331, 8.303043, 8.291055, 
    8.260824, 8.236291, 8.216876, 8.221387, 8.242724, 8.28148, 8.318274, 
    8.310204, 8.337285, 8.265747, 8.295688, 8.284106, 8.314329, 8.248217, 
    8.304501, 8.233881, 8.240052, 8.259167, 8.297724, 8.306268, 8.315405, 
    8.309765, 8.282465, 8.277997, 8.2587, 8.253381, 8.238708, 8.226578, 
    8.237661, 8.249314, 8.282475, 8.312451, 8.34523, 8.353265, 8.391731, 
    8.360414, 8.412149, 8.368156, 8.444421, 8.307766, 8.366858, 8.260036, 
    8.271491, 8.292246, 8.339996, 8.314187, 8.344376, 8.277822, 8.243464, 
    8.234588, 8.218056, 8.234966, 8.233589, 8.249795, 8.244584, 8.283578, 
    8.262613, 8.322277, 8.344136, 8.406104, 8.444273, 8.483258, 8.500517, 
    8.505774, 8.507974,
  12.6655, 12.72097, 12.71016, 12.75503, 12.73012, 12.75953, 12.67672, 
    12.72317, 12.6935, 12.67048, 12.84254, 12.75704, 12.9319, 12.87696, 
    13.01538, 12.92334, 13.03401, 13.01271, 13.07691, 13.05849, 13.14093, 
    13.08542, 13.18384, 13.12765, 13.13643, 13.08359, 12.7742, 12.83187, 
    12.77079, 12.779, 12.77531, 12.73064, 12.70819, 12.66126, 12.66977, 
    12.70424, 12.78269, 12.756, 12.82334, 12.82182, 12.89718, 12.86315, 
    12.99042, 12.95413, 13.05925, 13.03274, 13.05801, 13.05034, 13.05811, 
    13.01925, 13.03588, 13.00173, 12.86952, 12.90825, 12.79306, 12.72427, 
    12.67876, 12.64656, 12.6511, 12.65978, 12.70444, 12.74655, 12.77874, 
    12.80031, 12.8216, 12.88626, 12.92059, 12.99777, 12.98381, 13.00747, 
    13.03011, 13.0682, 13.06192, 13.07874, 13.00684, 13.05458, 12.97586, 
    12.99735, 12.82741, 12.7632, 12.73601, 12.71224, 12.6546, 12.69438, 
    12.67869, 12.71605, 12.73985, 12.72807, 12.8009, 12.77254, 12.92262, 
    12.85778, 13.02747, 12.98667, 13.03726, 13.01142, 13.05573, 13.01585, 
    13.08499, 13.1001, 13.08978, 13.12947, 13.01364, 13.05801, 12.72774, 
    12.72966, 12.73861, 12.69933, 12.69693, 12.66103, 12.69297, 12.70659, 
    12.74123, 12.76176, 12.7813, 12.82438, 12.87265, 12.94042, 12.98931, 
    13.02218, 13.00202, 13.01982, 12.99992, 12.9906, 13.09444, 13.03604, 
    13.12375, 13.11888, 13.07914, 13.11943, 12.73101, 12.71996, 12.68169, 
    12.71163, 12.65713, 12.68761, 12.70518, 12.77314, 12.78811, 12.80202, 
    12.82951, 12.86489, 12.92716, 12.98157, 13.03142, 13.02777, 13.02905, 
    13.04022, 13.01259, 13.04476, 13.05016, 13.03603, 13.11823, 13.0947, 
    13.11878, 13.10345, 12.72355, 12.74215, 12.7321, 12.751, 12.73768, 
    12.79702, 12.81486, 12.89864, 12.86419, 12.91906, 12.86975, 12.87848, 
    12.92086, 12.87241, 12.97857, 12.90652, 13.04065, 12.96838, 13.04519, 
    13.03121, 13.05436, 13.07514, 13.10131, 13.14973, 13.1385, 13.17909, 
    12.76991, 12.79412, 12.79198, 12.81735, 12.83615, 12.87697, 12.94269, 
    12.91794, 12.96341, 12.97256, 12.90349, 12.94586, 12.81034, 12.83215, 
    12.81916, 12.77182, 12.92365, 12.84552, 12.99012, 12.94754, 13.07217, 
    13.01006, 13.13233, 13.18493, 13.23459, 13.29288, 12.80734, 12.79088, 
    12.82037, 12.86129, 12.89936, 12.95014, 12.95534, 12.96488, 12.98961, 
    13.01044, 12.9679, 13.01567, 12.83722, 12.93045, 12.78466, 12.8284, 
    12.85888, 12.8455, 12.91511, 12.93157, 12.99866, 12.96394, 13.17193, 
    13.07953, 13.3374, 13.26487, 12.78513, 12.80729, 12.88469, 12.8478, 
    12.95353, 12.97968, 13.00097, 13.02824, 13.03119, 13.04737, 13.02086, 
    13.04632, 12.95025, 12.9931, 12.87581, 12.90427, 12.89117, 12.87682, 
    12.92116, 12.96857, 12.96958, 12.98481, 13.02785, 12.95396, 13.18391, 
    13.04147, 12.83149, 12.87435, 12.88048, 12.86385, 12.97706, 12.93593, 
    13.04698, 13.01688, 13.06623, 13.04168, 13.03808, 13.00662, 12.98708, 
    12.93782, 12.89786, 12.86626, 12.8736, 12.90834, 12.97147, 13.03146, 
    13.0183, 13.06247, 12.94584, 12.99463, 12.97575, 13.02502, 12.91728, 
    13.009, 12.89394, 12.90399, 12.93512, 12.99795, 13.01188, 13.02678, 
    13.01758, 12.97308, 12.9658, 12.93436, 12.92569, 12.9018, 12.88205, 
    12.90009, 12.91907, 12.97309, 13.02196, 13.07543, 13.08855, 13.15135, 
    13.10021, 13.18471, 13.11285, 13.23747, 13.01432, 13.11073, 12.93653, 
    12.9552, 12.98902, 13.06689, 13.02479, 13.07404, 12.96551, 12.90954, 
    12.89509, 12.86818, 12.89571, 12.89347, 12.91985, 12.91137, 12.97489, 
    12.94073, 13.03799, 13.07365, 13.17483, 13.23723, 13.30101, 13.32926, 
    13.33787, 13.34147,
  20.5999, 20.69597, 20.67725, 20.75503, 20.71184, 20.76283, 20.61933, 
    20.6998, 20.64838, 20.60852, 20.90694, 20.75851, 21.06235, 20.96676, 
    21.20782, 21.04745, 21.24033, 21.20317, 21.31521, 21.28304, 21.42711, 
    21.33008, 21.50221, 21.40389, 21.41924, 21.32689, 20.78827, 20.8884, 
    20.78236, 20.7966, 20.79021, 20.71273, 20.67382, 20.59257, 20.60729, 
    20.66698, 20.80301, 20.75671, 20.87359, 20.87094, 21.00193, 20.94275, 
    21.1643, 21.10106, 21.28439, 21.23811, 21.28221, 21.26883, 21.28238, 
    21.21457, 21.2436, 21.18402, 20.95382, 21.02118, 20.82101, 20.7017, 
    20.62285, 20.56712, 20.57499, 20.59, 20.66733, 20.74033, 20.79615, 
    20.8336, 20.87056, 20.98293, 21.04266, 21.17712, 21.15277, 21.19403, 
    21.23351, 21.30001, 21.28905, 21.31841, 21.19293, 21.27623, 21.13892, 
    21.17638, 20.88066, 20.76919, 20.72204, 20.68085, 20.58104, 20.64991, 
    20.62273, 20.68745, 20.7287, 20.70828, 20.83462, 20.7854, 21.04621, 
    20.93341, 21.2289, 21.15777, 21.246, 21.20092, 21.27822, 21.20864, 
    21.32934, 21.35573, 21.33769, 21.40706, 21.20479, 21.28222, 20.70771, 
    20.71104, 20.72655, 20.65848, 20.65432, 20.59217, 20.64746, 20.67106, 
    20.73109, 20.7667, 20.8006, 20.87538, 20.95926, 21.07719, 21.16237, 
    21.21969, 21.18452, 21.21556, 21.18086, 21.16462, 21.34584, 21.24387, 
    21.39707, 21.38856, 21.31911, 21.38952, 20.71338, 20.69423, 20.62794, 
    20.6798, 20.58541, 20.63819, 20.66861, 20.78644, 20.81242, 20.83655, 
    20.88431, 20.94578, 21.05411, 21.14888, 21.23581, 21.22943, 21.23168, 
    21.25115, 21.20295, 21.25908, 21.26852, 21.24385, 21.38742, 21.34629, 
    21.38838, 21.36159, 20.70045, 20.73269, 20.71526, 20.74804, 20.72495, 
    20.82788, 20.85885, 21.00448, 20.94457, 21.04, 20.95424, 20.9694, 
    21.04314, 20.95886, 21.14365, 21.01818, 21.25191, 21.1259, 21.25983, 
    21.23544, 21.27585, 21.31212, 21.35784, 21.44251, 21.42287, 21.49389, 
    20.78084, 20.82284, 20.81914, 20.86318, 20.89583, 20.96678, 21.08115, 
    21.03805, 21.11724, 21.13317, 21.0129, 21.08666, 20.851, 20.88888, 
    20.86632, 20.78415, 21.04798, 20.91212, 21.16378, 21.08959, 21.30694, 
    21.19854, 21.41207, 21.50411, 21.59112, 21.69336, 20.8458, 20.81721, 
    20.86843, 20.93953, 21.00573, 21.09411, 21.10317, 21.11979, 21.16289, 
    21.19921, 21.12505, 21.20832, 20.89769, 21.05982, 20.80643, 20.88237, 
    20.93533, 20.91207, 21.03313, 21.06178, 21.17867, 21.11815, 21.48136, 
    21.3198, 21.77154, 21.64421, 20.80724, 20.8457, 20.9802, 20.91608, 
    21.10002, 21.14558, 21.1827, 21.23026, 21.2354, 21.26364, 21.21738, 
    21.26181, 21.0943, 21.16897, 20.96477, 21.01427, 20.99148, 20.96651, 
    21.04366, 21.12622, 21.12798, 21.15453, 21.22958, 21.10077, 21.50233, 
    21.25334, 20.88773, 20.96223, 20.97288, 20.94397, 21.14101, 21.06938, 
    21.26295, 21.21043, 21.29656, 21.25371, 21.24742, 21.19255, 21.15847, 
    21.07266, 21.00312, 20.94816, 20.96092, 21.02135, 21.13128, 21.23587, 
    21.21291, 21.29, 21.08662, 21.17164, 21.13874, 21.22465, 21.03691, 
    21.19669, 20.9963, 21.01378, 21.06796, 21.17743, 21.20172, 21.22771, 
    21.21166, 21.13408, 21.12139, 21.06664, 21.05155, 21.00997, 20.97562, 
    21.007, 21.04002, 21.1341, 21.2193, 21.31264, 21.33554, 21.44535, 
    21.35593, 21.50373, 21.37802, 21.59616, 21.20598, 21.37431, 21.07042, 
    21.10292, 21.16186, 21.29772, 21.22424, 21.3102, 21.12089, 21.02344, 
    20.9983, 20.9515, 20.99937, 20.99547, 21.04138, 21.02662, 21.13724, 
    21.07773, 21.24726, 21.30952, 21.48644, 21.59573, 21.70762, 21.75724, 
    21.77237, 21.77869,
  34.64178, 34.82255, 34.7873, 34.9339, 34.85246, 34.94861, 34.67831, 
    34.82977, 34.73297, 34.65799, 35.22099, 34.94045, 35.51581, 35.33433, 
    35.79281, 35.48749, 35.85484, 35.78393, 35.99794, 35.93643, 36.21229, 
    36.02638, 36.3565, 36.16775, 36.19719, 36.02027, 34.99663, 35.18589, 
    34.98547, 35.01235, 35.00028, 34.85415, 34.78085, 34.62801, 34.65568, 
    34.76797, 35.02445, 34.93707, 35.15787, 35.15286, 35.40105, 35.28883, 
    35.70983, 35.58942, 35.939, 35.85061, 35.93484, 35.90927, 35.93517, 
    35.80567, 35.86107, 35.74742, 35.30981, 35.4376, 35.05845, 34.83335, 
    34.68494, 34.5802, 34.59498, 34.62318, 34.76862, 34.90616, 35.01151, 
    35.08224, 35.15214, 35.365, 35.47839, 35.73426, 35.68786, 35.76649, 
    35.84183, 35.96887, 35.94791, 36.00405, 35.7644, 35.92341, 35.66148, 
    35.73284, 35.17124, 34.96061, 34.87169, 34.79408, 34.60635, 34.73584, 
    34.68471, 34.80651, 34.88423, 34.84576, 35.08418, 34.99121, 35.48513, 
    35.27113, 35.83303, 35.69738, 35.86566, 35.77964, 35.92722, 35.79436, 
    36.02497, 36.07548, 36.04095, 36.17384, 35.78701, 35.93485, 34.84468, 
    34.85095, 34.88018, 34.75196, 34.74414, 34.62725, 34.73122, 34.77564, 
    34.88874, 34.9559, 35.01992, 35.16126, 35.32012, 35.54401, 35.70615, 
    35.81544, 35.74836, 35.80758, 35.74139, 35.71043, 36.05655, 35.8616, 
    36.15468, 36.13837, 36.00539, 36.14021, 34.85536, 34.81929, 34.6945, 
    34.7921, 34.61456, 34.71379, 34.77103, 34.99316, 35.04223, 35.08783, 
    35.17815, 35.29456, 35.50014, 35.68045, 35.84622, 35.83403, 35.83832, 
    35.8755, 35.78352, 35.89064, 35.90867, 35.86156, 36.13618, 36.05741, 
    36.13802, 36.0867, 34.83101, 34.89175, 34.85891, 34.92071, 34.87716, 
    35.07144, 35.13, 35.40589, 35.29227, 35.47334, 35.31059, 35.33935, 
    35.4793, 35.31936, 35.67049, 35.4319, 35.87695, 35.63669, 35.89209, 
    35.8455, 35.92268, 35.99202, 36.07952, 36.24183, 36.20415, 36.3405, 
    34.9826, 35.06193, 35.05492, 35.13819, 35.19995, 35.33437, 35.55154, 
    35.46964, 35.6202, 35.65054, 35.42188, 35.56203, 35.11515, 35.18681, 
    35.14411, 34.98885, 35.48851, 35.23079, 35.70884, 35.5676, 35.98212, 
    35.7751, 36.18343, 36.36015, 36.52758, 36.7248, 35.10532, 35.05129, 
    35.1481, 35.28272, 35.40826, 35.5762, 35.59344, 35.62506, 35.70713, 
    35.77637, 35.63507, 35.79375, 35.20348, 35.511, 35.03091, 35.17449, 
    35.27475, 35.23071, 35.4603, 35.51473, 35.73721, 35.62194, 36.31643, 
    36.00671, 36.876, 36.62993, 35.03245, 35.10513, 35.35982, 35.2383, 
    35.58744, 35.67417, 35.74489, 35.83562, 35.84542, 35.89936, 35.81104, 
    35.89586, 35.57656, 35.71872, 35.33056, 35.42447, 35.38122, 35.33387, 
    35.48029, 35.6373, 35.64064, 35.69121, 35.83432, 35.58887, 36.35673, 
    35.87968, 35.18463, 35.32574, 35.34594, 35.29114, 35.66546, 35.52916, 
    35.89804, 35.79779, 35.96227, 35.8804, 35.86837, 35.76368, 35.69872, 
    35.5354, 35.40331, 35.29908, 35.32327, 35.43792, 35.64693, 35.84632, 
    35.80251, 35.94973, 35.56196, 35.72381, 35.66113, 35.8249, 35.46747, 
    35.77157, 35.39036, 35.42354, 35.52646, 35.73484, 35.78116, 35.83075, 
    35.80013, 35.65226, 35.62811, 35.52395, 35.49529, 35.41631, 35.35114, 
    35.41068, 35.47338, 35.65231, 35.81471, 35.99301, 36.03684, 36.24728, 
    36.07586, 36.35942, 36.11818, 36.53728, 35.78928, 36.11107, 35.53115, 
    35.59296, 35.70518, 35.96449, 35.82413, 35.98835, 35.62716, 35.44189, 
    35.39416, 35.3054, 35.39619, 35.3888, 35.47597, 35.44792, 35.65827, 
    35.54505, 35.86808, 35.98705, 36.32619, 36.53647, 36.75237, 36.84832, 
    36.87759, 36.88984,
  60.67866, 61.07138, 60.99464, 61.31427, 61.13654, 61.34644, 60.75787, 
    61.08709, 60.87651, 60.71379, 61.94415, 61.3286, 62.59654, 62.19429, 
    63.21474, 62.53363, 63.35389, 63.19484, 63.67592, 63.53733, 64.16097, 
    63.74009, 64.48915, 64.05992, 64.12669, 63.72631, 61.45146, 61.86686, 
    61.42703, 61.48588, 61.45945, 61.14022, 60.9806, 60.64882, 60.70879, 
    60.95258, 61.51238, 61.32119, 61.80522, 61.7942, 62.34192, 62.09377, 
    63.02899, 62.76031, 63.54311, 63.34439, 63.53375, 63.4762, 63.5345, 
    63.24357, 63.36789, 63.11309, 62.1401, 62.42293, 61.58691, 61.09489, 
    60.77224, 60.54533, 60.5773, 60.63837, 60.95401, 61.2537, 61.48405, 
    61.6391, 61.79262, 62.26212, 62.51342, 63.08363, 62.97991, 63.15579, 
    63.32469, 63.61038, 63.56317, 63.68969, 63.15111, 63.50803, 62.92099, 
    63.08046, 61.83464, 61.37265, 61.17846, 61.00938, 60.60192, 60.88274, 
    60.77174, 61.03644, 61.20583, 61.12193, 61.64335, 61.4396, 62.52837, 
    62.05472, 63.30494, 63.00117, 63.37819, 63.18523, 63.5166, 63.21821, 
    63.7369, 63.85101, 63.77299, 64.07372, 63.20175, 63.53376, 61.11959, 
    61.13326, 61.197, 60.91779, 60.90078, 60.64719, 60.87272, 60.96927, 
    61.21567, 61.36237, 61.50245, 61.81269, 62.16289, 62.65925, 63.02077, 
    63.26548, 63.11519, 63.24784, 63.0996, 63.03035, 63.80822, 63.36906, 
    64.03029, 63.99333, 63.69271, 63.99749, 61.14286, 61.06427, 60.79298, 
    61.00508, 60.61969, 60.83485, 60.95924, 61.44387, 61.55134, 61.65136, 
    61.84983, 62.10643, 62.56173, 62.96335, 63.33453, 63.30719, 63.31681, 
    63.40031, 63.19391, 63.43432, 63.47487, 63.36899, 63.98838, 63.81017, 
    63.99254, 63.87637, 61.08979, 61.22225, 61.1506, 61.28547, 61.19041, 
    61.6154, 61.74396, 62.35265, 62.10136, 62.5022, 62.14183, 62.20539, 
    62.51543, 62.16119, 62.9411, 62.41028, 63.40356, 62.86567, 63.43758, 
    63.33292, 63.50638, 63.66257, 63.86015, 64.22809, 64.14249, 64.45267, 
    61.42075, 61.59453, 61.57916, 61.76195, 61.89783, 62.19437, 62.67599, 
    62.494, 62.8289, 62.89658, 62.38808, 62.69933, 61.71135, 61.86889, 
    61.77497, 61.43444, 62.53588, 61.96577, 63.02679, 62.71173, 63.64025, 
    63.17506, 64.09548, 64.49747, 64.88044, 65.3342, 61.68975, 61.57121, 
    61.78375, 62.08028, 62.35789, 62.73087, 62.76926, 62.83974, 63.02298, 
    63.1779, 62.86208, 63.21685, 61.9056, 62.58585, 61.52654, 61.84178, 
    62.06271, 61.96557, 62.47326, 62.59414, 63.09025, 62.83279, 64.3978, 
    63.6957, 65.68405, 65.11556, 61.5299, 61.68932, 62.25066, 61.98231, 
    62.75591, 62.94933, 63.10743, 63.31075, 63.33276, 63.45393, 63.25561, 
    63.44606, 62.73167, 63.04889, 62.18595, 62.39381, 62.298, 62.19328, 
    62.51765, 62.86703, 62.87449, 62.9874, 63.30784, 62.75908, 64.48967, 
    63.4097, 61.8641, 62.17531, 62.21996, 62.09887, 62.92989, 62.62622, 
    63.45097, 63.22589, 63.59551, 63.4113, 63.38429, 63.14947, 63.00418, 
    62.64008, 62.34694, 62.1164, 62.16985, 62.42362, 62.88852, 63.33477, 
    63.23648, 63.56726, 62.69917, 63.06026, 62.92022, 63.2867, 62.48919, 
    63.16716, 62.31825, 62.39175, 62.62022, 63.08494, 63.18863, 63.2998, 
    63.23115, 62.90041, 62.84653, 62.61464, 62.55093, 62.37573, 62.23145, 
    62.36326, 62.5023, 62.90052, 63.26383, 63.6648, 63.7637, 64.24046, 
    63.85188, 64.4958, 63.9476, 64.90269, 63.20683, 63.93153, 62.63064, 
    62.7682, 63.0186, 63.60052, 63.28497, 63.6543, 62.84442, 62.43243, 
    62.32666, 62.13037, 62.33117, 62.31479, 62.50804, 62.4458, 62.91383, 
    62.66155, 63.38363, 63.65136, 64.42004, 64.90083, 65.39787, 65.61987, 
    65.68774, 65.71616,
  116.3177, 117.5456, 117.3041, 118.3152, 117.7513, 118.4177, 116.5638, 
    117.5952, 116.9339, 116.4268, 120.3482, 118.3608, 122.5137, 121.1711, 
    124.6258, 122.3021, 125.1096, 124.5568, 126.2418, 125.7524, 127.9808, 
    126.4695, 129.1813, 127.6151, 127.8565, 126.4205, 118.7533, 120.0957, 
    118.6751, 118.8636, 118.7789, 117.7629, 117.26, 116.2252, 116.4112, 
    117.1721, 118.9487, 118.3372, 119.895, 119.8592, 121.661, 120.8393, 
    123.9848, 123.0674, 125.7727, 125.0765, 125.7398, 125.5376, 125.7424, 
    124.7258, 125.1585, 124.2743, 120.992, 121.9312, 119.1884, 117.6198, 
    116.6085, 115.9053, 116.004, 116.1928, 117.1766, 118.1225, 118.8577, 
    119.3567, 119.854, 121.3958, 122.2342, 124.1728, 123.8164, 124.4217, 
    125.0078, 126.01, 125.8434, 126.2906, 124.4056, 125.6494, 123.6147, 
    124.1619, 119.9907, 118.5013, 117.8839, 117.3505, 116.0801, 116.9533, 
    116.607, 117.4356, 117.9707, 117.7052, 119.3704, 118.7153, 122.2845, 
    120.7108, 124.9391, 123.8893, 125.1945, 124.5236, 125.6795, 124.6378, 
    126.4582, 126.8648, 126.5865, 127.6649, 124.5808, 125.7399, 117.6978, 
    117.741, 117.9427, 117.063, 117.0098, 116.2202, 116.922, 117.2245, 
    118.0018, 118.4685, 118.9168, 119.9193, 121.0672, 122.7252, 123.9566, 
    124.8018, 124.2816, 124.7406, 124.2278, 123.9895, 126.712, 125.1626, 
    127.5082, 127.3751, 126.3013, 127.3901, 117.7713, 117.5232, 116.6731, 
    117.337, 116.135, 116.8037, 117.193, 118.729, 119.0739, 119.3963, 
    120.0402, 120.881, 122.3966, 123.7596, 125.0421, 124.9469, 124.9804, 
    125.2718, 124.5536, 125.3908, 125.5329, 125.1623, 127.3573, 126.719, 
    127.3722, 126.9554, 117.6037, 118.0227, 117.7958, 118.2235, 117.9218, 
    119.2802, 119.696, 121.6967, 120.8643, 122.1966, 120.9977, 121.2078, 
    122.241, 121.0616, 123.6834, 121.889, 125.2831, 123.4258, 125.4022, 
    125.0365, 125.6436, 126.1945, 126.8974, 128.2247, 127.9138, 129.0469, 
    118.655, 119.2129, 119.1634, 119.7544, 120.1968, 121.1713, 122.7818, 
    122.1691, 123.3005, 123.5312, 121.8149, 122.8607, 119.5903, 120.1023, 
    119.7967, 118.6988, 122.3097, 120.4189, 123.9772, 122.9027, 126.1155, 
    124.4884, 127.7436, 129.212, 130.6391, 132.3671, 119.5204, 119.1378, 
    119.8252, 120.7949, 121.7142, 122.9675, 123.0978, 123.3374, 123.9641, 
    124.4982, 123.4135, 124.6331, 120.2221, 122.4777, 118.9941, 120.014, 
    120.7371, 120.4183, 122.0996, 122.5056, 124.1956, 123.3137, 128.8452, 
    126.3119, 133.7281, 131.5293, 119.005, 119.5191, 121.3577, 120.4731, 
    123.0524, 123.7116, 124.2548, 124.9593, 125.0359, 125.4595, 124.7676, 
    125.4319, 122.9702, 124.0532, 121.1435, 121.834, 121.5149, 121.1677, 
    122.2484, 123.4304, 123.4559, 123.842, 124.9492, 123.0632, 129.1832, 
    125.3046, 120.0867, 121.1083, 121.256, 120.8561, 123.6451, 122.6137, 
    125.4491, 124.6645, 125.9575, 125.3102, 125.2158, 124.3999, 123.8996, 
    122.6605, 121.6777, 120.9138, 121.0902, 121.9335, 123.5037, 125.043, 
    124.7011, 125.8578, 122.8602, 124.0923, 123.612, 124.8756, 122.153, 
    124.4611, 121.5822, 121.8271, 122.5935, 124.1773, 124.5353, 124.9212, 
    124.6827, 123.5443, 123.3605, 122.5747, 122.3602, 121.7737, 121.2941, 
    121.7321, 122.197, 123.5447, 124.7961, 126.2024, 126.5535, 128.2698, 
    126.8678, 129.2059, 127.2107, 130.7229, 124.5984, 127.153, 122.6286, 
    123.0941, 123.9491, 125.9752, 124.8696, 126.1653, 123.3533, 121.963, 
    121.6102, 120.9599, 121.6252, 121.5707, 122.2162, 122.0077, 123.5902, 
    122.733, 125.2134, 126.1548, 128.9268, 130.7158, 132.6129, 133.4765, 
    133.7426, 133.8544,
  366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 366.0466, 
    366.0466, 366.0466,
  603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 603.5089, 
    603.5089, 603.5089,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOILPSI =
  -0.02127072, -0.02092213, -0.02098943, -0.02071172, -0.02086529, 
    -0.02068414, -0.02119956, -0.02090842, -0.02109379, -0.02123909, 
    -0.02018379, -0.02069942, -0.01966258, -0.01998089, -0.01919145, 
    -0.01971175, -0.01908832, -0.01920626, -0.01885362, -0.01895394, 
    -0.01851038, -0.01880751, -0.01828482, -0.01858088, -0.01853423, 
    -0.0188174, -0.02059455, -0.02024723, -0.02061532, -0.02056536, 
    -0.02058777, -0.0208621, -0.0210018, -0.02129762, -0.02124359, 
    -0.02102648, -0.02054294, -0.02070576, -0.02029802, -0.02030713, 
    -0.01986295, -0.02006194, -0.01933073, -0.01953564, -0.01894974, 
    -0.01909531, -0.01895655, -0.01899851, -0.018956, -0.01916998, 
    -0.01907798, -0.01926742, -0.02002451, -0.01979879, -0.02048009, 
    -0.02090163, -0.0211867, -0.02139147, -0.02136239, -0.02130708, 
    -0.02102522, -0.02076381, -0.0205669, -0.02043628, -0.02030844, 
    -0.01992659, -0.01972758, -0.01928958, -0.01936786, -0.01923544, 
    -0.01910985, -0.01890094, -0.01893516, -0.01884371, -0.01923893, 
    -0.0189753, -0.0194126, -0.01929194, -0.0202738, -0.0206617, -0.02082891, 
    -0.02097647, -0.02134006, -0.02108827, -0.02118715, -0.02095271, 
    -0.02080516, -0.020878, -0.02043272, -0.02060463, -0.01971585, 
    -0.0200936, -0.01912446, -0.01935177, -0.0190704, -0.01921343, 
    -0.01896904, -0.01918884, -0.0188098, -0.01872832, -0.01878396, 
    -0.0185712, -0.0192011, -0.01895655, -0.02088004, -0.02086814, 
    -0.0208128, -0.02105722, -0.02107227, -0.0212991, -0.02109715, 
    -0.02101176, -0.02079664, -0.02067049, -0.02055132, -0.02029185, 
    -0.02000616, -0.01961379, -0.01933694, -0.01915369, -0.01926584, 
    -0.01916679, -0.01927755, -0.0193297, -0.01875881, -0.01907713, 
    -0.01860165, -0.01862762, -0.01884154, -0.0186247, -0.02085979, 
    -0.02092834, -0.02116816, -0.02098023, -0.02132396, -0.02113083, 
    -0.02102061, -0.02060101, -0.02051002, -0.02042602, -0.02026119, 
    -0.0200517, -0.01968973, -0.01938043, -0.01910258, -0.01912279, 
    -0.01911567, -0.01905413, -0.01920695, -0.01902917, -0.0189995, 
    -0.01907717, -0.01863111, -0.0187574, -0.01862818, -0.01871029, 
    -0.02090603, -0.02079096, -0.02085306, -0.02073645, -0.02081853, 
    -0.02045617, -0.02034884, -0.01985445, -0.0200558, -0.01973637, 
    -0.02002311, -0.01997198, -0.01972602, -0.0200075, -0.01939734, 
    -0.01980881, -0.01905174, -0.01945485, -0.01902678, -0.01910377, 
    -0.01897648, -0.01886325, -0.01872182, -0.0184638, -0.01852321, 
    -0.01830962, -0.02062066, -0.02047369, -0.02048659, -0.02033387, 
    -0.0202217, -0.01998082, -0.01960079, -0.01974279, -0.01948294, 
    -0.01943121, -0.01982632, -0.01958273, -0.02037595, -0.02024552, 
    -0.02032307, -0.02060903, -0.01970997, -0.02016606, -0.0193324, 
    -0.01957312, -0.01887935, -0.01922104, -0.018556, -0.01827919, 
    -0.01802273, -0.01772784, -0.02039395, -0.02049328, -0.02031579, 
    -0.02007288, -0.01985027, -0.01955835, -0.01952874, -0.01947464, 
    -0.01933527, -0.0192189, -0.01945757, -0.01918985, -0.02021538, 
    -0.0196709, -0.02053097, -0.02026786, -0.02008712, -0.0201662, 
    -0.01975909, -0.01966441, -0.01928459, -0.01947996, -0.0183471, 
    -0.01883941, -0.01750678, -0.01786875, -0.02052811, -0.0203943, 
    -0.01993571, -0.02015253, -0.01953902, -0.01939107, -0.01927167, 
    -0.01912017, -0.01910389, -0.01901481, -0.01916102, -0.01902056, 
    -0.01955773, -0.01931572, -0.01998758, -0.0198218, -0.01989789, 
    -0.01998169, -0.01972423, -0.01945378, -0.01944806, -0.0193622, 
    -0.0191224, -0.01953658, -0.01828454, -0.01904731, -0.02024943, 
    -0.01999617, -0.01996029, -0.0200578, -0.01940585, -0.01963944, 
    -0.01901698, -0.01918311, -0.0189117, -0.01904606, -0.01906591, 
    -0.01924015, -0.01934949, -0.01962866, -0.01985897, -0.02004363, 
    -0.02000053, -0.01979824, -0.01943737, -0.01910242, -0.01917526, 
    -0.01893218, -0.01958284, -0.01930716, -0.01941321, -0.01913796, 
    -0.01974658, -0.019227, -0.01988176, -0.01982342, -0.01964411, 
    -0.0192886, -0.01921089, -0.01912826, -0.0191792, -0.0194283, 
    -0.01946945, -0.01964845, -0.01969817, -0.01983611, -0.01995107, 
    -0.019846, -0.01973629, -0.0194282, -0.01915493, -0.01886164, -0.0187906, 
    -0.01845528, -0.01872774, -0.01828038, -0.01865996, -0.01800811, 
    -0.01919736, -0.01867127, -0.01963599, -0.01952956, -0.01933861, 
    -0.0189081, -0.01913925, -0.01886922, -0.01947106, -0.01979129, 
    -0.01987507, -0.02003235, -0.01987149, -0.01988452, -0.01973176, 
    -0.01978072, -0.01941806, -0.01961198, -0.0190664, -0.01887134, 
    -0.01833187, -0.0180093, -0.01768718, -0.01754692, -0.01750447, 
    -0.01748675,
  -0.05475521, -0.05370497, -0.05390748, -0.05307256, -0.05353404, 
    -0.05298977, -0.05454059, -0.05366368, -0.05422177, -0.05465984, 
    -0.05149094, -0.05303564, -0.0499371, -0.05088531, -0.04853887, 
    -0.05008336, -0.04823363, -0.0485828, -0.04754012, -0.04783639, 
    -0.04652847, -0.04740404, -0.04586561, -0.04673604, -0.04659869, 
    -0.04743321, -0.05272097, -0.0516806, -0.05278328, -0.0526334, 
    -0.05270062, -0.05352443, -0.05394467, -0.05483643, -0.0546734, 
    -0.05401903, -0.05256615, -0.05305471, -0.0518327, -0.05185997, 
    -0.05053369, -0.05112718, -0.04895167, -0.04955984, -0.04782398, 
    -0.04825436, -0.04784409, -0.04796811, -0.04784248, -0.04847534, 
    -0.0482031, -0.04876401, -0.05101545, -0.05034252, -0.05237779, 
    -0.05364321, -0.05450179, -0.05511978, -0.05503197, -0.05486495, 
    -0.05401522, -0.05322906, -0.05263806, -0.05224659, -0.05186389, 
    -0.05072324, -0.0501305, -0.04882961, -0.04906178, -0.04866921, 
    -0.0482974, -0.04767982, -0.0477809, -0.04751085, -0.04867958, 
    -0.04789946, -0.04919453, -0.04883666, -0.05176004, -0.05292245, 
    -0.05342458, -0.05386848, -0.05496455, -0.05420512, -0.05450315, 
    -0.05379701, -0.0533533, -0.05357228, -0.05223593, -0.05275121, 
    -0.0500956, -0.05122168, -0.04834061, -0.04901404, -0.04818067, 
    -0.04860404, -0.04788099, -0.04853121, -0.04741079, -0.04717045, 
    -0.04733454, -0.04670758, -0.04856752, -0.04784406, -0.05357841, 
    -0.05354263, -0.05337628, -0.05411159, -0.05415694, -0.05484089, 
    -0.05423189, -0.05397471, -0.05332772, -0.05294884, -0.05259133, 
    -0.05181424, -0.05096066, -0.04979204, -0.04897008, -0.04842716, 
    -0.04875933, -0.04846594, -0.04879403, -0.04894863, -0.04726033, 
    -0.04820056, -0.04679721, -0.04687373, -0.04750444, -0.0468651, 
    -0.05351752, -0.05372368, -0.0544459, -0.05387983, -0.05491593, 
    -0.05433336, -0.05400132, -0.05274032, -0.05246754, -0.05221583, 
    -0.05172253, -0.05109662, -0.05001792, -0.04909903, -0.04827587, 
    -0.04833569, -0.04831462, -0.04813255, -0.04858484, -0.04805873, 
    -0.047971, -0.0482007, -0.04688398, -0.04725622, -0.04687535, 
    -0.04711733, -0.05365658, -0.05331064, -0.05349728, -0.05314687, 
    -0.05339345, -0.0523061, -0.05198468, -0.0505083, -0.05110884, 
    -0.05015668, -0.05101128, -0.05085872, -0.05012581, -0.05096473, 
    -0.04914917, -0.05037231, -0.04812549, -0.04931979, -0.04805168, 
    -0.0482794, -0.04790301, -0.04756852, -0.04715129, -0.04639152, 
    -0.0465663, -0.04593844, -0.05279932, -0.05235861, -0.05239731, 
    -0.05193996, -0.05160443, -0.05088511, -0.04975344, -0.05017585, 
    -0.04940332, -0.04924974, -0.05042459, -0.04969972, -0.05206589, 
    -0.05167559, -0.05190764, -0.05276437, -0.05007809, -0.0514381, 
    -0.04895661, -0.0496712, -0.04761605, -0.04862654, -0.0466628, 
    -0.04584904, -0.04509719, -0.04423486, -0.0521198, -0.05241737, 
    -0.05188587, -0.0511598, -0.0504959, -0.04962729, -0.04953935, 
    -0.04937868, -0.04896513, -0.04862025, -0.04932794, -0.0485342, 
    -0.0515854, -0.04996188, -0.05253029, -0.0517424, -0.05120232, 
    -0.05143856, -0.05022439, -0.04994264, -0.04881486, -0.04939448, 
    -0.04604843, -0.04749811, -0.04359022, -0.0446466, -0.05252175, 
    -0.05212085, -0.05075054, -0.05139772, -0.0495699, -0.04913061, 
    -0.0487766, -0.0483279, -0.04827977, -0.04801627, -0.04844885, 
    -0.0480333, -0.04962546, -0.04890715, -0.05090529, -0.05041109, 
    -0.05063783, -0.05088774, -0.05012061, -0.04931669, -0.04929976, 
    -0.04904497, -0.04833429, -0.04956264, -0.04586461, -0.04811219, 
    -0.05168737, -0.05093084, -0.05082386, -0.05111485, -0.04917447, 
    -0.04986835, -0.04802269, -0.04851426, -0.04771161, -0.04810868, 
    -0.04816739, -0.04868321, -0.04900728, -0.04983629, -0.0505218, 
    -0.05107255, -0.05094393, -0.0503409, -0.04926799, -0.04827537, 
    -0.04849096, -0.04777212, -0.04970009, -0.04888174, -0.0491963, 
    -0.04838059, -0.05018711, -0.04864405, -0.05058976, -0.05041593, 
    -0.04988223, -0.04882669, -0.04859652, -0.04835186, -0.04850269, 
    -0.04924108, -0.04936323, -0.04989515, -0.05004304, -0.05045373, 
    -0.05079641, -0.0504832, -0.05015645, -0.04924081, -0.04843079, 
    -0.04756376, -0.04735414, -0.04636636, -0.04716865, -0.04585239, 
    -0.04696874, -0.04505423, -0.04855633, -0.04700219, -0.04985812, 
    -0.0495418, -0.04897496, -0.0477009, -0.04838439, -0.04758612, 
    -0.04936803, -0.05032018, -0.05056981, -0.05103887, -0.05055914, 
    -0.05059798, -0.05014303, -0.05028876, -0.04921072, -0.04978672, 
    -0.04816884, -0.04759239, -0.04600379, -0.04505782, -0.04411625, 
    -0.0437072, -0.04358351, -0.04353191,
  -0.07892327, -0.07726903, -0.07758781, -0.0762741, -0.07700003, 
    -0.07614392, -0.07858502, -0.07720403, -0.07808273, -0.07877295, 
    -0.07378995, -0.07621606, -0.07135536, -0.07284038, -0.0691697, 
    -0.07158427, -0.06869322, -0.06923831, -0.06761158, -0.0680735, 
    -0.06603594, -0.06739948, -0.06500509, -0.06635902, -0.06614523, 
    -0.06744494, -0.0757214, -0.07408752, -0.07581934, -0.07558377, 
    -0.07568941, -0.0769849, -0.07764634, -0.07905132, -0.07879434, 
    -0.07776343, -0.07547809, -0.07624605, -0.07432629, -0.07436909, 
    -0.07228945, -0.07321952, -0.06981447, -0.07076519, -0.06805416, 
    -0.06872559, -0.06808552, -0.06827897, -0.068083, -0.06907053, 
    -0.0686456, -0.06952131, -0.07304436, -0.07199004, -0.07518217, 
    -0.07717179, -0.07852388, -0.07949811, -0.07935962, -0.07909628, 
    -0.07775743, -0.07652025, -0.0755911, -0.0749761, -0.07437524, 
    -0.07258637, -0.07165807, -0.06962378, -0.06998654, -0.06937324, 
    -0.06879277, -0.06782936, -0.06798698, -0.06756595, -0.06938946, 
    -0.06817187, -0.07019402, -0.0696348, -0.07421219, -0.07603811, 
    -0.07682776, -0.07752641, -0.0792533, -0.07805649, -0.07852602, 
    -0.07741389, -0.07671566, -0.0770602, -0.07495936, -0.07576893, 
    -0.07160343, -0.07336769, -0.06886021, -0.06991193, -0.0686106, 
    -0.06927148, -0.06814307, -0.06915776, -0.06740999, -0.0670355, 
    -0.06729116, -0.06631473, -0.06921446, -0.06808547, -0.07706985, 
    -0.07701354, -0.07675182, -0.07790919, -0.07798062, -0.07905836, 
    -0.07809868, -0.07769365, -0.07667544, -0.07607958, -0.07551767, 
    -0.07429729, -0.07295846, -0.0711284, -0.06984325, -0.06899531, 
    -0.06951401, -0.06905586, -0.06956821, -0.06980973, -0.06717552, 
    -0.06864162, -0.06645425, -0.06657339, -0.06755595, -0.06655996, 
    -0.07697403, -0.07729848, -0.07843582, -0.07754429, -0.07917666, 
    -0.07825851, -0.07773555, -0.07575179, -0.07532317, -0.07492779, 
    -0.07415338, -0.07317162, -0.07148186, -0.07004475, -0.06875917, 
    -0.06885254, -0.06881965, -0.06853551, -0.06924149, -0.06842034, 
    -0.06828347, -0.06864186, -0.06658936, -0.06716914, -0.06657592, 
    -0.06695276, -0.07719287, -0.07664856, -0.07694218, -0.07639097, 
    -0.07677883, -0.07506956, -0.07456483, -0.07224966, -0.07319078, 
    -0.07169907, -0.07303783, -0.0727987, -0.07165071, -0.07296486, 
    -0.07012309, -0.07203666, -0.06852449, -0.07038979, -0.06840932, 
    -0.06876468, -0.06817742, -0.06765584, -0.06700566, -0.06582288, 
    -0.06609484, -0.06511831, -0.07584454, -0.07515204, -0.07521285, 
    -0.07449465, -0.07396806, -0.07284007, -0.07106801, -0.07172909, 
    -0.07052042, -0.07028031, -0.07211858, -0.07098397, -0.07469233, 
    -0.0740797, -0.07444391, -0.07578961, -0.07157604, -0.0737071, 
    -0.06982219, -0.07093937, -0.06772994, -0.0693066, -0.06624503, 
    -0.06497931, -0.06381156, -0.0624741, -0.07477698, -0.07524436, 
    -0.07440975, -0.07327065, -0.07223026, -0.07087068, -0.07073314, 
    -0.07048189, -0.06983552, -0.06929679, -0.07040254, -0.06916243, 
    -0.07393815, -0.07139417, -0.07542175, -0.07418454, -0.07333734, 
    -0.07370784, -0.07180508, -0.07136407, -0.06960073, -0.0705066, 
    -0.06528925, -0.06754606, -0.06147569, -0.06311243, -0.07540835, 
    -0.07477865, -0.07262918, -0.07364379, -0.07078093, -0.07009412, 
    -0.06954098, -0.06884037, -0.06876525, -0.06835409, -0.06902918, 
    -0.06838066, -0.07086781, -0.06974492, -0.07287171, -0.07209742, 
    -0.07245259, -0.07284419, -0.07164261, -0.07038496, -0.07035851, 
    -0.06996026, -0.06885028, -0.07076957, -0.06500346, -0.06850368, 
    -0.0740982, -0.07291172, -0.07274409, -0.0732002, -0.07016265, 
    -0.0712478, -0.0683641, -0.0691313, -0.06787894, -0.06849827, 
    -0.06858987, -0.06939512, -0.06990137, -0.07119764, -0.07227083, 
    -0.07313389, -0.07293227, -0.07198751, -0.07030883, -0.06875837, 
    -0.06909491, -0.06797329, -0.07098456, -0.06970521, -0.07019676, 
    -0.06892261, -0.07174671, -0.0693339, -0.07237729, -0.07210502, 
    -0.07126952, -0.0696192, -0.06925974, -0.06887776, -0.06911324, 
    -0.07026678, -0.07045774, -0.07128975, -0.07152118, -0.07216422, 
    -0.07270107, -0.07221036, -0.07169871, -0.07026635, -0.06900097, 
    -0.06764842, -0.06732172, -0.06578372, -0.06703268, -0.06498447, 
    -0.06672126, -0.06374483, -0.06919695, -0.06677338, -0.0712318, 
    -0.07073697, -0.06985085, -0.06786221, -0.06892855, -0.06768326, 
    -0.07046524, -0.07195505, -0.07234604, -0.07308108, -0.07232933, 
    -0.07239018, -0.07167772, -0.07190588, -0.07021932, -0.07112009, 
    -0.06859213, -0.06769304, -0.06521988, -0.06375043, -0.06229033, 
    -0.06165679, -0.06146532, -0.06138545,
  -0.08614822, -0.08423896, -0.08460679, -0.08309133, -0.08392864, 
    -0.08294121, -0.08575772, -0.08416398, -0.08517794, -0.08597468, 
    -0.08022813, -0.0830244, -0.07742523, -0.07913451, -0.07491172, 
    -0.07768863, -0.07436414, -0.07499059, -0.07312156, -0.07365213, 
    -0.07131277, -0.072878, -0.07013018, -0.07168353, -0.07143818, 
    -0.07293019, -0.08245402, -0.08057093, -0.08256693, -0.08229534, 
    -0.08241714, -0.08391119, -0.08467433, -0.08629607, -0.08599936, 
    -0.08480944, -0.08217351, -0.08305899, -0.08084603, -0.08089534, 
    -0.07850024, -0.07957111, -0.07565293, -0.07674626, -0.07362992, 
    -0.07440133, -0.07366594, -0.07388817, -0.07366305, -0.07479773, 
    -0.07430942, -0.07531589, -0.0793694, -0.07815561, -0.08183239, 
    -0.08412679, -0.08568715, -0.08681199, -0.08665206, -0.08634797, 
    -0.08480252, -0.08337522, -0.08230379, -0.08159487, -0.08090243, 
    -0.07884206, -0.07777355, -0.07543368, -0.07585076, -0.07514568, 
    -0.07447852, -0.07337169, -0.07355274, -0.07306916, -0.07516432, 
    -0.07376513, -0.07608935, -0.07544635, -0.08071456, -0.08281919, 
    -0.08372992, -0.08453593, -0.08652929, -0.08514766, -0.0856896, 
    -0.08440612, -0.08360061, -0.08399805, -0.08157557, -0.08250882, 
    -0.07771068, -0.07974175, -0.07455603, -0.07576498, -0.0742692, 
    -0.07502871, -0.07373205, -0.074898, -0.07289007, -0.07246006, 
    -0.07275362, -0.07163269, -0.07496317, -0.07366588, -0.08400919, 
    -0.08394422, -0.08364232, -0.08497766, -0.08506008, -0.08630419, 
    -0.08519635, -0.08472892, -0.08355421, -0.08286703, -0.08221913, 
    -0.08081263, -0.07927049, -0.0771641, -0.07568601, -0.07471129, 
    -0.0753075, -0.07478088, -0.0753698, -0.07564747, -0.07262084, 
    -0.07430484, -0.07179283, -0.07192957, -0.07305768, -0.07191415, 
    -0.08389865, -0.08427295, -0.08558548, -0.08455656, -0.08644079, 
    -0.08538082, -0.08477727, -0.08248906, -0.08199492, -0.08153919, 
    -0.0806468, -0.07951594, -0.07757078, -0.0759177, -0.07443992, 
    -0.07454721, -0.07450942, -0.07418292, -0.07499424, -0.07405059, 
    -0.07389334, -0.07430512, -0.0719479, -0.0726135, -0.07193249, 
    -0.07236508, -0.08415111, -0.08352321, -0.0838619, -0.08322612, 
    -0.08367347, -0.08170259, -0.08112089, -0.07845444, -0.07953801, 
    -0.07782073, -0.07936188, -0.07908653, -0.07776508, -0.07927786, 
    -0.07600778, -0.07820927, -0.07417026, -0.07631449, -0.07403793, 
    -0.07444625, -0.07377151, -0.0731724, -0.07242581, -0.07106829, 
    -0.07138035, -0.07026003, -0.082596, -0.08179766, -0.08186775, 
    -0.08104002, -0.0804333, -0.07913416, -0.07709462, -0.07785529, 
    -0.07646473, -0.07618859, -0.07830356, -0.07699794, -0.08126783, 
    -0.08056192, -0.08098155, -0.08253267, -0.07767916, -0.08013269, 
    -0.0756618, -0.07694663, -0.07325751, -0.07506908, -0.0715527, 
    -0.07010062, -0.06876182, -0.06722952, -0.08136538, -0.08190408, 
    -0.08094219, -0.07962999, -0.07843211, -0.07686761, -0.0767094, 
    -0.07642041, -0.07567713, -0.0750578, -0.07632916, -0.07490336, 
    -0.08039885, -0.07746988, -0.08210856, -0.08068271, -0.0797068, 
    -0.08013354, -0.07794274, -0.07743525, -0.07540718, -0.07644883, 
    -0.07045611, -0.07304633, -0.06608645, -0.06796069, -0.0820931, 
    -0.0813673, -0.07889135, -0.08005976, -0.07676437, -0.07597446, 
    -0.07533851, -0.07453323, -0.0744469, -0.07397447, -0.07475021, 
    -0.074005, -0.07686431, -0.07557297, -0.07917059, -0.0782792, 
    -0.07868805, -0.0791389, -0.07775576, -0.07630894, -0.07627852, 
    -0.07582054, -0.07454462, -0.0767513, -0.07012832, -0.07414635, 
    -0.08058324, -0.07921667, -0.07902364, -0.07954886, -0.07605328, 
    -0.07730147, -0.07398597, -0.07486759, -0.07342865, -0.07414012, 
    -0.07424538, -0.07517082, -0.07575284, -0.07724375, -0.07847881, 
    -0.07947249, -0.07924032, -0.07815269, -0.07622138, -0.074439, 
    -0.07482576, -0.07353701, -0.07699861, -0.07552731, -0.0760925, 
    -0.07462774, -0.07787556, -0.07510046, -0.07860136, -0.07828794, 
    -0.07732646, -0.07542843, -0.07501521, -0.0745762, -0.07484683, 
    -0.07617301, -0.07639264, -0.07734973, -0.07761603, -0.07835609, 
    -0.07897411, -0.07840921, -0.07782032, -0.07617253, -0.07471779, 
    -0.07316388, -0.0727887, -0.07102335, -0.07245683, -0.07010654, 
    -0.07209932, -0.06868534, -0.07494304, -0.07215916, -0.07728305, 
    -0.07671381, -0.07569475, -0.07340942, -0.07463456, -0.07320389, 
    -0.07640126, -0.07811534, -0.07856539, -0.07941168, -0.07854614, 
    -0.07861619, -0.07779617, -0.07805874, -0.07611843, -0.07715453, 
    -0.07424798, -0.07321513, -0.07037654, -0.06869176, -0.06701908, 
    -0.06629374, -0.06607457, -0.06598315,
  -0.0672486, -0.0657028, -0.06600061, -0.0647736, -0.06545154, -0.06465206, 
    -0.06693244, -0.06564209, -0.06646304, -0.06710809, -0.06245528, 
    -0.06471941, -0.0601857, -0.06156976, -0.05815042, -0.06039899, 
    -0.05770702, -0.05821428, -0.05670086, -0.05713048, -0.05523624, 
    -0.05650363, -0.05427869, -0.05553645, -0.05533779, -0.0565459, 
    -0.06425758, -0.06273286, -0.06434901, -0.06412911, -0.06422772, 
    -0.06543741, -0.0660553, -0.0673683, -0.06712808, -0.06616469, 
    -0.06403046, -0.06474742, -0.0629556, -0.06299553, -0.06105617, 
    -0.06192328, -0.0587506, -0.05963592, -0.05711249, -0.05773713, 
    -0.05714166, -0.0573216, -0.05713932, -0.05805812, -0.05766271, 
    -0.05847768, -0.06175995, -0.06077711, -0.06375425, -0.06561197, 
    -0.0668753, -0.06778599, -0.06765652, -0.06741033, -0.06615909, 
    -0.06500345, -0.06413595, -0.06356194, -0.06300128, -0.06133295, 
    -0.06046775, -0.05857307, -0.0589108, -0.05833986, -0.05779964, 
    -0.0569034, -0.05705, -0.05665843, -0.05835495, -0.05722198, -0.05910399, 
    -0.05858333, -0.06284916, -0.06455325, -0.06529065, -0.06594324, 
    -0.06755712, -0.06643852, -0.0668773, -0.06583814, -0.06518595, 
    -0.06550774, -0.06354631, -0.06430195, -0.06041684, -0.06206146, 
    -0.0578624, -0.05884134, -0.05763014, -0.05824515, -0.05719519, 
    -0.05813931, -0.05651341, -0.05616523, -0.05640293, -0.05549529, 
    -0.05819207, -0.05714161, -0.06551675, -0.06546416, -0.06521972, 
    -0.06630088, -0.06636762, -0.06737487, -0.06647794, -0.06609949, 
    -0.06514838, -0.06459199, -0.0640674, -0.06292855, -0.06167986, 
    -0.05997426, -0.05877739, -0.05798812, -0.05847089, -0.05804447, 
    -0.05852134, -0.05874618, -0.05629541, -0.057659, -0.05562495, 
    -0.05573568, -0.05664914, -0.05572319, -0.06542726, -0.06573032, 
    -0.06679299, -0.06595995, -0.06748547, -0.0666273, -0.06613865, 
    -0.06428596, -0.06388585, -0.06351686, -0.06279428, -0.06187861, 
    -0.06030356, -0.058965, -0.05776838, -0.05785526, -0.05782466, 
    -0.05756028, -0.05821724, -0.05745313, -0.0573258, -0.05765922, 
    -0.05575052, -0.05628947, -0.05573803, -0.05608831, -0.06563167, 
    -0.06512328, -0.06539751, -0.06488274, -0.06524494, -0.06364916, 
    -0.06317817, -0.06101909, -0.06189648, -0.06050595, -0.06175387, 
    -0.0615309, -0.0604609, -0.06168583, -0.05903795, -0.06082057, 
    -0.05755003, -0.0592863, -0.05744288, -0.0577735, -0.05722714, 
    -0.05674203, -0.05613749, -0.05503828, -0.05529096, -0.05438383, 
    -0.06437254, -0.06372613, -0.06378289, -0.06311268, -0.06262141, 
    -0.06156947, -0.05991799, -0.06053393, -0.05940795, -0.05918434, 
    -0.06089691, -0.0598397, -0.06329714, -0.06272556, -0.06306534, 
    -0.06432126, -0.06039132, -0.062378, -0.05875779, -0.05979816, 
    -0.05681094, -0.05827783, -0.05543052, -0.05425476, -0.05317075, 
    -0.05193013, -0.06337613, -0.0638123, -0.06303346, -0.06197096, 
    -0.061001, -0.05973418, -0.05960607, -0.05937206, -0.05877019, 
    -0.0582687, -0.05929817, -0.05814365, -0.06259353, -0.06022185, 
    -0.06397787, -0.06282336, -0.06203315, -0.0623787, -0.06060474, 
    -0.06019381, -0.05855162, -0.05939507, -0.0545426, -0.05663994, 
    -0.05100467, -0.05252211, -0.06396536, -0.06337767, -0.06137286, 
    -0.06231895, -0.05965057, -0.05901096, -0.058496, -0.05784394, 
    -0.05777403, -0.05739149, -0.05801964, -0.05741621, -0.05973151, 
    -0.05868585, -0.06159898, -0.06087719, -0.06120824, -0.06157332, 
    -0.06045334, -0.0592818, -0.05925716, -0.05888633, -0.05785317, -0.05964, 
    -0.05427719, -0.05753067, -0.06274281, -0.06163628, -0.06147999, 
    -0.06190526, -0.05907478, -0.06008549, -0.0574008, -0.05811468, 
    -0.05694951, -0.05752562, -0.05761085, -0.05836022, -0.0588315, 
    -0.06003875, -0.06103882, -0.06184343, -0.06165543, -0.06077475, 
    -0.0592109, -0.05776764, -0.05808081, -0.05703726, -0.05984025, 
    -0.05864888, -0.05910654, -0.05792047, -0.06055035, -0.05830325, 
    -0.06113805, -0.06088427, -0.06010572, -0.05856882, -0.05823422, 
    -0.05787873, -0.05809787, -0.05917174, -0.05934957, -0.06012457, 
    -0.0603402, -0.06093945, -0.06143988, -0.06098246, -0.06050562, 
    -0.05917135, -0.05799338, -0.05673513, -0.05643133, -0.0550019, 
    -0.05616261, -0.05425955, -0.05587313, -0.05310883, -0.05817578, 
    -0.05592158, -0.06007058, -0.05960964, -0.05878447, -0.05693395, 
    -0.05792599, -0.05676753, -0.05935656, -0.06074451, -0.06110892, 
    -0.06179419, -0.06109335, -0.06115006, -0.06048606, -0.06069868, 
    -0.05912754, -0.05996651, -0.05761296, -0.05677662, -0.05447816, 
    -0.05311403, -0.05175973, -0.05117249, -0.05099505, -0.05092105,
  -0.0638878, -0.06219571, -0.06252145, -0.06118011, -0.06192097, 
    -0.06104734, -0.06354146, -0.06212931, -0.06302749, -0.06373387, 
    -0.05865141, -0.0611209, -0.05618335, -0.05768754, -0.0539767, 
    -0.05641496, -0.05349683, -0.05404584, -0.05240909, -0.05287335, 
    -0.05082871, -0.05219607, -0.04979745, -0.05115236, -0.05093816, 
    -0.05224172, -0.06061661, -0.05895377, -0.06071642, -0.06047637, 
    -0.06058401, -0.06190552, -0.06258129, -0.06401896, -0.06375577, 
    -0.06270097, -0.06036871, -0.0611515, -0.05919648, -0.05924, -0.05712904, 
    -0.0580722, -0.05462674, -0.05558664, -0.0528539, -0.05352941, 
    -0.05288543, -0.05307997, -0.0528829, -0.05387678, -0.05344889, 
    -0.05433109, -0.05789446, -0.05682575, -0.06006733, -0.06209638, 
    -0.06347889, -0.06447678, -0.06433484, -0.06406501, -0.06269485, 
    -0.06143122, -0.06048384, -0.05985754, -0.05924626, -0.05742998, 
    -0.05648965, -0.05443441, -0.05480035, -0.05418183, -0.05359704, 
    -0.05262792, -0.05278635, -0.05236326, -0.05419816, -0.05297226, 
    -0.05500976, -0.05444552, -0.05908049, -0.06093944, -0.06174509, 
    -0.06245869, -0.06422589, -0.06300066, -0.06348107, -0.06234372, 
    -0.06163065, -0.06198241, -0.0598405, -0.06066505, -0.05643435, 
    -0.05822259, -0.05366496, -0.05472507, -0.05341366, -0.05407926, 
    -0.0529433, -0.05396467, -0.05220662, -0.0518307, -0.05208732, 
    -0.05110797, -0.0540218, -0.05288538, -0.06199227, -0.06193476, 
    -0.06166755, -0.06285001, -0.06292305, -0.06402616, -0.06304381, 
    -0.06262964, -0.06158959, -0.06098174, -0.06040902, -0.05916701, 
    -0.05780732, -0.0559538, -0.05465577, -0.05380102, -0.05432373, 
    -0.05386201, -0.05437837, -0.05462196, -0.05197123, -0.05344488, 
    -0.05124779, -0.05136721, -0.05235322, -0.05135375, -0.06189442, 
    -0.0622258, -0.06338875, -0.06247697, -0.06414735, -0.06320732, 
    -0.06267248, -0.06064758, -0.06021091, -0.05980837, -0.05902069, 
    -0.05802358, -0.05631132, -0.05485909, -0.05356322, -0.05365723, 
    -0.05362411, -0.0533381, -0.05404904, -0.05322219, -0.0530845, 
    -0.05344512, -0.05138322, -0.05196482, -0.05136975, -0.05174769, 
    -0.06211792, -0.06156216, -0.0618619, -0.06129932, -0.06169512, 
    -0.05995268, -0.05943907, -0.05708873, -0.05804303, -0.05653114, 
    -0.05788784, -0.05764527, -0.0564822, -0.05781381, -0.05493817, 
    -0.05687296, -0.05332701, -0.05520742, -0.05321112, -0.05356877, 
    -0.05297784, -0.05245356, -0.05180077, -0.05061537, -0.05088769, 
    -0.0499106, -0.06074211, -0.06003665, -0.06009857, -0.05936769, 
    -0.05883235, -0.05768723, -0.05589274, -0.05656153, -0.05533936, 
    -0.05509688, -0.05695593, -0.05580777, -0.05956878, -0.05894582, 
    -0.05931609, -0.06068613, -0.05640663, -0.05856724, -0.05463453, 
    -0.05576269, -0.05252801, -0.05411466, -0.05103813, -0.04977169, 
    -0.04860622, -0.04727496, -0.05965491, -0.06013065, -0.05928134, 
    -0.0581241, -0.05706907, -0.05569325, -0.05555426, -0.05530043, 
    -0.05464798, -0.05410476, -0.0552203, -0.05396937, -0.05880198, 
    -0.0562226, -0.06031131, -0.05905238, -0.05819178, -0.05856799, 
    -0.05663846, -0.05619216, -0.05441117, -0.05532539, -0.05008151, 
    -0.05234329, -0.04628376, -0.04790984, -0.06029766, -0.05965659, 
    -0.05747338, -0.05850293, -0.05560255, -0.05490891, -0.05435093, 
    -0.05364498, -0.05356934, -0.05315554, -0.05383513, -0.05318227, 
    -0.05569036, -0.05455659, -0.05771932, -0.0569345, -0.05729437, 
    -0.05769141, -0.056474, -0.05520255, -0.05517584, -0.05477383, 
    -0.05365497, -0.05559107, -0.04979584, -0.05330606, -0.05896461, 
    -0.05775991, -0.05758988, -0.05805259, -0.05497809, -0.05607455, 
    -0.05316561, -0.05393801, -0.05267775, -0.05330061, -0.0533928, 
    -0.05420387, -0.05471441, -0.05602381, -0.05711018, -0.05798529, 
    -0.05778074, -0.05682318, -0.05512566, -0.05356242, -0.05390135, 
    -0.05277259, -0.05580836, -0.05451654, -0.05501252, -0.05372779, 
    -0.05657937, -0.05414218, -0.05721806, -0.05694219, -0.05609652, 
    -0.0544298, -0.05406743, -0.05368263, -0.05391981, -0.05508321, 
    -0.05527604, -0.05611697, -0.05635111, -0.05700216, -0.05754626, 
    -0.05704891, -0.05653078, -0.05508278, -0.05380671, -0.05244611, 
    -0.05211799, -0.05057618, -0.05182788, -0.04977685, -0.05151549, 
    -0.04853971, -0.05400416, -0.05156777, -0.05605836, -0.05555813, 
    -0.05466345, -0.05266094, -0.05373377, -0.05248111, -0.05528362, 
    -0.05679032, -0.05718638, -0.05793171, -0.05716945, -0.05723111, 
    -0.05650954, -0.05674052, -0.05503529, -0.05594539, -0.05339507, 
    -0.05249094, -0.05001215, -0.04854529, -0.04709235, -0.04646339, 
    -0.04627347, -0.04619428,
  -0.04035017, -0.03907184, -0.03931778, -0.03830553, -0.03886447, 
    -0.0382054, -0.04008836, -0.03902173, -0.03969999, -0.0402338, 
    -0.03640078, -0.03826088, -0.03454657, -0.03567605, -0.0328932, 
    -0.03472036, -0.03253425, -0.03294493, -0.03172141, -0.03206819, 
    -0.03054259, -0.03156237, -0.0297748, -0.03078379, -0.03062415, 
    -0.03159644, -0.03788066, -0.03662828, -0.0379559, -0.03777496, 
    -0.03785609, -0.03885281, -0.03936297, -0.04044933, -0.04025035, 
    -0.03945336, -0.03769382, -0.03828395, -0.03681095, -0.03684371, 
    -0.03525646, -0.03596519, -0.0333798, -0.03409905, -0.03205366, 
    -0.03255861, -0.03207722, -0.0322226, -0.03207533, -0.03281844, 
    -0.0324984, -0.03315843, -0.03583157, -0.0350287, -0.03746673, 
    -0.03899687, -0.04004107, -0.04079557, -0.04068821, -0.04048416, 
    -0.03944873, -0.03849493, -0.03778059, -0.03730871, -0.03684842, 
    -0.03548251, -0.03477641, -0.03323578, -0.03350982, -0.03304671, 
    -0.03260919, -0.03188484, -0.03200319, -0.03168719, -0.03305893, 
    -0.03214211, -0.03366669, -0.0332441, -0.03672365, -0.03812404, 
    -0.03873174, -0.0392704, -0.04060581, -0.03967972, -0.04004272, 
    -0.03918359, -0.03864539, -0.03891084, -0.03729587, -0.03791717, 
    -0.03473491, -0.03607827, -0.03265998, -0.03345343, -0.03247205, 
    -0.03296995, -0.03212046, -0.0328842, -0.03157025, -0.03128969, 
    -0.03148119, -0.0307507, -0.03292695, -0.03207719, -0.03891828, 
    -0.03887488, -0.03867324, -0.03956592, -0.0396211, -0.04045478, 
    -0.03971232, -0.03939948, -0.03861441, -0.03815594, -0.0377242, 
    -0.03678877, -0.03576607, -0.03437437, -0.03340153, -0.03276176, 
    -0.03315292, -0.03280739, -0.03319383, -0.03337621, -0.03139455, 
    -0.0324954, -0.03085493, -0.03094397, -0.03167969, -0.03093393, 
    -0.03884443, -0.03909456, -0.03997295, -0.03928419, -0.04054642, 
    -0.03983586, -0.03943183, -0.03790401, -0.03757491, -0.03727167, 
    -0.03667865, -0.03592864, -0.03464259, -0.03355382, -0.03258389, 
    -0.0326542, -0.03262943, -0.03241555, -0.03294734, -0.03232891, 
    -0.03222599, -0.03249558, -0.03095591, -0.03138977, -0.03094587, 
    -0.03122775, -0.03901313, -0.03859372, -0.03881989, -0.03839545, 
    -0.03869404, -0.03738037, -0.03699358, -0.03522618, -0.03594326, 
    -0.03480756, -0.03582659, -0.03564429, -0.03477082, -0.03577095, 
    -0.03361305, -0.03506416, -0.03240727, -0.0338148, -0.03232063, 
    -0.03258804, -0.03214628, -0.03175462, -0.03126735, -0.03038366, 
    -0.03058653, -0.02985898, -0.03797527, -0.03744363, -0.03749027, 
    -0.03693983, -0.03653692, -0.03567582, -0.03432857, -0.03483037, 
    -0.03391368, -0.03373196, -0.03512646, -0.03426485, -0.03709124, 
    -0.0366223, -0.03690099, -0.03793306, -0.03471411, -0.03633747, 
    -0.03338563, -0.03423104, -0.03181022, -0.03299643, -0.03069865, 
    -0.02975564, -0.0288894, -0.02790193, -0.03715609, -0.03751444, 
    -0.03687483, -0.0360042, -0.03521141, -0.03417898, -0.03407476, 
    -0.0338845, -0.0333957, -0.03298903, -0.03382445, -0.03288772, 
    -0.03651407, -0.03457602, -0.03765057, -0.0367025, -0.0360551, 
    -0.03633804, -0.03488811, -0.03455318, -0.03321838, -0.03390321, 
    -0.02998617, -0.03167228, -0.02716813, -0.02837259, -0.03764028, 
    -0.03715736, -0.03551513, -0.0362891, -0.03411097, -0.03359114, 
    -0.03317328, -0.03264504, -0.03258847, -0.03227909, -0.03278728, 
    -0.03229907, -0.03417681, -0.03332726, -0.03569993, -0.03511037, 
    -0.03538064, -0.03567896, -0.03476467, -0.03381115, -0.03379113, 
    -0.03348995, -0.03265251, -0.03410237, -0.0297736, -0.03239161, 
    -0.03663645, -0.03573044, -0.03560267, -0.03595044, -0.03364296, 
    -0.03446495, -0.03228661, -0.03286425, -0.03192206, -0.03238753, 
    -0.03245645, -0.0330632, -0.03344545, -0.03442689, -0.03524229, 
    -0.03589985, -0.03574609, -0.03502678, -0.03375353, -0.03258329, 
    -0.03283682, -0.03199291, -0.03426529, -0.03329727, -0.03366876, 
    -0.03270698, -0.03484375, -0.03301704, -0.03532331, -0.03511614, 
    -0.03448142, -0.03323233, -0.03296109, -0.0326732, -0.03285063, 
    -0.03372172, -0.03386622, -0.03449677, -0.03467245, -0.03516117, 
    -0.03556988, -0.03519628, -0.03480728, -0.0337214, -0.03276602, 
    -0.03174906, -0.03150408, -0.03035447, -0.03128758, -0.02975948, 
    -0.03105455, -0.02884002, -0.03291374, -0.03109354, -0.0344528, 
    -0.03407767, -0.03340728, -0.03190951, -0.03271146, -0.0317752, 
    -0.0338719, -0.0350021, -0.03529953, -0.03585957, -0.03528681, 
    -0.03533312, -0.03479134, -0.03496472, -0.03368582, -0.03436807, 
    -0.03245816, -0.03178254, -0.02993454, -0.02884416, -0.02776664, 
    -0.02730101, -0.02716052, -0.02710195,
  -0.01970495, -0.01870051, -0.01889313, -0.01810233, -0.01853834, 
    -0.01802441, -0.01949858, -0.0186613, -0.01919307, -0.01961318, 
    -0.01662921, -0.01806758, -0.01521542, -0.01607413, -0.01397334, 
    -0.01534703, -0.01370616, -0.01401192, -0.01310461, -0.01336065, 
    -0.01224113, -0.01298748, -0.01168475, -0.01241691, -0.01230052, 
    -0.01301256, -0.01777202, -0.01680408, -0.01783044, -0.01768999, 
    -0.01775294, -0.01852923, -0.01892854, -0.0197832, -0.01962623, 
    -0.01899943, -0.01762706, -0.01808554, -0.01694472, -0.01696996, 
    -0.0157542, -0.01629521, -0.01433697, -0.01487742, -0.01334991, 
    -0.01372426, -0.01336733, -0.01347495, -0.01336593, -0.01391762, 
    -0.01367953, -0.01417134, -0.01619298, -0.015581, -0.01745114, 
    -0.01864185, -0.01946134, -0.02005678, -0.01997189, -0.01981069, 
    -0.0189958, -0.0182499, -0.01769435, -0.01732889, -0.01697359, 
    -0.01592643, -0.01538952, -0.01422918, -0.01443441, -0.01408788, 
    -0.01376187, -0.01322516, -0.01331259, -0.01307939, -0.01409701, 
    -0.01341534, -0.01455213, -0.0142354, -0.01687748, -0.01796112, 
    -0.01843466, -0.01885599, -0.01990677, -0.01917714, -0.01946264, 
    -0.01878799, -0.01836725, -0.01857458, -0.01731896, -0.01780037, 
    -0.01535806, -0.0163818, -0.01379965, -0.01439214, -0.01365996, 
    -0.01403058, -0.01339933, -0.01396663, -0.01299328, -0.01278711, 
    -0.01292777, -0.01239277, -0.0139985, -0.0133673, -0.0185804, 
    -0.01854647, -0.01838898, -0.01908777, -0.01913109, -0.0197875, 
    -0.01920275, -0.01895718, -0.01834308, -0.01798592, -0.01765062, 
    -0.01692763, -0.01614291, -0.01508521, -0.01435325, -0.0138754, 
    -0.01416722, -0.01390938, -0.0141978, -0.01433429, -0.0128641, 
    -0.0136773, -0.01246885, -0.01253391, -0.01307387, -0.01252657, 
    -0.01852268, -0.01871829, -0.01940772, -0.0188668, -0.01985986, 
    -0.01929986, -0.01898255, -0.01779014, -0.01753491, -0.01730026, 
    -0.01684284, -0.01626723, -0.01528811, -0.01446741, -0.01374306, 
    -0.01379535, -0.01377692, -0.01361802, -0.01401371, -0.01355374, 
    -0.01347746, -0.01367744, -0.01254264, -0.01286059, -0.0125353, 
    -0.01274168, -0.01865457, -0.01832693, -0.0185035, -0.01817236, 
    -0.01840522, -0.01738431, -0.01708551, -0.01573116, -0.01627842, 
    -0.01541313, -0.01618917, -0.01604987, -0.01538528, -0.01614663, 
    -0.01451186, -0.01560794, -0.01361187, -0.01466342, -0.0135476, 
    -0.01374614, -0.01341843, -0.01312909, -0.01277073, -0.01212556, 
    -0.01227312, -0.01174552, -0.01784549, -0.01743325, -0.01746936, 
    -0.01704405, -0.01673382, -0.01607395, -0.01505061, -0.01543043, 
    -0.0147378, -0.01460116, -0.0156553, -0.0150025, -0.01716087, 
    -0.01679948, -0.0170141, -0.0178127, -0.01534229, -0.01658059, 
    -0.01434134, -0.01497698, -0.0131701, -0.01405035, -0.01235481, 
    -0.01167093, -0.01104941, -0.0103492, -0.01721095, -0.01748808, 
    -0.01699394, -0.01632508, -0.01571992, -0.0149377, -0.01485912, 
    -0.01471585, -0.01434888, -0.01404482, -0.01467068, -0.01396925, 
    -0.01671625, -0.01523771, -0.01759354, -0.01686119, -0.01636406, 
    -0.01658102, -0.01547424, -0.01522042, -0.01421617, -0.01472993, 
    -0.01183743, -0.0130684, -0.009834953, -0.01068181, -0.01758556, 
    -0.01721193, -0.0159513, -0.01654346, -0.01488641, -0.01449541, 
    -0.01418244, -0.01378853, -0.01374646, -0.0135168, -0.01389441, 
    -0.01353161, -0.01493606, -0.01429764, -0.01609237, -0.01564306, 
    -0.01584878, -0.01607635, -0.01538061, -0.01466068, -0.01464562, 
    -0.01441952, -0.01379409, -0.01487992, -0.01168389, -0.01360025, 
    -0.01681037, -0.01611568, -0.0160181, -0.01628392, -0.01453431, 
    -0.01515368, -0.01352238, -0.01395176, -0.01325265, -0.01359722, 
    -0.01364838, -0.0141002, -0.01438616, -0.0151249, -0.01574342, 
    -0.01624521, -0.01612764, -0.01557954, -0.01461737, -0.01374261, 
    -0.01393131, -0.01330499, -0.01500283, -0.01427519, -0.01455368, 
    -0.01383462, -0.01544059, -0.01406572, -0.01580511, -0.01564746, 
    -0.01516614, -0.0142266, -0.01402398, -0.01380948, -0.01394161, 
    -0.01459346, -0.0147021, -0.01517775, -0.01531073, -0.0156817, 
    -0.01599308, -0.01570841, -0.01541293, -0.01459322, -0.01387857, 
    -0.01312499, -0.0129446, -0.01210436, -0.01278557, -0.0116737, 
    -0.0126148, -0.01101418, -0.01398866, -0.01264334, -0.0151445, 
    -0.01486131, -0.01435756, -0.01324338, -0.01383795, -0.01314426, 
    -0.01470637, -0.01556079, -0.01578699, -0.0162144, -0.01577731, 
    -0.01581258, -0.01540083, -0.0155324, -0.01456649, -0.01508045, 
    -0.01364964, -0.01314967, -0.01180011, -0.01101713, -0.01025399, 
    -0.009927681, -0.009829647, -0.009788836,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, 
    -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659, -0.0008999659,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15,
  -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, 
    -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15, -15 ;

 SOILWATER_10CM =
  363.8103, 365.636, 365.2806, 366.7545, 365.9372, 366.9021, 364.1799, 
    365.7088, 364.7322, 363.9743, 369.6232, 366.8203, 372.5483, 370.75, 
    375.2776, 372.2682, 375.8862, 375.1903, 377.2867, 376.6854, 379.3756, 
    377.5645, 380.7745, 378.9424, 379.2288, 377.5049, 367.383, 369.2736, 
    367.2712, 367.5403, 367.4195, 365.9542, 365.2156, 363.6708, 363.9509, 
    365.0855, 367.6614, 366.7862, 368.994, 368.944, 371.412, 370.2979, 
    374.4618, 373.2752, 376.7104, 375.8447, 376.6698, 376.4194, 376.6731, 
    375.4038, 375.9473, 374.8316, 370.5064, 371.7743, 368.0014, 365.7449, 
    364.2469, 363.1865, 363.3363, 363.622, 365.0922, 366.4763, 367.5319, 
    368.2391, 368.9368, 371.0547, 372.1781, 374.7022, 374.2456, 375.0191, 
    375.7586, 377.0026, 376.7976, 377.3464, 374.9985, 376.558, 373.9857, 
    374.6882, 369.1276, 367.0222, 366.1305, 365.3489, 363.4515, 364.7612, 
    364.2445, 365.4742, 366.2563, 365.8698, 368.2585, 367.3287, 372.2448, 
    370.122, 375.6723, 374.3393, 375.9922, 375.1481, 376.5952, 375.2927, 
    377.5508, 378.0437, 377.7068, 379.0016, 375.2206, 376.6699, 365.859, 
    365.9221, 366.2156, 364.924, 364.845, 363.6632, 364.7146, 365.163, 
    366.3015, 366.975, 367.616, 369.0279, 370.609, 372.827, 374.4256, 
    375.4997, 374.8408, 375.4225, 374.7723, 374.4677, 377.859, 375.9524, 
    378.8152, 378.6564, 377.3595, 378.6743, 365.9663, 365.6031, 364.3435, 
    365.329, 363.5346, 364.5385, 365.1165, 367.3483, 367.8392, 368.295, 
    369.1962, 370.3549, 372.3933, 374.1727, 375.8016, 375.6821, 375.7242, 
    376.0887, 375.1862, 376.237, 376.4137, 375.9521, 378.6352, 377.8674, 
    378.653, 378.153, 365.7212, 366.3318, 366.002, 366.6223, 366.1853, 
    368.1313, 368.7161, 371.4601, 370.3321, 372.1281, 370.5142, 370.7999, 
    372.1872, 370.6013, 374.0746, 371.7179, 376.1029, 373.7416, 376.2512, 
    375.7946, 376.5508, 377.2289, 378.083, 379.6626, 379.2964, 380.6196, 
    367.2425, 368.0362, 367.9661, 368.7977, 369.4135, 370.7504, 372.9013, 
    372.0915, 373.5789, 373.878, 371.6185, 373.0049, 368.5678, 369.2826, 
    368.8568, 367.3051, 372.2782, 369.7207, 374.4521, 373.0599, 377.1322, 
    375.1036, 379.095, 380.8099, 382.4183, 384.3004, 368.4696, 367.9298, 
    368.8966, 370.2372, 371.4835, 373.1448, 373.3149, 373.6268, 374.4353, 
    375.116, 373.7256, 375.2867, 369.4488, 372.5007, 367.726, 369.1598, 
    370.1581, 369.7197, 371.9989, 372.5375, 374.7312, 373.5961, 380.3864, 
    377.3725, 385.7368, 383.3962, 367.7413, 368.4677, 371.0031, 369.7953, 
    373.2557, 374.1108, 374.8066, 375.6977, 375.7938, 376.3225, 375.4565, 
    376.2882, 373.1483, 374.5493, 370.7125, 371.6441, 371.2153, 370.7454, 
    372.1969, 373.7476, 373.7804, 374.2786, 375.6853, 373.2698, 380.777, 
    376.13, 369.2608, 370.6648, 370.8653, 370.3209, 374.025, 372.6801, 
    376.3095, 375.3264, 376.9381, 376.1367, 376.0189, 374.9913, 374.3525, 
    372.7418, 371.4345, 370.3997, 370.6402, 371.7773, 373.8425, 375.8027, 
    375.3728, 376.8154, 373.0042, 374.5994, 373.9824, 375.5925, 372.07, 
    375.0692, 371.306, 371.6349, 372.6535, 374.708, 375.1631, 375.6499, 
    375.3494, 373.8949, 373.6569, 372.6286, 372.3452, 371.5633, 370.9168, 
    371.5075, 372.1285, 373.8954, 375.4925, 377.2386, 377.6666, 379.7156, 
    378.0475, 380.8031, 378.4601, 382.5114, 375.243, 378.3908, 372.6998, 
    373.3102, 374.4161, 376.96, 375.5849, 377.1932, 373.6475, 371.8168, 
    371.3437, 370.4627, 371.3638, 371.2905, 372.1541, 371.8764, 373.9542, 
    372.8371, 376.016, 377.1804, 380.4809, 382.5034, 384.5626, 385.4741, 
    385.7518, 385.8679 ;

 SOMC_FIRE =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SOMHR =
  6.191113e-08, 6.218415e-08, 6.213108e-08, 6.235129e-08, 6.222914e-08, 
    6.237333e-08, 6.196649e-08, 6.219499e-08, 6.204912e-08, 6.193572e-08, 
    6.277865e-08, 6.236112e-08, 6.321246e-08, 6.294614e-08, 6.361521e-08, 
    6.317101e-08, 6.370478e-08, 6.360241e-08, 6.391058e-08, 6.382229e-08, 
    6.421644e-08, 6.395133e-08, 6.44208e-08, 6.415313e-08, 6.4195e-08, 
    6.394257e-08, 6.244515e-08, 6.272666e-08, 6.242847e-08, 6.246862e-08, 
    6.24506e-08, 6.223166e-08, 6.212131e-08, 6.189027e-08, 6.193222e-08, 
    6.210192e-08, 6.248666e-08, 6.235607e-08, 6.268525e-08, 6.267781e-08, 
    6.304429e-08, 6.287905e-08, 6.349508e-08, 6.331999e-08, 6.382597e-08, 
    6.369872e-08, 6.382e-08, 6.378323e-08, 6.382047e-08, 6.363384e-08, 
    6.37138e-08, 6.354958e-08, 6.290999e-08, 6.309795e-08, 6.253738e-08, 
    6.220033e-08, 6.197651e-08, 6.181767e-08, 6.184013e-08, 6.188293e-08, 
    6.210291e-08, 6.230976e-08, 6.246739e-08, 6.257284e-08, 6.267674e-08, 
    6.299121e-08, 6.31577e-08, 6.353047e-08, 6.346321e-08, 6.357717e-08, 
    6.368606e-08, 6.386886e-08, 6.383878e-08, 6.391931e-08, 6.357418e-08, 
    6.380355e-08, 6.34249e-08, 6.352845e-08, 6.270493e-08, 6.23913e-08, 
    6.225795e-08, 6.214128e-08, 6.185739e-08, 6.205343e-08, 6.197615e-08, 
    6.216003e-08, 6.227686e-08, 6.221908e-08, 6.257572e-08, 6.243706e-08, 
    6.316757e-08, 6.285291e-08, 6.367335e-08, 6.347702e-08, 6.372042e-08, 
    6.359622e-08, 6.380903e-08, 6.361751e-08, 6.394929e-08, 6.402153e-08, 
    6.397217e-08, 6.416183e-08, 6.360688e-08, 6.381999e-08, 6.221745e-08, 
    6.222687e-08, 6.227079e-08, 6.207778e-08, 6.206597e-08, 6.188912e-08, 
    6.204649e-08, 6.21135e-08, 6.228363e-08, 6.238426e-08, 6.247993e-08, 
    6.269027e-08, 6.292518e-08, 6.32537e-08, 6.348974e-08, 6.364797e-08, 
    6.355095e-08, 6.363661e-08, 6.354085e-08, 6.349597e-08, 6.399446e-08, 
    6.371454e-08, 6.413455e-08, 6.411131e-08, 6.392123e-08, 6.411393e-08, 
    6.22335e-08, 6.217927e-08, 6.199097e-08, 6.213833e-08, 6.186986e-08, 
    6.202013e-08, 6.210653e-08, 6.243995e-08, 6.251322e-08, 6.258114e-08, 
    6.271532e-08, 6.288751e-08, 6.318957e-08, 6.345243e-08, 6.36924e-08, 
    6.367481e-08, 6.3681e-08, 6.373461e-08, 6.360182e-08, 6.375641e-08, 
    6.378234e-08, 6.371452e-08, 6.410819e-08, 6.399572e-08, 6.411081e-08, 
    6.403759e-08, 6.21969e-08, 6.228814e-08, 6.223884e-08, 6.233156e-08, 
    6.226623e-08, 6.255671e-08, 6.264381e-08, 6.305137e-08, 6.288411e-08, 
    6.315032e-08, 6.291116e-08, 6.295353e-08, 6.315899e-08, 6.292409e-08, 
    6.343792e-08, 6.308954e-08, 6.373669e-08, 6.338875e-08, 6.375849e-08, 
    6.369136e-08, 6.380252e-08, 6.390207e-08, 6.402733e-08, 6.425844e-08, 
    6.420493e-08, 6.439821e-08, 6.242419e-08, 6.254255e-08, 6.253214e-08, 
    6.265601e-08, 6.274763e-08, 6.294621e-08, 6.326471e-08, 6.314495e-08, 
    6.336484e-08, 6.340898e-08, 6.307491e-08, 6.328001e-08, 6.262177e-08, 
    6.272811e-08, 6.26648e-08, 6.243353e-08, 6.317253e-08, 6.279325e-08, 
    6.349364e-08, 6.328816e-08, 6.388787e-08, 6.358961e-08, 6.417547e-08, 
    6.44259e-08, 6.466167e-08, 6.493715e-08, 6.260716e-08, 6.252674e-08, 
    6.267075e-08, 6.286999e-08, 6.305489e-08, 6.33007e-08, 6.332585e-08, 
    6.33719e-08, 6.349119e-08, 6.359149e-08, 6.338645e-08, 6.361663e-08, 
    6.275275e-08, 6.320546e-08, 6.249633e-08, 6.270984e-08, 6.285825e-08, 
    6.279316e-08, 6.313125e-08, 6.321094e-08, 6.353477e-08, 6.336737e-08, 
    6.436409e-08, 6.392309e-08, 6.514694e-08, 6.480489e-08, 6.249864e-08, 
    6.260689e-08, 6.298366e-08, 6.280439e-08, 6.331711e-08, 6.344332e-08, 
    6.354593e-08, 6.367708e-08, 6.369125e-08, 6.376896e-08, 6.364161e-08, 
    6.376393e-08, 6.330121e-08, 6.350799e-08, 6.29406e-08, 6.307869e-08, 
    6.301516e-08, 6.294548e-08, 6.316055e-08, 6.338968e-08, 6.339459e-08, 
    6.346806e-08, 6.367506e-08, 6.331919e-08, 6.442097e-08, 6.374049e-08, 
    6.272494e-08, 6.293345e-08, 6.296325e-08, 6.288247e-08, 6.343066e-08, 
    6.323202e-08, 6.376707e-08, 6.362246e-08, 6.38594e-08, 6.374166e-08, 
    6.372434e-08, 6.357312e-08, 6.347897e-08, 6.324113e-08, 6.304762e-08, 
    6.289419e-08, 6.292986e-08, 6.309841e-08, 6.34037e-08, 6.369253e-08, 
    6.362925e-08, 6.384139e-08, 6.327993e-08, 6.351534e-08, 6.342435e-08, 
    6.366162e-08, 6.314175e-08, 6.35844e-08, 6.302862e-08, 6.307734e-08, 
    6.322809e-08, 6.35313e-08, 6.359841e-08, 6.367004e-08, 6.362585e-08, 
    6.341145e-08, 6.337633e-08, 6.322442e-08, 6.318248e-08, 6.306674e-08, 
    6.297091e-08, 6.305846e-08, 6.31504e-08, 6.341154e-08, 6.364689e-08, 
    6.390349e-08, 6.39663e-08, 6.426609e-08, 6.402202e-08, 6.442477e-08, 
    6.408233e-08, 6.467514e-08, 6.361008e-08, 6.407228e-08, 6.323495e-08, 
    6.332515e-08, 6.34883e-08, 6.386253e-08, 6.366051e-08, 6.389678e-08, 
    6.337496e-08, 6.310422e-08, 6.303419e-08, 6.290352e-08, 6.303718e-08, 
    6.302631e-08, 6.315422e-08, 6.311311e-08, 6.342022e-08, 6.325525e-08, 
    6.37239e-08, 6.389492e-08, 6.437795e-08, 6.467408e-08, 6.497555e-08, 
    6.510865e-08, 6.514917e-08, 6.51661e-08 ;

 SOM_C_LEACHED =
  6.657648e-21, 3.039822e-20, 5.200039e-20, -2.03758e-20, 5.574121e-20, 
    1.492206e-20, -1.561889e-20, 4.428614e-20, -8.652879e-21, 5.61541e-20, 
    3.059099e-20, 4.22108e-20, -1.695172e-20, 1.82915e-20, -7.109433e-20, 
    1.158868e-20, -6.064935e-20, 5.66068e-20, -1.812884e-20, -4.377217e-21, 
    -3.013369e-20, 1.638766e-20, -8.849536e-21, 2.986745e-21, -7.517207e-21, 
    1.835956e-20, -1.474935e-20, 2.99211e-21, 8.249317e-20, -6.120689e-20, 
    -7.533984e-20, -4.564115e-20, -3.096286e-20, 1.416125e-20, 9.985265e-21, 
    -2.757441e-21, 4.945248e-21, -4.332511e-20, -4.89707e-20, -2.974236e-20, 
    -3.397118e-20, 1.846426e-21, 2.868701e-20, 8.28873e-20, 6.397629e-21, 
    9.377487e-22, -1.425182e-21, -6.558464e-20, -1.717759e-20, 2.005233e-20, 
    2.399132e-20, -1.56084e-20, 9.083962e-20, -3.250207e-20, -1.38633e-20, 
    1.111775e-20, 1.389309e-21, -3.8568e-20, 2.001616e-20, 3.138819e-21, 
    -2.398639e-20, -3.183206e-20, -5.059036e-20, -3.114727e-21, 4.586286e-20, 
    -3.035182e-20, 8.644366e-20, 4.016519e-20, -1.892729e-20, 1.141729e-20, 
    -1.482125e-20, -5.032271e-20, -6.959532e-23, 5.639702e-20, 8.248853e-21, 
    1.167437e-20, -1.762498e-20, 3.214592e-20, 1.762543e-20, -5.992074e-20, 
    8.421782e-21, 2.127394e-21, 4.13221e-20, -4.310748e-20, -7.461423e-21, 
    1.188337e-20, -2.115255e-20, -7.743329e-20, 4.635999e-20, 2.76523e-20, 
    -2.592629e-20, 2.817687e-20, -6.387813e-20, 3.344197e-20, 2.189698e-20, 
    -2.06842e-21, -7.41293e-21, -1.087593e-19, 6.879248e-21, 4.550485e-20, 
    1.459818e-20, -5.30042e-20, 1.845436e-20, -1.631172e-20, -3.939492e-20, 
    -7.499873e-20, 1.463317e-20, 4.167118e-20, 5.453739e-20, 5.502157e-21, 
    3.450963e-20, 3.583629e-20, 2.004864e-21, 3.640138e-20, -5.200511e-20, 
    7.96408e-21, -4.043587e-20, -1.621425e-20, -2.959982e-20, 3.444836e-20, 
    1.069272e-20, 7.942012e-20, 7.111012e-20, 3.403563e-20, 2.335646e-20, 
    9.168804e-21, -7.670029e-21, 1.009991e-20, 2.006832e-20, 1.777887e-20, 
    -4.07633e-21, 3.393858e-20, -1.827358e-20, 3.772533e-20, 2.498536e-20, 
    8.175131e-20, -4.007458e-20, 8.040823e-20, -2.283666e-20, -1.444605e-20, 
    -7.684224e-20, -2.848146e-20, 9.348851e-21, -2.884586e-20, 2.776217e-20, 
    -2.782957e-20, -1.944125e-20, -9.448025e-21, -3.898638e-20, 
    -4.547635e-21, -2.373381e-20, 3.323341e-20, 3.440055e-20, -2.857653e-20, 
    5.61646e-21, 9.772121e-21, -1.916269e-20, 5.186e-21, -7.205079e-23, 
    -4.204013e-21, -2.233145e-20, -4.554e-20, -2.206438e-20, 3.499556e-20, 
    1.239575e-20, -2.470792e-20, -1.829226e-20, -3.48238e-21, -2.666211e-20, 
    -1.52781e-20, -2.857212e-20, -7.351045e-21, 3.485153e-22, 2.282711e-21, 
    -7.780807e-20, 1.989674e-20, 5.101242e-20, 3.557692e-20, 1.436729e-21, 
    -7.367761e-21, -2.538598e-20, -2.077053e-20, -2.685027e-20, 2.957197e-20, 
    4.368627e-20, 7.406494e-20, 2.29796e-20, 2.115373e-20, 1.401451e-20, 
    -2.884041e-20, 2.909515e-20, -1.998245e-21, 2.899389e-20, 2.14882e-20, 
    4.33754e-21, 4.239214e-20, 9.754966e-20, -3.653635e-20, -8.048204e-20, 
    -2.882958e-20, -2.967465e-20, 2.40871e-20, 7.646506e-20, 3.410087e-20, 
    4.988607e-20, -1.407674e-20, 2.473295e-20, -4.326298e-20, 5.004951e-20, 
    2.228475e-20, 8.148906e-21, 2.283374e-20, -2.496867e-20, -1.735347e-21, 
    -1.190973e-20, 5.050898e-20, 3.509064e-20, 7.430893e-22, 6.069374e-20, 
    2.460226e-21, 2.227606e-20, 4.957216e-20, 2.815242e-20, -4.827562e-20, 
    5.219333e-20, -1.161311e-20, 1.832984e-21, 3.945207e-20, 1.865998e-20, 
    3.64541e-20, -1.184974e-20, -1.810585e-21, -3.810753e-20, 6.348742e-20, 
    -1.652272e-20, -2.925065e-20, -5.724356e-20, -3.476509e-20, 4.921742e-20, 
    6.587955e-20, 2.494048e-20, -4.218126e-21, -1.845564e-20, -1.142723e-20, 
    -1.757401e-20, 1.608307e-20, -4.321702e-20, -2.208232e-20, -1.784726e-20, 
    -2.343215e-20, -2.060463e-20, 5.742045e-20, 5.736216e-21, 4.02224e-20, 
    -3.036512e-20, -2.053614e-20, -4.625486e-20, 2.311636e-20, -3.46999e-20, 
    2.419441e-20, 4.31964e-20, 3.11294e-20, -1.072736e-20, -2.998775e-20, 
    5.556651e-20, 8.888771e-21, 2.861457e-20, -3.073492e-20, -3.679506e-20, 
    5.037674e-20, -8.113181e-20, 6.28956e-20, 8.477449e-20, -3.307498e-20, 
    2.516808e-20, 1.926103e-20, -2.817033e-21, 4.152434e-20, 1.392474e-20, 
    2.791535e-20, -3.322734e-20, -5.263906e-20, 2.78325e-20, -2.30044e-20, 
    -5.119578e-21, -3.744333e-20, -1.936367e-20, 2.077072e-20, -5.849072e-21, 
    5.129816e-20, -1.535525e-20, -1.097237e-20, 1.841254e-20, -2.713964e-20, 
    3.162929e-20, -1.680854e-20, -1.605227e-20, 1.841599e-20, -7.504367e-20, 
    1.685996e-20, -1.996504e-20, -4.700038e-20, -6.696237e-20, -6.770071e-21, 
    3.088982e-20, 4.585941e-20, 5.066639e-20, 2.168741e-20, -1.123256e-20, 
    -3.693876e-21, 2.679999e-21, 6.245959e-20, -1.794455e-21, 4.824228e-20, 
    3.351146e-20, 5.133601e-20, -3.846757e-20, 3.225811e-20, 1.384046e-20, 
    1.200112e-20, -4.529867e-20, 1.169699e-20, 1.595541e-20, -6.536584e-21, 
    4.252089e-20, -1.519833e-20, -3.945135e-20, -4.844152e-20, 1.59701e-20, 
    8.19501e-20, -4.733438e-20, 1.036044e-19, 3.475347e-20, 2.097446e-20, 
    9.633883e-21, -6.30339e-20, 8.493184e-21, -3.675565e-20 ;

 SR =
  6.191209e-08, 6.218511e-08, 6.213204e-08, 6.235225e-08, 6.22301e-08, 
    6.237429e-08, 6.196745e-08, 6.219594e-08, 6.205008e-08, 6.193667e-08, 
    6.277961e-08, 6.236208e-08, 6.321343e-08, 6.29471e-08, 6.361618e-08, 
    6.317198e-08, 6.370576e-08, 6.360339e-08, 6.391155e-08, 6.382326e-08, 
    6.421742e-08, 6.39523e-08, 6.442178e-08, 6.415411e-08, 6.419598e-08, 
    6.394355e-08, 6.244612e-08, 6.272763e-08, 6.242944e-08, 6.246958e-08, 
    6.245157e-08, 6.223262e-08, 6.212228e-08, 6.189123e-08, 6.193318e-08, 
    6.210288e-08, 6.248763e-08, 6.235703e-08, 6.26862e-08, 6.267877e-08, 
    6.304526e-08, 6.288002e-08, 6.349605e-08, 6.332096e-08, 6.382695e-08, 
    6.369969e-08, 6.382097e-08, 6.37842e-08, 6.382145e-08, 6.363481e-08, 
    6.371478e-08, 6.355055e-08, 6.291096e-08, 6.309892e-08, 6.253835e-08, 
    6.220129e-08, 6.197747e-08, 6.181863e-08, 6.184109e-08, 6.188389e-08, 
    6.210387e-08, 6.231072e-08, 6.246836e-08, 6.25738e-08, 6.267771e-08, 
    6.299219e-08, 6.315867e-08, 6.353144e-08, 6.346419e-08, 6.357814e-08, 
    6.368703e-08, 6.386984e-08, 6.383975e-08, 6.392029e-08, 6.357515e-08, 
    6.380452e-08, 6.342587e-08, 6.352943e-08, 6.27059e-08, 6.239227e-08, 
    6.225892e-08, 6.214224e-08, 6.185834e-08, 6.205439e-08, 6.19771e-08, 
    6.216099e-08, 6.227782e-08, 6.222004e-08, 6.257669e-08, 6.243803e-08, 
    6.316854e-08, 6.285387e-08, 6.367434e-08, 6.347799e-08, 6.372139e-08, 
    6.359719e-08, 6.381001e-08, 6.361848e-08, 6.395027e-08, 6.402251e-08, 
    6.397314e-08, 6.41628e-08, 6.360786e-08, 6.382096e-08, 6.221842e-08, 
    6.222784e-08, 6.227175e-08, 6.207874e-08, 6.206693e-08, 6.189008e-08, 
    6.204745e-08, 6.211446e-08, 6.22846e-08, 6.238523e-08, 6.248089e-08, 
    6.269123e-08, 6.292615e-08, 6.325467e-08, 6.349072e-08, 6.364895e-08, 
    6.355192e-08, 6.363758e-08, 6.354183e-08, 6.349695e-08, 6.399544e-08, 
    6.371552e-08, 6.413553e-08, 6.411229e-08, 6.39222e-08, 6.411491e-08, 
    6.223446e-08, 6.218023e-08, 6.199193e-08, 6.213929e-08, 6.187082e-08, 
    6.202109e-08, 6.210749e-08, 6.244091e-08, 6.251418e-08, 6.258211e-08, 
    6.271628e-08, 6.288847e-08, 6.319055e-08, 6.34534e-08, 6.369337e-08, 
    6.367579e-08, 6.368198e-08, 6.373558e-08, 6.36028e-08, 6.375738e-08, 
    6.378333e-08, 6.371549e-08, 6.410917e-08, 6.39967e-08, 6.411179e-08, 
    6.403856e-08, 6.219786e-08, 6.228911e-08, 6.22398e-08, 6.233252e-08, 
    6.22672e-08, 6.255767e-08, 6.264477e-08, 6.305234e-08, 6.288508e-08, 
    6.315129e-08, 6.291213e-08, 6.29545e-08, 6.315996e-08, 6.292505e-08, 
    6.34389e-08, 6.30905e-08, 6.373767e-08, 6.338972e-08, 6.375947e-08, 
    6.369233e-08, 6.38035e-08, 6.390305e-08, 6.402831e-08, 6.425942e-08, 
    6.420591e-08, 6.43992e-08, 6.242516e-08, 6.254352e-08, 6.25331e-08, 
    6.265698e-08, 6.27486e-08, 6.294718e-08, 6.326568e-08, 6.314591e-08, 
    6.33658e-08, 6.340995e-08, 6.307588e-08, 6.328098e-08, 6.262274e-08, 
    6.272907e-08, 6.266577e-08, 6.243449e-08, 6.317349e-08, 6.279422e-08, 
    6.349462e-08, 6.328914e-08, 6.388886e-08, 6.359058e-08, 6.417645e-08, 
    6.442689e-08, 6.466265e-08, 6.493813e-08, 6.260812e-08, 6.25277e-08, 
    6.267172e-08, 6.287096e-08, 6.305586e-08, 6.330166e-08, 6.332682e-08, 
    6.337287e-08, 6.349217e-08, 6.359246e-08, 6.338743e-08, 6.361761e-08, 
    6.275372e-08, 6.320642e-08, 6.249729e-08, 6.27108e-08, 6.285921e-08, 
    6.279412e-08, 6.313223e-08, 6.321191e-08, 6.353574e-08, 6.336835e-08, 
    6.436507e-08, 6.392407e-08, 6.514793e-08, 6.480587e-08, 6.249959e-08, 
    6.260785e-08, 6.298463e-08, 6.280536e-08, 6.331808e-08, 6.344429e-08, 
    6.35469e-08, 6.367805e-08, 6.369222e-08, 6.376993e-08, 6.364259e-08, 
    6.376491e-08, 6.330219e-08, 6.350896e-08, 6.294157e-08, 6.307966e-08, 
    6.301614e-08, 6.294646e-08, 6.316152e-08, 6.339064e-08, 6.339556e-08, 
    6.346902e-08, 6.367603e-08, 6.332016e-08, 6.442196e-08, 6.374147e-08, 
    6.27259e-08, 6.293441e-08, 6.296421e-08, 6.288344e-08, 6.343164e-08, 
    6.3233e-08, 6.376804e-08, 6.362344e-08, 6.386038e-08, 6.374263e-08, 
    6.372531e-08, 6.357409e-08, 6.347994e-08, 6.32421e-08, 6.304859e-08, 
    6.289515e-08, 6.293084e-08, 6.309938e-08, 6.340467e-08, 6.36935e-08, 
    6.363022e-08, 6.384236e-08, 6.32809e-08, 6.351632e-08, 6.342533e-08, 
    6.36626e-08, 6.314273e-08, 6.358538e-08, 6.302958e-08, 6.307831e-08, 
    6.322905e-08, 6.353228e-08, 6.359939e-08, 6.367102e-08, 6.362682e-08, 
    6.341242e-08, 6.33773e-08, 6.322539e-08, 6.318344e-08, 6.30677e-08, 
    6.297188e-08, 6.305942e-08, 6.315137e-08, 6.341251e-08, 6.364786e-08, 
    6.390447e-08, 6.396727e-08, 6.426707e-08, 6.4023e-08, 6.442575e-08, 
    6.40833e-08, 6.467612e-08, 6.361105e-08, 6.407326e-08, 6.323592e-08, 
    6.332613e-08, 6.348927e-08, 6.386351e-08, 6.366148e-08, 6.389776e-08, 
    6.337593e-08, 6.310519e-08, 6.303516e-08, 6.290448e-08, 6.303815e-08, 
    6.302728e-08, 6.315518e-08, 6.311409e-08, 6.342119e-08, 6.325622e-08, 
    6.372487e-08, 6.38959e-08, 6.437893e-08, 6.467506e-08, 6.497654e-08, 
    6.510964e-08, 6.515015e-08, 6.516709e-08 ;

 STORVEGC =
  0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 0.7217545, 
    0.7217545, 0.7217545 ;

 STORVEGN =
  0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 0.02887061, 
    0.02887061, 0.02887061 ;

 SUPPLEMENT_TO_SMINN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 SoilAlpha =
  0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999958, 0.9999957, 0.9999958, 0.9999958, 
    0.9999958, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999958, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999958, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999958, 
    0.9999958, 0.9999958, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999958, 0.9999958, 0.9999958, 0.9999958, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999958, 0.9999957, 0.9999958, 0.9999958, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999958, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999958, 0.9999957, 0.9999958, 0.9999957, 0.9999958, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 0.9999957, 
    0.9999957, 0.9999957, 0.9999958, 0.9999958, 0.9999958, 0.9999958, 
    0.9999958, 0.9999958 ;

 SoilAlpha_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TAUX =
  -0.3396222, -0.339627, -0.3396261, -0.3396298, -0.3396278, -0.3396302, 
    -0.3396232, -0.3396271, -0.3396247, -0.3396227, -0.3396372, -0.33963, 
    -0.3396453, -0.3396405, -0.3396526, -0.3396445, -0.3396542, -0.3396524, 
    -0.3396581, -0.3396565, -0.3396635, -0.3396588, -0.3396673, -0.3396624, 
    -0.3396631, -0.3396586, -0.3396315, -0.3396363, -0.3396312, -0.3396319, 
    -0.3396316, -0.3396278, -0.3396258, -0.3396219, -0.3396226, -0.3396255, 
    -0.3396322, -0.33963, -0.3396358, -0.3396357, -0.3396423, -0.3396393, 
    -0.3396505, -0.3396473, -0.3396565, -0.3396542, -0.3396564, -0.3396558, 
    -0.3396564, -0.339653, -0.3396544, -0.3396515, -0.3396399, -0.3396432, 
    -0.3396331, -0.3396271, -0.3396234, -0.3396207, -0.3396211, -0.3396218, 
    -0.3396255, -0.3396292, -0.3396319, -0.3396338, -0.3396357, -0.3396412, 
    -0.3396443, -0.3396511, -0.3396499, -0.3396519, -0.339654, -0.3396573, 
    -0.3396567, -0.3396582, -0.3396519, -0.3396561, -0.3396493, -0.3396511, 
    -0.3396359, -0.3396306, -0.3396281, -0.3396262, -0.3396213, -0.3396247, 
    -0.3396234, -0.3396266, -0.3396286, -0.3396276, -0.3396339, -0.3396314, 
    -0.3396445, -0.3396388, -0.3396537, -0.3396502, -0.3396546, -0.3396524, 
    -0.3396562, -0.3396527, -0.3396588, -0.33966, -0.3396592, -0.3396626, 
    -0.3396525, -0.3396564, -0.3396276, -0.3396277, -0.3396285, -0.3396251, 
    -0.3396249, -0.3396219, -0.3396246, -0.3396257, -0.3396288, -0.3396305, 
    -0.3396322, -0.3396359, -0.3396401, -0.3396461, -0.3396504, -0.3396533, 
    -0.3396515, -0.3396531, -0.3396513, -0.3396505, -0.3396595, -0.3396544, 
    -0.3396621, -0.3396617, -0.3396582, -0.3396618, -0.3396279, -0.3396269, 
    -0.3396237, -0.3396262, -0.3396216, -0.3396241, -0.3396256, -0.3396314, 
    -0.3396327, -0.3396339, -0.3396364, -0.3396395, -0.3396449, -0.3396497, 
    -0.3396541, -0.3396538, -0.3396539, -0.3396549, -0.3396524, -0.3396553, 
    -0.3396557, -0.3396545, -0.3396617, -0.3396596, -0.3396617, -0.3396604, 
    -0.3396272, -0.3396288, -0.339628, -0.3396295, -0.3396284, -0.3396334, 
    -0.339635, -0.3396423, -0.3396394, -0.3396442, -0.3396399, -0.3396406, 
    -0.3396442, -0.3396402, -0.3396493, -0.339643, -0.3396549, -0.3396484, 
    -0.3396553, -0.3396541, -0.3396561, -0.3396579, -0.3396602, -0.3396643, 
    -0.3396634, -0.3396669, -0.3396312, -0.3396332, -0.3396331, -0.3396353, 
    -0.339637, -0.3396406, -0.3396463, -0.3396442, -0.3396482, -0.3396489, 
    -0.3396429, -0.3396465, -0.3396347, -0.3396365, -0.3396354, -0.3396313, 
    -0.3396446, -0.3396377, -0.3396505, -0.3396467, -0.3396576, -0.3396522, 
    -0.3396628, -0.3396673, -0.3396717, -0.3396766, -0.3396344, -0.339633, 
    -0.3396356, -0.3396391, -0.3396425, -0.339647, -0.3396474, -0.3396482, 
    -0.3396505, -0.3396523, -0.3396485, -0.3396527, -0.3396368, -0.3396452, 
    -0.3396324, -0.3396361, -0.3396389, -0.3396378, -0.3396439, -0.3396454, 
    -0.3396512, -0.3396482, -0.3396661, -0.3396582, -0.3396806, -0.3396742, 
    -0.3396325, -0.3396344, -0.3396412, -0.339638, -0.3396473, -0.3396496, 
    -0.3396514, -0.3396538, -0.3396541, -0.3396555, -0.3396532, -0.3396554, 
    -0.339647, -0.3396508, -0.3396405, -0.3396429, -0.3396418, -0.3396406, 
    -0.3396445, -0.3396485, -0.3396487, -0.33965, -0.3396534, -0.3396473, 
    -0.339667, -0.3396547, -0.3396366, -0.3396402, -0.3396409, -0.3396394, 
    -0.3396493, -0.3396457, -0.3396554, -0.3396528, -0.3396571, -0.339655, 
    -0.3396547, -0.3396519, -0.3396502, -0.3396459, -0.3396423, -0.3396396, 
    -0.3396403, -0.3396433, -0.3396488, -0.3396541, -0.3396529, -0.3396568, 
    -0.3396466, -0.3396508, -0.3396492, -0.3396535, -0.3396441, -0.3396518, 
    -0.3396421, -0.3396429, -0.3396457, -0.339651, -0.3396524, -0.3396536, 
    -0.3396529, -0.3396489, -0.3396483, -0.3396456, -0.3396448, -0.3396428, 
    -0.339641, -0.3396426, -0.3396442, -0.339649, -0.3396532, -0.3396579, 
    -0.3396591, -0.3396643, -0.3396599, -0.339667, -0.3396608, -0.3396717, 
    -0.3396524, -0.3396608, -0.3396458, -0.3396474, -0.3396503, -0.3396571, 
    -0.3396535, -0.3396577, -0.3396483, -0.3396433, -0.3396422, -0.3396398, 
    -0.3396422, -0.339642, -0.3396443, -0.3396436, -0.3396491, -0.3396462, 
    -0.3396546, -0.3396577, -0.3396665, -0.3396719, -0.3396775, -0.3396799, 
    -0.3396807, -0.339681 ;

 TAUY =
  -0.3396222, -0.339627, -0.3396261, -0.3396298, -0.3396278, -0.3396302, 
    -0.3396232, -0.3396271, -0.3396247, -0.3396227, -0.3396372, -0.33963, 
    -0.3396453, -0.3396405, -0.3396526, -0.3396445, -0.3396542, -0.3396524, 
    -0.3396581, -0.3396565, -0.3396635, -0.3396588, -0.3396673, -0.3396624, 
    -0.3396631, -0.3396586, -0.3396315, -0.3396363, -0.3396312, -0.3396319, 
    -0.3396316, -0.3396278, -0.3396258, -0.3396219, -0.3396226, -0.3396255, 
    -0.3396322, -0.33963, -0.3396358, -0.3396357, -0.3396423, -0.3396393, 
    -0.3396505, -0.3396473, -0.3396565, -0.3396542, -0.3396564, -0.3396558, 
    -0.3396564, -0.339653, -0.3396544, -0.3396515, -0.3396399, -0.3396432, 
    -0.3396331, -0.3396271, -0.3396234, -0.3396207, -0.3396211, -0.3396218, 
    -0.3396255, -0.3396292, -0.3396319, -0.3396338, -0.3396357, -0.3396412, 
    -0.3396443, -0.3396511, -0.3396499, -0.3396519, -0.339654, -0.3396573, 
    -0.3396567, -0.3396582, -0.3396519, -0.3396561, -0.3396493, -0.3396511, 
    -0.3396359, -0.3396306, -0.3396281, -0.3396262, -0.3396213, -0.3396247, 
    -0.3396234, -0.3396266, -0.3396286, -0.3396276, -0.3396339, -0.3396314, 
    -0.3396445, -0.3396388, -0.3396537, -0.3396502, -0.3396546, -0.3396524, 
    -0.3396562, -0.3396527, -0.3396588, -0.33966, -0.3396592, -0.3396626, 
    -0.3396525, -0.3396564, -0.3396276, -0.3396277, -0.3396285, -0.3396251, 
    -0.3396249, -0.3396219, -0.3396246, -0.3396257, -0.3396288, -0.3396305, 
    -0.3396322, -0.3396359, -0.3396401, -0.3396461, -0.3396504, -0.3396533, 
    -0.3396515, -0.3396531, -0.3396513, -0.3396505, -0.3396595, -0.3396544, 
    -0.3396621, -0.3396617, -0.3396582, -0.3396618, -0.3396279, -0.3396269, 
    -0.3396237, -0.3396262, -0.3396216, -0.3396241, -0.3396256, -0.3396314, 
    -0.3396327, -0.3396339, -0.3396364, -0.3396395, -0.3396449, -0.3396497, 
    -0.3396541, -0.3396538, -0.3396539, -0.3396549, -0.3396524, -0.3396553, 
    -0.3396557, -0.3396545, -0.3396617, -0.3396596, -0.3396617, -0.3396604, 
    -0.3396272, -0.3396288, -0.339628, -0.3396295, -0.3396284, -0.3396334, 
    -0.339635, -0.3396423, -0.3396394, -0.3396442, -0.3396399, -0.3396406, 
    -0.3396442, -0.3396402, -0.3396493, -0.339643, -0.3396549, -0.3396484, 
    -0.3396553, -0.3396541, -0.3396561, -0.3396579, -0.3396602, -0.3396643, 
    -0.3396634, -0.3396669, -0.3396312, -0.3396332, -0.3396331, -0.3396353, 
    -0.339637, -0.3396406, -0.3396463, -0.3396442, -0.3396482, -0.3396489, 
    -0.3396429, -0.3396465, -0.3396347, -0.3396365, -0.3396354, -0.3396313, 
    -0.3396446, -0.3396377, -0.3396505, -0.3396467, -0.3396576, -0.3396522, 
    -0.3396628, -0.3396673, -0.3396717, -0.3396766, -0.3396344, -0.339633, 
    -0.3396356, -0.3396391, -0.3396425, -0.339647, -0.3396474, -0.3396482, 
    -0.3396505, -0.3396523, -0.3396485, -0.3396527, -0.3396368, -0.3396452, 
    -0.3396324, -0.3396361, -0.3396389, -0.3396378, -0.3396439, -0.3396454, 
    -0.3396512, -0.3396482, -0.3396661, -0.3396582, -0.3396806, -0.3396742, 
    -0.3396325, -0.3396344, -0.3396412, -0.339638, -0.3396473, -0.3396496, 
    -0.3396514, -0.3396538, -0.3396541, -0.3396555, -0.3396532, -0.3396554, 
    -0.339647, -0.3396508, -0.3396405, -0.3396429, -0.3396418, -0.3396406, 
    -0.3396445, -0.3396485, -0.3396487, -0.33965, -0.3396534, -0.3396473, 
    -0.339667, -0.3396547, -0.3396366, -0.3396402, -0.3396409, -0.3396394, 
    -0.3396493, -0.3396457, -0.3396554, -0.3396528, -0.3396571, -0.339655, 
    -0.3396547, -0.3396519, -0.3396502, -0.3396459, -0.3396423, -0.3396396, 
    -0.3396403, -0.3396433, -0.3396488, -0.3396541, -0.3396529, -0.3396568, 
    -0.3396466, -0.3396508, -0.3396492, -0.3396535, -0.3396441, -0.3396518, 
    -0.3396421, -0.3396429, -0.3396457, -0.339651, -0.3396524, -0.3396536, 
    -0.3396529, -0.3396489, -0.3396483, -0.3396456, -0.3396448, -0.3396428, 
    -0.339641, -0.3396426, -0.3396442, -0.339649, -0.3396532, -0.3396579, 
    -0.3396591, -0.3396643, -0.3396599, -0.339667, -0.3396608, -0.3396717, 
    -0.3396524, -0.3396608, -0.3396458, -0.3396474, -0.3396503, -0.3396571, 
    -0.3396535, -0.3396577, -0.3396483, -0.3396433, -0.3396422, -0.3396398, 
    -0.3396422, -0.339642, -0.3396443, -0.3396436, -0.3396491, -0.3396462, 
    -0.3396546, -0.3396577, -0.3396665, -0.3396719, -0.3396775, -0.3396799, 
    -0.3396807, -0.339681 ;

 TBOT =
  253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605 ;

 TBUILD =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TG =
  261.0567, 261.0778, 261.0737, 261.0907, 261.0813, 261.0924, 261.061, 
    261.0786, 261.0674, 261.0586, 261.1237, 261.0915, 261.1573, 261.1367, 
    261.1883, 261.154, 261.1953, 261.1874, 261.2112, 261.2043, 261.2347, 
    261.2143, 261.2505, 261.2299, 261.2331, 261.2136, 261.098, 261.1197, 
    261.0967, 261.0998, 261.0984, 261.0815, 261.073, 261.0551, 261.0584, 
    261.0715, 261.1012, 261.0911, 261.1165, 261.116, 261.1443, 261.1315, 
    261.1791, 261.1656, 261.2046, 261.1948, 261.2042, 261.2013, 261.2042, 
    261.1898, 261.196, 261.1833, 261.1339, 261.1484, 261.1051, 261.079, 
    261.0618, 261.0495, 261.0512, 261.0546, 261.0715, 261.0875, 261.0997, 
    261.1078, 261.1159, 261.1401, 261.153, 261.1818, 261.1766, 261.1854, 
    261.1938, 261.2079, 261.2056, 261.2118, 261.1852, 261.2029, 261.1737, 
    261.1817, 261.118, 261.0938, 261.0835, 261.0745, 261.0526, 261.0677, 
    261.0618, 261.076, 261.085, 261.0805, 261.1081, 261.0974, 261.1538, 
    261.1295, 261.1928, 261.1777, 261.1965, 261.1869, 261.2033, 261.1885, 
    261.2141, 261.2197, 261.2159, 261.2305, 261.1877, 261.2042, 261.0804, 
    261.0811, 261.0845, 261.0696, 261.0687, 261.055, 261.0672, 261.0724, 
    261.0855, 261.0933, 261.1007, 261.1169, 261.1351, 261.1604, 261.1787, 
    261.1909, 261.1834, 261.19, 261.1826, 261.1792, 261.2176, 261.196, 
    261.2284, 261.2267, 261.212, 261.2268, 261.0816, 261.0775, 261.0629, 
    261.0743, 261.0536, 261.0652, 261.0718, 261.0976, 261.1033, 261.1085, 
    261.1189, 261.1322, 261.1555, 261.1758, 261.1943, 261.193, 261.1935, 
    261.1976, 261.1873, 261.1992, 261.2013, 261.196, 261.2264, 261.2177, 
    261.2266, 261.2209, 261.0788, 261.0859, 261.0821, 261.0892, 261.0842, 
    261.1066, 261.1133, 261.1448, 261.1319, 261.1525, 261.134, 261.1373, 
    261.1531, 261.135, 261.1747, 261.1477, 261.1977, 261.1708, 261.1994, 
    261.1942, 261.2028, 261.2105, 261.2202, 261.238, 261.2339, 261.2488, 
    261.0964, 261.1055, 261.1047, 261.1143, 261.1214, 261.1367, 261.1613, 
    261.152, 261.169, 261.1724, 261.1466, 261.1625, 261.1116, 261.1198, 
    261.115, 261.0971, 261.1542, 261.1249, 261.179, 261.1631, 261.2094, 
    261.1864, 261.2316, 261.2509, 261.2691, 261.2903, 261.1105, 261.1043, 
    261.1154, 261.1308, 261.1451, 261.1641, 261.166, 261.1696, 261.1788, 
    261.1865, 261.1707, 261.1885, 261.1217, 261.1567, 261.102, 261.1184, 
    261.1299, 261.1249, 261.151, 261.1571, 261.1821, 261.1692, 261.2461, 
    261.2121, 261.3065, 261.2801, 261.1021, 261.1105, 261.1396, 261.1257, 
    261.1653, 261.1751, 261.183, 261.1931, 261.1942, 261.2002, 261.1904, 
    261.1998, 261.1641, 261.1801, 261.1363, 261.1469, 261.142, 261.1367, 
    261.1533, 261.1709, 261.1713, 261.177, 261.1929, 261.1655, 261.2505, 
    261.198, 261.1196, 261.1357, 261.138, 261.1318, 261.1741, 261.1588, 
    261.2001, 261.1889, 261.2072, 261.1981, 261.1968, 261.1851, 261.1778, 
    261.1595, 261.1445, 261.1327, 261.1354, 261.1484, 261.172, 261.1943, 
    261.1894, 261.2058, 261.1625, 261.1806, 261.1736, 261.1919, 261.1518, 
    261.1859, 261.1431, 261.1468, 261.1585, 261.1819, 261.1871, 261.1926, 
    261.1892, 261.1726, 261.1699, 261.1582, 261.1549, 261.146, 261.1386, 
    261.1454, 261.1525, 261.1726, 261.1908, 261.2106, 261.2155, 261.2386, 
    261.2197, 261.2508, 261.2243, 261.2701, 261.1879, 261.2236, 261.159, 
    261.166, 261.1786, 261.2074, 261.1919, 261.2101, 261.1698, 261.1489, 
    261.1435, 261.1334, 261.1437, 261.1429, 261.1528, 261.1496, 261.1733, 
    261.1606, 261.1967, 261.2099, 261.2472, 261.27, 261.2933, 261.3036, 
    261.3067, 261.308 ;

 TG_R =
  261.0567, 261.0778, 261.0737, 261.0907, 261.0813, 261.0924, 261.061, 
    261.0786, 261.0674, 261.0586, 261.1237, 261.0915, 261.1573, 261.1367, 
    261.1883, 261.154, 261.1953, 261.1874, 261.2112, 261.2043, 261.2347, 
    261.2143, 261.2505, 261.2299, 261.2331, 261.2136, 261.098, 261.1197, 
    261.0967, 261.0998, 261.0984, 261.0815, 261.073, 261.0551, 261.0584, 
    261.0715, 261.1012, 261.0911, 261.1165, 261.116, 261.1443, 261.1315, 
    261.1791, 261.1656, 261.2046, 261.1948, 261.2042, 261.2013, 261.2042, 
    261.1898, 261.196, 261.1833, 261.1339, 261.1484, 261.1051, 261.079, 
    261.0618, 261.0495, 261.0512, 261.0546, 261.0715, 261.0875, 261.0997, 
    261.1078, 261.1159, 261.1401, 261.153, 261.1818, 261.1766, 261.1854, 
    261.1938, 261.2079, 261.2056, 261.2118, 261.1852, 261.2029, 261.1737, 
    261.1817, 261.118, 261.0938, 261.0835, 261.0745, 261.0526, 261.0677, 
    261.0618, 261.076, 261.085, 261.0805, 261.1081, 261.0974, 261.1538, 
    261.1295, 261.1928, 261.1777, 261.1965, 261.1869, 261.2033, 261.1885, 
    261.2141, 261.2197, 261.2159, 261.2305, 261.1877, 261.2042, 261.0804, 
    261.0811, 261.0845, 261.0696, 261.0687, 261.055, 261.0672, 261.0724, 
    261.0855, 261.0933, 261.1007, 261.1169, 261.1351, 261.1604, 261.1787, 
    261.1909, 261.1834, 261.19, 261.1826, 261.1792, 261.2176, 261.196, 
    261.2284, 261.2267, 261.212, 261.2268, 261.0816, 261.0775, 261.0629, 
    261.0743, 261.0536, 261.0652, 261.0718, 261.0976, 261.1033, 261.1085, 
    261.1189, 261.1322, 261.1555, 261.1758, 261.1943, 261.193, 261.1935, 
    261.1976, 261.1873, 261.1992, 261.2013, 261.196, 261.2264, 261.2177, 
    261.2266, 261.2209, 261.0788, 261.0859, 261.0821, 261.0892, 261.0842, 
    261.1066, 261.1133, 261.1448, 261.1319, 261.1525, 261.134, 261.1373, 
    261.1531, 261.135, 261.1747, 261.1477, 261.1977, 261.1708, 261.1994, 
    261.1942, 261.2028, 261.2105, 261.2202, 261.238, 261.2339, 261.2488, 
    261.0964, 261.1055, 261.1047, 261.1143, 261.1214, 261.1367, 261.1613, 
    261.152, 261.169, 261.1724, 261.1466, 261.1625, 261.1116, 261.1198, 
    261.115, 261.0971, 261.1542, 261.1249, 261.179, 261.1631, 261.2094, 
    261.1864, 261.2316, 261.2509, 261.2691, 261.2903, 261.1105, 261.1043, 
    261.1154, 261.1308, 261.1451, 261.1641, 261.166, 261.1696, 261.1788, 
    261.1865, 261.1707, 261.1885, 261.1217, 261.1567, 261.102, 261.1184, 
    261.1299, 261.1249, 261.151, 261.1571, 261.1821, 261.1692, 261.2461, 
    261.2121, 261.3065, 261.2801, 261.1021, 261.1105, 261.1396, 261.1257, 
    261.1653, 261.1751, 261.183, 261.1931, 261.1942, 261.2002, 261.1904, 
    261.1998, 261.1641, 261.1801, 261.1363, 261.1469, 261.142, 261.1367, 
    261.1533, 261.1709, 261.1713, 261.177, 261.1929, 261.1655, 261.2505, 
    261.198, 261.1196, 261.1357, 261.138, 261.1318, 261.1741, 261.1588, 
    261.2001, 261.1889, 261.2072, 261.1981, 261.1968, 261.1851, 261.1778, 
    261.1595, 261.1445, 261.1327, 261.1354, 261.1484, 261.172, 261.1943, 
    261.1894, 261.2058, 261.1625, 261.1806, 261.1736, 261.1919, 261.1518, 
    261.1859, 261.1431, 261.1468, 261.1585, 261.1819, 261.1871, 261.1926, 
    261.1892, 261.1726, 261.1699, 261.1582, 261.1549, 261.146, 261.1386, 
    261.1454, 261.1525, 261.1726, 261.1908, 261.2106, 261.2155, 261.2386, 
    261.2197, 261.2508, 261.2243, 261.2701, 261.1879, 261.2236, 261.159, 
    261.166, 261.1786, 261.2074, 261.1919, 261.2101, 261.1698, 261.1489, 
    261.1435, 261.1334, 261.1437, 261.1429, 261.1528, 261.1496, 261.1733, 
    261.1606, 261.1967, 261.2099, 261.2472, 261.27, 261.2933, 261.3036, 
    261.3067, 261.308 ;

 TG_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TH2OSFC =
  254.483, 254.4845, 254.4842, 254.4854, 254.4848, 254.4855, 254.4833, 
    254.4846, 254.4838, 254.4832, 254.4877, 254.4855, 254.4901, 254.4887, 
    254.4923, 254.4899, 254.4928, 254.4923, 254.494, 254.4935, 254.4956, 
    254.4942, 254.4968, 254.4953, 254.4955, 254.4942, 254.4859, 254.4874, 
    254.4858, 254.4861, 254.486, 254.4848, 254.4841, 254.4829, 254.4831, 
    254.4841, 254.4861, 254.4854, 254.4872, 254.4872, 254.4892, 254.4883, 
    254.4917, 254.4907, 254.4935, 254.4928, 254.4935, 254.4933, 254.4935, 
    254.4924, 254.4929, 254.492, 254.4885, 254.4895, 254.4864, 254.4846, 
    254.4834, 254.4825, 254.4826, 254.4829, 254.4841, 254.4852, 254.4861, 
    254.4866, 254.4872, 254.4889, 254.4898, 254.4919, 254.4915, 254.4921, 
    254.4927, 254.4937, 254.4936, 254.494, 254.4921, 254.4934, 254.4913, 
    254.4919, 254.4873, 254.4856, 254.4849, 254.4843, 254.4827, 254.4838, 
    254.4834, 254.4844, 254.485, 254.4847, 254.4866, 254.4859, 254.4899, 
    254.4881, 254.4927, 254.4916, 254.4929, 254.4922, 254.4934, 254.4924, 
    254.4942, 254.4946, 254.4943, 254.4954, 254.4923, 254.4935, 254.4847, 
    254.4847, 254.485, 254.4839, 254.4839, 254.4829, 254.4838, 254.4841, 
    254.4851, 254.4856, 254.4861, 254.4873, 254.4885, 254.4903, 254.4917, 
    254.4925, 254.492, 254.4925, 254.4919, 254.4917, 254.4944, 254.4929, 
    254.4952, 254.4951, 254.494, 254.4951, 254.4848, 254.4845, 254.4835, 
    254.4843, 254.4828, 254.4836, 254.4841, 254.4859, 254.4863, 254.4867, 
    254.4874, 254.4883, 254.49, 254.4914, 254.4928, 254.4927, 254.4927, 
    254.493, 254.4923, 254.4931, 254.4933, 254.4929, 254.4951, 254.4944, 
    254.4951, 254.4947, 254.4846, 254.4851, 254.4848, 254.4853, 254.485, 
    254.4865, 254.487, 254.4892, 254.4883, 254.4898, 254.4885, 254.4887, 
    254.4898, 254.4886, 254.4913, 254.4894, 254.493, 254.4911, 254.4931, 
    254.4928, 254.4934, 254.4939, 254.4946, 254.4959, 254.4956, 254.4967, 
    254.4858, 254.4865, 254.4864, 254.4871, 254.4876, 254.4887, 254.4904, 
    254.4898, 254.491, 254.4912, 254.4894, 254.4905, 254.4869, 254.4875, 
    254.4871, 254.4859, 254.4899, 254.4878, 254.4917, 254.4905, 254.4939, 
    254.4922, 254.4954, 254.4968, 254.4981, 254.4996, 254.4868, 254.4864, 
    254.4872, 254.4882, 254.4893, 254.4906, 254.4908, 254.491, 254.4917, 
    254.4922, 254.4911, 254.4924, 254.4876, 254.4901, 254.4862, 254.4874, 
    254.4882, 254.4878, 254.4897, 254.4901, 254.4919, 254.491, 254.4964, 
    254.494, 254.5008, 254.4989, 254.4862, 254.4868, 254.4889, 254.4879, 
    254.4907, 254.4914, 254.492, 254.4927, 254.4928, 254.4932, 254.4925, 
    254.4932, 254.4906, 254.4918, 254.4886, 254.4894, 254.489, 254.4887, 
    254.4899, 254.4911, 254.4911, 254.4915, 254.4926, 254.4907, 254.4967, 
    254.493, 254.4875, 254.4886, 254.4888, 254.4883, 254.4913, 254.4902, 
    254.4932, 254.4924, 254.4937, 254.493, 254.493, 254.4921, 254.4916, 
    254.4903, 254.4892, 254.4884, 254.4886, 254.4895, 254.4912, 254.4928, 
    254.4924, 254.4936, 254.4905, 254.4918, 254.4913, 254.4926, 254.4897, 
    254.4921, 254.4891, 254.4894, 254.4902, 254.4919, 254.4922, 254.4926, 
    254.4924, 254.4912, 254.491, 254.4902, 254.49, 254.4893, 254.4888, 
    254.4893, 254.4898, 254.4912, 254.4925, 254.4939, 254.4943, 254.4959, 
    254.4946, 254.4967, 254.4948, 254.4982, 254.4923, 254.4948, 254.4902, 
    254.4908, 254.4916, 254.4937, 254.4926, 254.4939, 254.491, 254.4895, 
    254.4892, 254.4884, 254.4892, 254.4891, 254.4898, 254.4896, 254.4913, 
    254.4904, 254.4929, 254.4939, 254.4966, 254.4982, 254.4999, 254.5006, 
    254.5008, 254.5009 ;

 THBOT =
  253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 253.8605, 
    253.8605, 253.8605 ;

 TKE1 =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TLAI =
  0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312, 0.001119312, 0.001119312, 
    0.001119312, 0.001119312, 0.001119312 ;

 TLAKE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TOTCOLC =
  18.24019, 18.24018, 18.24018, 18.24017, 18.24018, 18.24017, 18.24019, 
    18.24018, 18.24018, 18.24019, 18.24015, 18.24017, 18.24013, 18.24014, 
    18.24011, 18.24013, 18.2401, 18.24011, 18.24009, 18.2401, 18.24008, 
    18.24009, 18.24007, 18.24008, 18.24008, 18.24009, 18.24016, 18.24015, 
    18.24017, 18.24016, 18.24016, 18.24018, 18.24018, 18.24019, 18.24019, 
    18.24018, 18.24016, 18.24017, 18.24015, 18.24015, 18.24014, 18.24014, 
    18.24011, 18.24012, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 
    18.24011, 18.2401, 18.24011, 18.24014, 18.24013, 18.24016, 18.24018, 
    18.24019, 18.24019, 18.24019, 18.24019, 18.24018, 18.24017, 18.24016, 
    18.24016, 18.24015, 18.24014, 18.24013, 18.24011, 18.24012, 18.24011, 
    18.2401, 18.2401, 18.2401, 18.24009, 18.24011, 18.2401, 18.24012, 
    18.24011, 18.24015, 18.24017, 18.24017, 18.24018, 18.24019, 18.24018, 
    18.24019, 18.24018, 18.24017, 18.24018, 18.24016, 18.24016, 18.24013, 
    18.24014, 18.2401, 18.24011, 18.2401, 18.24011, 18.2401, 18.24011, 
    18.24009, 18.24009, 18.24009, 18.24008, 18.24011, 18.2401, 18.24018, 
    18.24018, 18.24017, 18.24018, 18.24018, 18.24019, 18.24018, 18.24018, 
    18.24017, 18.24017, 18.24016, 18.24015, 18.24014, 18.24013, 18.24011, 
    18.24011, 18.24011, 18.24011, 18.24011, 18.24011, 18.24009, 18.2401, 
    18.24008, 18.24008, 18.24009, 18.24008, 18.24017, 18.24018, 18.24019, 
    18.24018, 18.24019, 18.24018, 18.24018, 18.24016, 18.24016, 18.24016, 
    18.24015, 18.24014, 18.24013, 18.24012, 18.2401, 18.2401, 18.2401, 
    18.2401, 18.24011, 18.2401, 18.2401, 18.2401, 18.24008, 18.24009, 
    18.24008, 18.24009, 18.24018, 18.24017, 18.24017, 18.24017, 18.24017, 
    18.24016, 18.24015, 18.24014, 18.24014, 18.24013, 18.24014, 18.24014, 
    18.24013, 18.24014, 18.24012, 18.24013, 18.2401, 18.24012, 18.2401, 
    18.2401, 18.2401, 18.2401, 18.24009, 18.24008, 18.24008, 18.24007, 
    18.24017, 18.24016, 18.24016, 18.24015, 18.24015, 18.24014, 18.24013, 
    18.24013, 18.24012, 18.24012, 18.24013, 18.24012, 18.24016, 18.24015, 
    18.24015, 18.24016, 18.24013, 18.24015, 18.24011, 18.24012, 18.2401, 
    18.24011, 18.24008, 18.24007, 18.24006, 18.24005, 18.24016, 18.24016, 
    18.24015, 18.24014, 18.24014, 18.24012, 18.24012, 18.24012, 18.24011, 
    18.24011, 18.24012, 18.24011, 18.24015, 18.24013, 18.24016, 18.24015, 
    18.24014, 18.24015, 18.24013, 18.24013, 18.24011, 18.24012, 18.24007, 
    18.24009, 18.24003, 18.24005, 18.24016, 18.24016, 18.24014, 18.24015, 
    18.24012, 18.24012, 18.24011, 18.2401, 18.2401, 18.2401, 18.24011, 
    18.2401, 18.24012, 18.24011, 18.24014, 18.24013, 18.24014, 18.24014, 
    18.24013, 18.24012, 18.24012, 18.24011, 18.2401, 18.24012, 18.24007, 
    18.2401, 18.24015, 18.24014, 18.24014, 18.24014, 18.24012, 18.24013, 
    18.2401, 18.24011, 18.2401, 18.2401, 18.2401, 18.24011, 18.24011, 
    18.24013, 18.24014, 18.24014, 18.24014, 18.24013, 18.24012, 18.2401, 
    18.24011, 18.2401, 18.24012, 18.24011, 18.24012, 18.24011, 18.24013, 
    18.24011, 18.24014, 18.24013, 18.24013, 18.24011, 18.24011, 18.2401, 
    18.24011, 18.24012, 18.24012, 18.24013, 18.24013, 18.24014, 18.24014, 
    18.24014, 18.24013, 18.24012, 18.24011, 18.2401, 18.24009, 18.24008, 
    18.24009, 18.24007, 18.24009, 18.24006, 18.24011, 18.24009, 18.24013, 
    18.24012, 18.24011, 18.2401, 18.24011, 18.2401, 18.24012, 18.24013, 
    18.24014, 18.24014, 18.24014, 18.24014, 18.24013, 18.24013, 18.24012, 
    18.24013, 18.2401, 18.2401, 18.24007, 18.24006, 18.24004, 18.24004, 
    18.24003, 18.24003 ;

 TOTCOLCH4 =
  4.605777e-06, 4.466226e-06, 4.493206e-06, 4.38175e-06, 4.443425e-06, 
    4.370667e-06, 4.577334e-06, 4.46072e-06, 4.535011e-06, 4.593142e-06, 
    4.169084e-06, 4.376809e-06, 3.958301e-06, 4.087137e-06, 3.767189e-06, 
    3.978217e-06, 3.725299e-06, 3.773212e-06, 3.629914e-06, 3.670697e-06, 
    3.490287e-06, 3.611165e-06, 3.398511e-06, 3.518981e-06, 3.499997e-06, 
    3.615185e-06, 4.334646e-06, 4.194689e-06, 4.343001e-06, 4.322898e-06, 
    4.331916e-06, 4.442144e-06, 4.498158e-06, 4.61653e-06, 4.59494e-06, 
    4.508053e-06, 4.313873e-06, 4.379361e-06, 4.215201e-06, 4.218877e-06, 
    4.039437e-06, 4.119896e-06, 3.823744e-06, 3.906865e-06, 3.66899e-06, 
    3.728144e-06, 3.671757e-06, 3.688813e-06, 3.671535e-06, 3.758474e-06, 
    3.721106e-06, 3.798046e-06, 4.104769e-06, 4.013466e-06, 4.288572e-06, 
    4.457991e-06, 4.572189e-06, 4.654e-06, 4.642395e-06, 4.620305e-06, 
    4.507546e-06, 4.402686e-06, 4.323523e-06, 4.270933e-06, 4.219406e-06, 
    4.065164e-06, 3.984632e-06, 3.807033e-06, 3.838812e-06, 3.785058e-06, 
    3.734054e-06, 3.649151e-06, 3.663063e-06, 3.625883e-06, 3.786478e-06, 
    3.679373e-06, 3.856966e-06, 3.807997e-06, 4.205407e-06, 4.361651e-06, 
    4.428813e-06, 4.488013e-06, 4.63348e-06, 4.532798e-06, 4.572369e-06, 
    4.478491e-06, 4.419291e-06, 4.448527e-06, 4.269499e-06, 4.338701e-06, 
    3.979882e-06, 4.132684e-06, 3.739986e-06, 3.83228e-06, 3.718024e-06, 
    3.776123e-06, 3.676834e-06, 3.766137e-06, 3.612095e-06, 3.578957e-06, 
    3.601586e-06, 3.515046e-06, 3.771116e-06, 3.671754e-06, 4.449346e-06, 
    4.444571e-06, 4.422361e-06, 4.520365e-06, 4.526394e-06, 4.617121e-06, 
    4.536357e-06, 4.502155e-06, 4.415873e-06, 4.365186e-06, 4.317252e-06, 
    4.212712e-06, 4.097348e-06, 3.938536e-06, 3.826264e-06, 3.751863e-06, 
    3.797405e-06, 3.757184e-06, 3.802159e-06, 3.823327e-06, 3.591354e-06, 
    3.720756e-06, 3.527431e-06, 3.538e-06, 3.625e-06, 3.536808e-06, 
    4.44122e-06, 4.468719e-06, 4.564773e-06, 4.489524e-06, 4.62705e-06, 
    4.549835e-06, 4.505698e-06, 4.337241e-06, 4.30063e-06, 4.266796e-06, 
    4.200343e-06, 4.11576e-06, 3.969307e-06, 3.843908e-06, 3.731099e-06, 
    3.739311e-06, 3.736418e-06, 3.711415e-06, 3.773491e-06, 3.701271e-06, 
    3.689211e-06, 3.720776e-06, 3.539417e-06, 3.590787e-06, 3.538225e-06, 
    3.571628e-06, 4.459773e-06, 4.41359e-06, 4.438518e-06, 4.391693e-06, 
    4.424655e-06, 4.278937e-06, 4.235683e-06, 4.03599e-06, 4.117415e-06, 
    3.988194e-06, 4.104204e-06, 4.083533e-06, 3.983994e-06, 4.097898e-06, 
    3.850765e-06, 4.017515e-06, 3.710444e-06, 3.874088e-06, 3.7003e-06, 
    3.731583e-06, 3.679861e-06, 3.633827e-06, 3.576314e-06, 3.471342e-06, 
    3.495517e-06, 3.408605e-06, 4.345151e-06, 4.285995e-06, 4.291196e-06, 
    4.229657e-06, 4.184407e-06, 4.08711e-06, 3.933273e-06, 3.990801e-06, 
    3.885497e-06, 3.864513e-06, 4.024619e-06, 3.925948e-06, 4.246618e-06, 
    4.194012e-06, 4.225303e-06, 4.340467e-06, 3.9775e-06, 4.161944e-06, 
    3.82442e-06, 3.922059e-06, 3.640372e-06, 3.779209e-06, 3.508858e-06, 
    3.396215e-06, 3.291864e-06, 3.171903e-06, 4.253875e-06, 4.293891e-06, 
    4.222369e-06, 4.124312e-06, 4.034305e-06, 3.916069e-06, 3.904069e-06, 
    3.882131e-06, 3.825587e-06, 3.778345e-06, 3.8752e-06, 3.766547e-06, 
    4.18184e-06, 3.961677e-06, 4.309058e-06, 4.203026e-06, 4.130065e-06, 
    4.162006e-06, 3.997403e-06, 3.959056e-06, 3.805012e-06, 3.884289e-06, 
    3.423845e-06, 3.624129e-06, 3.082055e-06, 3.229216e-06, 4.307911e-06, 
    4.254015e-06, 4.068866e-06, 4.156487e-06, 3.908238e-06, 3.848227e-06, 
    3.799771e-06, 3.738242e-06, 3.731633e-06, 3.695434e-06, 3.75484e-06, 
    3.697775e-06, 3.915819e-06, 3.81765e-06, 4.089846e-06, 4.022784e-06, 
    4.053573e-06, 4.087466e-06, 3.983284e-06, 3.873664e-06, 3.871349e-06, 
    3.836512e-06, 3.739123e-06, 3.907247e-06, 3.398376e-06, 3.70862e-06, 
    4.1956e-06, 4.093309e-06, 4.078808e-06, 4.118227e-06, 3.854223e-06, 
    3.948935e-06, 3.696316e-06, 3.763813e-06, 3.653528e-06, 3.708134e-06, 
    3.7162e-06, 3.786975e-06, 3.831355e-06, 3.944566e-06, 4.037823e-06, 
    4.112501e-06, 4.095081e-06, 4.013246e-06, 3.867008e-06, 3.731029e-06, 
    3.760617e-06, 3.661855e-06, 3.925998e-06, 3.814171e-06, 3.857208e-06, 
    3.745473e-06, 3.992333e-06, 3.781612e-06, 4.047049e-06, 4.023442e-06, 
    3.950826e-06, 3.806634e-06, 3.775092e-06, 3.74153e-06, 3.762226e-06, 
    3.863331e-06, 3.880021e-06, 3.952586e-06, 3.972727e-06, 4.028577e-06, 
    4.075085e-06, 4.03258e-06, 3.988162e-06, 3.863293e-06, 3.752362e-06, 
    3.633171e-06, 3.604288e-06, 3.467864e-06, 3.578712e-06, 3.396682e-06, 
    3.551126e-06, 3.285898e-06, 3.769584e-06, 3.55574e-06, 3.94754e-06, 
    3.904403e-06, 3.826933e-06, 3.652055e-06, 3.745995e-06, 3.636251e-06, 
    3.880677e-06, 4.01043e-06, 4.044341e-06, 4.10794e-06, 4.042893e-06, 
    4.048165e-06, 3.986336e-06, 4.006158e-06, 3.859179e-06, 3.93781e-06, 
    3.7164e-06, 3.637115e-06, 3.417659e-06, 3.286395e-06, 3.155379e-06, 
    3.098368e-06, 3.081119e-06, 3.073922e-06 ;

 TOTCOLN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTECOSYSC =
  18.24019, 18.24018, 18.24018, 18.24017, 18.24018, 18.24017, 18.24019, 
    18.24018, 18.24018, 18.24019, 18.24015, 18.24017, 18.24013, 18.24014, 
    18.24011, 18.24013, 18.2401, 18.24011, 18.24009, 18.2401, 18.24008, 
    18.24009, 18.24007, 18.24008, 18.24008, 18.24009, 18.24016, 18.24015, 
    18.24017, 18.24016, 18.24016, 18.24018, 18.24018, 18.24019, 18.24019, 
    18.24018, 18.24016, 18.24017, 18.24015, 18.24015, 18.24014, 18.24014, 
    18.24011, 18.24012, 18.2401, 18.2401, 18.2401, 18.2401, 18.2401, 
    18.24011, 18.2401, 18.24011, 18.24014, 18.24013, 18.24016, 18.24018, 
    18.24019, 18.24019, 18.24019, 18.24019, 18.24018, 18.24017, 18.24016, 
    18.24016, 18.24015, 18.24014, 18.24013, 18.24011, 18.24012, 18.24011, 
    18.2401, 18.2401, 18.2401, 18.24009, 18.24011, 18.2401, 18.24012, 
    18.24011, 18.24015, 18.24017, 18.24017, 18.24018, 18.24019, 18.24018, 
    18.24019, 18.24018, 18.24017, 18.24018, 18.24016, 18.24016, 18.24013, 
    18.24014, 18.2401, 18.24011, 18.2401, 18.24011, 18.2401, 18.24011, 
    18.24009, 18.24009, 18.24009, 18.24008, 18.24011, 18.2401, 18.24018, 
    18.24018, 18.24017, 18.24018, 18.24018, 18.24019, 18.24018, 18.24018, 
    18.24017, 18.24017, 18.24016, 18.24015, 18.24014, 18.24013, 18.24011, 
    18.24011, 18.24011, 18.24011, 18.24011, 18.24011, 18.24009, 18.2401, 
    18.24008, 18.24008, 18.24009, 18.24008, 18.24017, 18.24018, 18.24019, 
    18.24018, 18.24019, 18.24018, 18.24018, 18.24016, 18.24016, 18.24016, 
    18.24015, 18.24014, 18.24013, 18.24012, 18.2401, 18.2401, 18.2401, 
    18.2401, 18.24011, 18.2401, 18.2401, 18.2401, 18.24008, 18.24009, 
    18.24008, 18.24009, 18.24018, 18.24017, 18.24017, 18.24017, 18.24017, 
    18.24016, 18.24015, 18.24014, 18.24014, 18.24013, 18.24014, 18.24014, 
    18.24013, 18.24014, 18.24012, 18.24013, 18.2401, 18.24012, 18.2401, 
    18.2401, 18.2401, 18.2401, 18.24009, 18.24008, 18.24008, 18.24007, 
    18.24017, 18.24016, 18.24016, 18.24015, 18.24015, 18.24014, 18.24013, 
    18.24013, 18.24012, 18.24012, 18.24013, 18.24012, 18.24016, 18.24015, 
    18.24015, 18.24016, 18.24013, 18.24015, 18.24011, 18.24012, 18.2401, 
    18.24011, 18.24008, 18.24007, 18.24006, 18.24005, 18.24016, 18.24016, 
    18.24015, 18.24014, 18.24014, 18.24012, 18.24012, 18.24012, 18.24011, 
    18.24011, 18.24012, 18.24011, 18.24015, 18.24013, 18.24016, 18.24015, 
    18.24014, 18.24015, 18.24013, 18.24013, 18.24011, 18.24012, 18.24007, 
    18.24009, 18.24003, 18.24005, 18.24016, 18.24016, 18.24014, 18.24015, 
    18.24012, 18.24012, 18.24011, 18.2401, 18.2401, 18.2401, 18.24011, 
    18.2401, 18.24012, 18.24011, 18.24014, 18.24013, 18.24014, 18.24014, 
    18.24013, 18.24012, 18.24012, 18.24011, 18.2401, 18.24012, 18.24007, 
    18.2401, 18.24015, 18.24014, 18.24014, 18.24014, 18.24012, 18.24013, 
    18.2401, 18.24011, 18.2401, 18.2401, 18.2401, 18.24011, 18.24011, 
    18.24013, 18.24014, 18.24014, 18.24014, 18.24013, 18.24012, 18.2401, 
    18.24011, 18.2401, 18.24012, 18.24011, 18.24012, 18.24011, 18.24013, 
    18.24011, 18.24014, 18.24013, 18.24013, 18.24011, 18.24011, 18.2401, 
    18.24011, 18.24012, 18.24012, 18.24013, 18.24013, 18.24014, 18.24014, 
    18.24014, 18.24013, 18.24012, 18.24011, 18.2401, 18.24009, 18.24008, 
    18.24009, 18.24007, 18.24009, 18.24006, 18.24011, 18.24009, 18.24013, 
    18.24012, 18.24011, 18.2401, 18.24011, 18.2401, 18.24012, 18.24013, 
    18.24014, 18.24014, 18.24014, 18.24014, 18.24013, 18.24013, 18.24012, 
    18.24013, 18.2401, 18.2401, 18.24007, 18.24006, 18.24004, 18.24004, 
    18.24003, 18.24003 ;

 TOTECOSYSN =
  1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 1.806727, 
    1.806727, 1.806727 ;

 TOTLITC =
  5.976298e-05, 5.976283e-05, 5.976286e-05, 5.976274e-05, 5.976281e-05, 
    5.976273e-05, 5.976295e-05, 5.976282e-05, 5.97629e-05, 5.976297e-05, 
    5.976251e-05, 5.976273e-05, 5.976227e-05, 5.976242e-05, 5.976206e-05, 
    5.97623e-05, 5.976201e-05, 5.976206e-05, 5.97619e-05, 5.976194e-05, 
    5.976173e-05, 5.976187e-05, 5.976162e-05, 5.976177e-05, 5.976174e-05, 
    5.976188e-05, 5.976269e-05, 5.976254e-05, 5.97627e-05, 5.976267e-05, 
    5.976269e-05, 5.976281e-05, 5.976286e-05, 5.976299e-05, 5.976297e-05, 
    5.976288e-05, 5.976267e-05, 5.976274e-05, 5.976256e-05, 5.976256e-05, 
    5.976236e-05, 5.976245e-05, 5.976212e-05, 5.976221e-05, 5.976194e-05, 
    5.976201e-05, 5.976194e-05, 5.976197e-05, 5.976194e-05, 5.976205e-05, 
    5.9762e-05, 5.976209e-05, 5.976243e-05, 5.976234e-05, 5.976264e-05, 
    5.976282e-05, 5.976294e-05, 5.976303e-05, 5.976302e-05, 5.9763e-05, 
    5.976288e-05, 5.976276e-05, 5.976267e-05, 5.976262e-05, 5.976256e-05, 
    5.976239e-05, 5.97623e-05, 5.97621e-05, 5.976214e-05, 5.976207e-05, 
    5.976202e-05, 5.976192e-05, 5.976193e-05, 5.976189e-05, 5.976208e-05, 
    5.976195e-05, 5.976216e-05, 5.97621e-05, 5.976255e-05, 5.976272e-05, 
    5.976279e-05, 5.976285e-05, 5.976301e-05, 5.97629e-05, 5.976294e-05, 
    5.976284e-05, 5.976278e-05, 5.976281e-05, 5.976262e-05, 5.976269e-05, 
    5.97623e-05, 5.976247e-05, 5.976202e-05, 5.976213e-05, 5.9762e-05, 
    5.976206e-05, 5.976195e-05, 5.976205e-05, 5.976187e-05, 5.976183e-05, 
    5.976186e-05, 5.976176e-05, 5.976206e-05, 5.976194e-05, 5.976281e-05, 
    5.976281e-05, 5.976278e-05, 5.976289e-05, 5.976289e-05, 5.976299e-05, 
    5.97629e-05, 5.976287e-05, 5.976278e-05, 5.976272e-05, 5.976267e-05, 
    5.976255e-05, 5.976243e-05, 5.976225e-05, 5.976212e-05, 5.976204e-05, 
    5.976209e-05, 5.976204e-05, 5.97621e-05, 5.976212e-05, 5.976185e-05, 
    5.9762e-05, 5.976178e-05, 5.976179e-05, 5.976189e-05, 5.976179e-05, 
    5.97628e-05, 5.976283e-05, 5.976293e-05, 5.976285e-05, 5.9763e-05, 
    5.976292e-05, 5.976287e-05, 5.976269e-05, 5.976265e-05, 5.976261e-05, 
    5.976254e-05, 5.976245e-05, 5.976229e-05, 5.976214e-05, 5.976201e-05, 
    5.976202e-05, 5.976202e-05, 5.976199e-05, 5.976206e-05, 5.976198e-05, 
    5.976197e-05, 5.9762e-05, 5.976179e-05, 5.976185e-05, 5.976179e-05, 
    5.976183e-05, 5.976282e-05, 5.976277e-05, 5.97628e-05, 5.976275e-05, 
    5.976278e-05, 5.976263e-05, 5.976258e-05, 5.976236e-05, 5.976245e-05, 
    5.976231e-05, 5.976243e-05, 5.976241e-05, 5.97623e-05, 5.976243e-05, 
    5.976215e-05, 5.976234e-05, 5.976199e-05, 5.976218e-05, 5.976198e-05, 
    5.976201e-05, 5.976195e-05, 5.97619e-05, 5.976183e-05, 5.976171e-05, 
    5.976174e-05, 5.976163e-05, 5.97627e-05, 5.976263e-05, 5.976264e-05, 
    5.976257e-05, 5.976253e-05, 5.976242e-05, 5.976225e-05, 5.976231e-05, 
    5.976219e-05, 5.976217e-05, 5.976235e-05, 5.976223e-05, 5.976259e-05, 
    5.976254e-05, 5.976257e-05, 5.976269e-05, 5.976229e-05, 5.97625e-05, 
    5.976212e-05, 5.976223e-05, 5.976191e-05, 5.976207e-05, 5.976175e-05, 
    5.976162e-05, 5.976149e-05, 5.976134e-05, 5.97626e-05, 5.976265e-05, 
    5.976257e-05, 5.976246e-05, 5.976236e-05, 5.976222e-05, 5.976221e-05, 
    5.976219e-05, 5.976212e-05, 5.976207e-05, 5.976218e-05, 5.976205e-05, 
    5.976252e-05, 5.976228e-05, 5.976266e-05, 5.976254e-05, 5.976246e-05, 
    5.97625e-05, 5.976232e-05, 5.976227e-05, 5.97621e-05, 5.976219e-05, 
    5.976165e-05, 5.976189e-05, 5.976123e-05, 5.976141e-05, 5.976266e-05, 
    5.97626e-05, 5.97624e-05, 5.976249e-05, 5.976222e-05, 5.976215e-05, 
    5.976209e-05, 5.976202e-05, 5.976201e-05, 5.976197e-05, 5.976204e-05, 
    5.976198e-05, 5.976222e-05, 5.976211e-05, 5.976242e-05, 5.976234e-05, 
    5.976238e-05, 5.976242e-05, 5.97623e-05, 5.976218e-05, 5.976217e-05, 
    5.976213e-05, 5.976202e-05, 5.976222e-05, 5.976162e-05, 5.976199e-05, 
    5.976254e-05, 5.976242e-05, 5.976241e-05, 5.976245e-05, 5.976215e-05, 
    5.976226e-05, 5.976197e-05, 5.976205e-05, 5.976192e-05, 5.976199e-05, 
    5.976199e-05, 5.976208e-05, 5.976213e-05, 5.976226e-05, 5.976236e-05, 
    5.976245e-05, 5.976243e-05, 5.976233e-05, 5.976217e-05, 5.976201e-05, 
    5.976205e-05, 5.976193e-05, 5.976223e-05, 5.976211e-05, 5.976216e-05, 
    5.976203e-05, 5.976231e-05, 5.976207e-05, 5.976237e-05, 5.976235e-05, 
    5.976226e-05, 5.97621e-05, 5.976206e-05, 5.976202e-05, 5.976205e-05, 
    5.976217e-05, 5.976218e-05, 5.976227e-05, 5.976229e-05, 5.976235e-05, 
    5.97624e-05, 5.976235e-05, 5.976231e-05, 5.976217e-05, 5.976204e-05, 
    5.97619e-05, 5.976186e-05, 5.97617e-05, 5.976183e-05, 5.976162e-05, 
    5.97618e-05, 5.976148e-05, 5.976206e-05, 5.976181e-05, 5.976226e-05, 
    5.976221e-05, 5.976212e-05, 5.976192e-05, 5.976203e-05, 5.97619e-05, 
    5.976218e-05, 5.976233e-05, 5.976237e-05, 5.976244e-05, 5.976237e-05, 
    5.976237e-05, 5.97623e-05, 5.976233e-05, 5.976216e-05, 5.976225e-05, 
    5.976199e-05, 5.97619e-05, 5.976164e-05, 5.976149e-05, 5.976132e-05, 
    5.976125e-05, 5.976123e-05, 5.976122e-05 ;

 TOTLITC_1m =
  5.976298e-05, 5.976283e-05, 5.976286e-05, 5.976274e-05, 5.976281e-05, 
    5.976273e-05, 5.976295e-05, 5.976282e-05, 5.97629e-05, 5.976297e-05, 
    5.976251e-05, 5.976273e-05, 5.976227e-05, 5.976242e-05, 5.976206e-05, 
    5.97623e-05, 5.976201e-05, 5.976206e-05, 5.97619e-05, 5.976194e-05, 
    5.976173e-05, 5.976187e-05, 5.976162e-05, 5.976177e-05, 5.976174e-05, 
    5.976188e-05, 5.976269e-05, 5.976254e-05, 5.97627e-05, 5.976267e-05, 
    5.976269e-05, 5.976281e-05, 5.976286e-05, 5.976299e-05, 5.976297e-05, 
    5.976288e-05, 5.976267e-05, 5.976274e-05, 5.976256e-05, 5.976256e-05, 
    5.976236e-05, 5.976245e-05, 5.976212e-05, 5.976221e-05, 5.976194e-05, 
    5.976201e-05, 5.976194e-05, 5.976197e-05, 5.976194e-05, 5.976205e-05, 
    5.9762e-05, 5.976209e-05, 5.976243e-05, 5.976234e-05, 5.976264e-05, 
    5.976282e-05, 5.976294e-05, 5.976303e-05, 5.976302e-05, 5.9763e-05, 
    5.976288e-05, 5.976276e-05, 5.976267e-05, 5.976262e-05, 5.976256e-05, 
    5.976239e-05, 5.97623e-05, 5.97621e-05, 5.976214e-05, 5.976207e-05, 
    5.976202e-05, 5.976192e-05, 5.976193e-05, 5.976189e-05, 5.976208e-05, 
    5.976195e-05, 5.976216e-05, 5.97621e-05, 5.976255e-05, 5.976272e-05, 
    5.976279e-05, 5.976285e-05, 5.976301e-05, 5.97629e-05, 5.976294e-05, 
    5.976284e-05, 5.976278e-05, 5.976281e-05, 5.976262e-05, 5.976269e-05, 
    5.97623e-05, 5.976247e-05, 5.976202e-05, 5.976213e-05, 5.9762e-05, 
    5.976206e-05, 5.976195e-05, 5.976205e-05, 5.976187e-05, 5.976183e-05, 
    5.976186e-05, 5.976176e-05, 5.976206e-05, 5.976194e-05, 5.976281e-05, 
    5.976281e-05, 5.976278e-05, 5.976289e-05, 5.976289e-05, 5.976299e-05, 
    5.97629e-05, 5.976287e-05, 5.976278e-05, 5.976272e-05, 5.976267e-05, 
    5.976255e-05, 5.976243e-05, 5.976225e-05, 5.976212e-05, 5.976204e-05, 
    5.976209e-05, 5.976204e-05, 5.97621e-05, 5.976212e-05, 5.976185e-05, 
    5.9762e-05, 5.976178e-05, 5.976179e-05, 5.976189e-05, 5.976179e-05, 
    5.97628e-05, 5.976283e-05, 5.976293e-05, 5.976285e-05, 5.9763e-05, 
    5.976292e-05, 5.976287e-05, 5.976269e-05, 5.976265e-05, 5.976261e-05, 
    5.976254e-05, 5.976245e-05, 5.976229e-05, 5.976214e-05, 5.976201e-05, 
    5.976202e-05, 5.976202e-05, 5.976199e-05, 5.976206e-05, 5.976198e-05, 
    5.976197e-05, 5.9762e-05, 5.976179e-05, 5.976185e-05, 5.976179e-05, 
    5.976183e-05, 5.976282e-05, 5.976277e-05, 5.97628e-05, 5.976275e-05, 
    5.976278e-05, 5.976263e-05, 5.976258e-05, 5.976236e-05, 5.976245e-05, 
    5.976231e-05, 5.976243e-05, 5.976241e-05, 5.97623e-05, 5.976243e-05, 
    5.976215e-05, 5.976234e-05, 5.976199e-05, 5.976218e-05, 5.976198e-05, 
    5.976201e-05, 5.976195e-05, 5.97619e-05, 5.976183e-05, 5.976171e-05, 
    5.976174e-05, 5.976163e-05, 5.97627e-05, 5.976263e-05, 5.976264e-05, 
    5.976257e-05, 5.976253e-05, 5.976242e-05, 5.976225e-05, 5.976231e-05, 
    5.976219e-05, 5.976217e-05, 5.976235e-05, 5.976223e-05, 5.976259e-05, 
    5.976254e-05, 5.976257e-05, 5.976269e-05, 5.976229e-05, 5.97625e-05, 
    5.976212e-05, 5.976223e-05, 5.976191e-05, 5.976207e-05, 5.976175e-05, 
    5.976162e-05, 5.976149e-05, 5.976134e-05, 5.97626e-05, 5.976265e-05, 
    5.976257e-05, 5.976246e-05, 5.976236e-05, 5.976222e-05, 5.976221e-05, 
    5.976219e-05, 5.976212e-05, 5.976207e-05, 5.976218e-05, 5.976205e-05, 
    5.976252e-05, 5.976228e-05, 5.976266e-05, 5.976254e-05, 5.976246e-05, 
    5.97625e-05, 5.976232e-05, 5.976227e-05, 5.97621e-05, 5.976219e-05, 
    5.976165e-05, 5.976189e-05, 5.976123e-05, 5.976141e-05, 5.976266e-05, 
    5.97626e-05, 5.97624e-05, 5.976249e-05, 5.976222e-05, 5.976215e-05, 
    5.976209e-05, 5.976202e-05, 5.976201e-05, 5.976197e-05, 5.976204e-05, 
    5.976198e-05, 5.976222e-05, 5.976211e-05, 5.976242e-05, 5.976234e-05, 
    5.976238e-05, 5.976242e-05, 5.97623e-05, 5.976218e-05, 5.976217e-05, 
    5.976213e-05, 5.976202e-05, 5.976222e-05, 5.976162e-05, 5.976199e-05, 
    5.976254e-05, 5.976242e-05, 5.976241e-05, 5.976245e-05, 5.976215e-05, 
    5.976226e-05, 5.976197e-05, 5.976205e-05, 5.976192e-05, 5.976199e-05, 
    5.976199e-05, 5.976208e-05, 5.976213e-05, 5.976226e-05, 5.976236e-05, 
    5.976245e-05, 5.976243e-05, 5.976233e-05, 5.976217e-05, 5.976201e-05, 
    5.976205e-05, 5.976193e-05, 5.976223e-05, 5.976211e-05, 5.976216e-05, 
    5.976203e-05, 5.976231e-05, 5.976207e-05, 5.976237e-05, 5.976235e-05, 
    5.976226e-05, 5.97621e-05, 5.976206e-05, 5.976202e-05, 5.976205e-05, 
    5.976217e-05, 5.976218e-05, 5.976227e-05, 5.976229e-05, 5.976235e-05, 
    5.97624e-05, 5.976235e-05, 5.976231e-05, 5.976217e-05, 5.976204e-05, 
    5.97619e-05, 5.976186e-05, 5.97617e-05, 5.976183e-05, 5.976162e-05, 
    5.97618e-05, 5.976148e-05, 5.976206e-05, 5.976181e-05, 5.976226e-05, 
    5.976221e-05, 5.976212e-05, 5.976192e-05, 5.976203e-05, 5.97619e-05, 
    5.976218e-05, 5.976233e-05, 5.976237e-05, 5.976244e-05, 5.976237e-05, 
    5.976237e-05, 5.97623e-05, 5.976233e-05, 5.976216e-05, 5.976225e-05, 
    5.976199e-05, 5.97619e-05, 5.976164e-05, 5.976149e-05, 5.976132e-05, 
    5.976125e-05, 5.976123e-05, 5.976122e-05 ;

 TOTLITN =
  1.375956e-06, 1.375952e-06, 1.375952e-06, 1.375949e-06, 1.375951e-06, 
    1.375949e-06, 1.375955e-06, 1.375951e-06, 1.375954e-06, 1.375955e-06, 
    1.375942e-06, 1.375949e-06, 1.375936e-06, 1.37594e-06, 1.37593e-06, 
    1.375936e-06, 1.375928e-06, 1.37593e-06, 1.375925e-06, 1.375927e-06, 
    1.375921e-06, 1.375925e-06, 1.375917e-06, 1.375922e-06, 1.375921e-06, 
    1.375925e-06, 1.375948e-06, 1.375943e-06, 1.375948e-06, 1.375947e-06, 
    1.375947e-06, 1.375951e-06, 1.375952e-06, 1.375956e-06, 1.375955e-06, 
    1.375953e-06, 1.375947e-06, 1.375949e-06, 1.375944e-06, 1.375944e-06, 
    1.375938e-06, 1.375941e-06, 1.375932e-06, 1.375934e-06, 1.375927e-06, 
    1.375928e-06, 1.375927e-06, 1.375927e-06, 1.375927e-06, 1.375929e-06, 
    1.375928e-06, 1.375931e-06, 1.37594e-06, 1.375938e-06, 1.375946e-06, 
    1.375951e-06, 1.375955e-06, 1.375957e-06, 1.375957e-06, 1.375956e-06, 
    1.375953e-06, 1.37595e-06, 1.375947e-06, 1.375946e-06, 1.375944e-06, 
    1.375939e-06, 1.375937e-06, 1.375931e-06, 1.375932e-06, 1.37593e-06, 
    1.375929e-06, 1.375926e-06, 1.375926e-06, 1.375925e-06, 1.37593e-06, 
    1.375927e-06, 1.375933e-06, 1.375931e-06, 1.375944e-06, 1.375948e-06, 
    1.37595e-06, 1.375952e-06, 1.375957e-06, 1.375954e-06, 1.375955e-06, 
    1.375952e-06, 1.37595e-06, 1.375951e-06, 1.375946e-06, 1.375948e-06, 
    1.375937e-06, 1.375941e-06, 1.375929e-06, 1.375932e-06, 1.375928e-06, 
    1.37593e-06, 1.375927e-06, 1.37593e-06, 1.375925e-06, 1.375923e-06, 
    1.375924e-06, 1.375921e-06, 1.37593e-06, 1.375927e-06, 1.375951e-06, 
    1.375951e-06, 1.37595e-06, 1.375953e-06, 1.375953e-06, 1.375956e-06, 
    1.375954e-06, 1.375953e-06, 1.37595e-06, 1.375949e-06, 1.375947e-06, 
    1.375944e-06, 1.37594e-06, 1.375935e-06, 1.375932e-06, 1.375929e-06, 
    1.375931e-06, 1.375929e-06, 1.375931e-06, 1.375932e-06, 1.375924e-06, 
    1.375928e-06, 1.375922e-06, 1.375922e-06, 1.375925e-06, 1.375922e-06, 
    1.375951e-06, 1.375952e-06, 1.375955e-06, 1.375952e-06, 1.375956e-06, 
    1.375954e-06, 1.375953e-06, 1.375948e-06, 1.375946e-06, 1.375945e-06, 
    1.375943e-06, 1.375941e-06, 1.375936e-06, 1.375932e-06, 1.375928e-06, 
    1.375929e-06, 1.375929e-06, 1.375928e-06, 1.37593e-06, 1.375928e-06, 
    1.375927e-06, 1.375928e-06, 1.375922e-06, 1.375924e-06, 1.375922e-06, 
    1.375923e-06, 1.375951e-06, 1.37595e-06, 1.375951e-06, 1.375949e-06, 
    1.37595e-06, 1.375946e-06, 1.375945e-06, 1.375938e-06, 1.375941e-06, 
    1.375937e-06, 1.37594e-06, 1.37594e-06, 1.375937e-06, 1.37594e-06, 
    1.375932e-06, 1.375938e-06, 1.375928e-06, 1.375933e-06, 1.375928e-06, 
    1.375929e-06, 1.375927e-06, 1.375925e-06, 1.375923e-06, 1.37592e-06, 
    1.375921e-06, 1.375918e-06, 1.375948e-06, 1.375946e-06, 1.375946e-06, 
    1.375944e-06, 1.375943e-06, 1.37594e-06, 1.375935e-06, 1.375937e-06, 
    1.375933e-06, 1.375933e-06, 1.375938e-06, 1.375935e-06, 1.375945e-06, 
    1.375943e-06, 1.375944e-06, 1.375948e-06, 1.375936e-06, 1.375942e-06, 
    1.375932e-06, 1.375935e-06, 1.375926e-06, 1.37593e-06, 1.375921e-06, 
    1.375917e-06, 1.375914e-06, 1.37591e-06, 1.375945e-06, 1.375946e-06, 
    1.375944e-06, 1.375941e-06, 1.375938e-06, 1.375935e-06, 1.375934e-06, 
    1.375933e-06, 1.375932e-06, 1.37593e-06, 1.375933e-06, 1.37593e-06, 
    1.375943e-06, 1.375936e-06, 1.375947e-06, 1.375943e-06, 1.375941e-06, 
    1.375942e-06, 1.375937e-06, 1.375936e-06, 1.375931e-06, 1.375933e-06, 
    1.375918e-06, 1.375925e-06, 1.375906e-06, 1.375912e-06, 1.375947e-06, 
    1.375945e-06, 1.375939e-06, 1.375942e-06, 1.375934e-06, 1.375932e-06, 
    1.375931e-06, 1.375929e-06, 1.375929e-06, 1.375927e-06, 1.375929e-06, 
    1.375927e-06, 1.375935e-06, 1.375931e-06, 1.37594e-06, 1.375938e-06, 
    1.375939e-06, 1.37594e-06, 1.375937e-06, 1.375933e-06, 1.375933e-06, 
    1.375932e-06, 1.375929e-06, 1.375934e-06, 1.375917e-06, 1.375928e-06, 
    1.375943e-06, 1.37594e-06, 1.37594e-06, 1.375941e-06, 1.375932e-06, 
    1.375936e-06, 1.375927e-06, 1.37593e-06, 1.375926e-06, 1.375928e-06, 
    1.375928e-06, 1.37593e-06, 1.375932e-06, 1.375935e-06, 1.375938e-06, 
    1.375941e-06, 1.37594e-06, 1.375938e-06, 1.375933e-06, 1.375928e-06, 
    1.37593e-06, 1.375926e-06, 1.375935e-06, 1.375931e-06, 1.375933e-06, 
    1.375929e-06, 1.375937e-06, 1.37593e-06, 1.375939e-06, 1.375938e-06, 
    1.375936e-06, 1.375931e-06, 1.37593e-06, 1.375929e-06, 1.37593e-06, 
    1.375933e-06, 1.375933e-06, 1.375936e-06, 1.375936e-06, 1.375938e-06, 
    1.37594e-06, 1.375938e-06, 1.375937e-06, 1.375933e-06, 1.375929e-06, 
    1.375925e-06, 1.375924e-06, 1.37592e-06, 1.375923e-06, 1.375917e-06, 
    1.375923e-06, 1.375914e-06, 1.37593e-06, 1.375923e-06, 1.375936e-06, 
    1.375934e-06, 1.375932e-06, 1.375926e-06, 1.375929e-06, 1.375925e-06, 
    1.375933e-06, 1.375937e-06, 1.375939e-06, 1.375941e-06, 1.375938e-06, 
    1.375939e-06, 1.375937e-06, 1.375937e-06, 1.375933e-06, 1.375935e-06, 
    1.375928e-06, 1.375925e-06, 1.375918e-06, 1.375914e-06, 1.375909e-06, 
    1.375907e-06, 1.375906e-06, 1.375906e-06 ;

 TOTLITN_1m =
  1.375956e-06, 1.375952e-06, 1.375952e-06, 1.375949e-06, 1.375951e-06, 
    1.375949e-06, 1.375955e-06, 1.375951e-06, 1.375954e-06, 1.375955e-06, 
    1.375942e-06, 1.375949e-06, 1.375936e-06, 1.37594e-06, 1.37593e-06, 
    1.375936e-06, 1.375928e-06, 1.37593e-06, 1.375925e-06, 1.375927e-06, 
    1.375921e-06, 1.375925e-06, 1.375917e-06, 1.375922e-06, 1.375921e-06, 
    1.375925e-06, 1.375948e-06, 1.375943e-06, 1.375948e-06, 1.375947e-06, 
    1.375947e-06, 1.375951e-06, 1.375952e-06, 1.375956e-06, 1.375955e-06, 
    1.375953e-06, 1.375947e-06, 1.375949e-06, 1.375944e-06, 1.375944e-06, 
    1.375938e-06, 1.375941e-06, 1.375932e-06, 1.375934e-06, 1.375927e-06, 
    1.375928e-06, 1.375927e-06, 1.375927e-06, 1.375927e-06, 1.375929e-06, 
    1.375928e-06, 1.375931e-06, 1.37594e-06, 1.375938e-06, 1.375946e-06, 
    1.375951e-06, 1.375955e-06, 1.375957e-06, 1.375957e-06, 1.375956e-06, 
    1.375953e-06, 1.37595e-06, 1.375947e-06, 1.375946e-06, 1.375944e-06, 
    1.375939e-06, 1.375937e-06, 1.375931e-06, 1.375932e-06, 1.37593e-06, 
    1.375929e-06, 1.375926e-06, 1.375926e-06, 1.375925e-06, 1.37593e-06, 
    1.375927e-06, 1.375933e-06, 1.375931e-06, 1.375944e-06, 1.375948e-06, 
    1.37595e-06, 1.375952e-06, 1.375957e-06, 1.375954e-06, 1.375955e-06, 
    1.375952e-06, 1.37595e-06, 1.375951e-06, 1.375946e-06, 1.375948e-06, 
    1.375937e-06, 1.375941e-06, 1.375929e-06, 1.375932e-06, 1.375928e-06, 
    1.37593e-06, 1.375927e-06, 1.37593e-06, 1.375925e-06, 1.375923e-06, 
    1.375924e-06, 1.375921e-06, 1.37593e-06, 1.375927e-06, 1.375951e-06, 
    1.375951e-06, 1.37595e-06, 1.375953e-06, 1.375953e-06, 1.375956e-06, 
    1.375954e-06, 1.375953e-06, 1.37595e-06, 1.375949e-06, 1.375947e-06, 
    1.375944e-06, 1.37594e-06, 1.375935e-06, 1.375932e-06, 1.375929e-06, 
    1.375931e-06, 1.375929e-06, 1.375931e-06, 1.375932e-06, 1.375924e-06, 
    1.375928e-06, 1.375922e-06, 1.375922e-06, 1.375925e-06, 1.375922e-06, 
    1.375951e-06, 1.375952e-06, 1.375955e-06, 1.375952e-06, 1.375956e-06, 
    1.375954e-06, 1.375953e-06, 1.375948e-06, 1.375946e-06, 1.375945e-06, 
    1.375943e-06, 1.375941e-06, 1.375936e-06, 1.375932e-06, 1.375928e-06, 
    1.375929e-06, 1.375929e-06, 1.375928e-06, 1.37593e-06, 1.375928e-06, 
    1.375927e-06, 1.375928e-06, 1.375922e-06, 1.375924e-06, 1.375922e-06, 
    1.375923e-06, 1.375951e-06, 1.37595e-06, 1.375951e-06, 1.375949e-06, 
    1.37595e-06, 1.375946e-06, 1.375945e-06, 1.375938e-06, 1.375941e-06, 
    1.375937e-06, 1.37594e-06, 1.37594e-06, 1.375937e-06, 1.37594e-06, 
    1.375932e-06, 1.375938e-06, 1.375928e-06, 1.375933e-06, 1.375928e-06, 
    1.375929e-06, 1.375927e-06, 1.375925e-06, 1.375923e-06, 1.37592e-06, 
    1.375921e-06, 1.375918e-06, 1.375948e-06, 1.375946e-06, 1.375946e-06, 
    1.375944e-06, 1.375943e-06, 1.37594e-06, 1.375935e-06, 1.375937e-06, 
    1.375933e-06, 1.375933e-06, 1.375938e-06, 1.375935e-06, 1.375945e-06, 
    1.375943e-06, 1.375944e-06, 1.375948e-06, 1.375936e-06, 1.375942e-06, 
    1.375932e-06, 1.375935e-06, 1.375926e-06, 1.37593e-06, 1.375921e-06, 
    1.375917e-06, 1.375914e-06, 1.37591e-06, 1.375945e-06, 1.375946e-06, 
    1.375944e-06, 1.375941e-06, 1.375938e-06, 1.375935e-06, 1.375934e-06, 
    1.375933e-06, 1.375932e-06, 1.37593e-06, 1.375933e-06, 1.37593e-06, 
    1.375943e-06, 1.375936e-06, 1.375947e-06, 1.375943e-06, 1.375941e-06, 
    1.375942e-06, 1.375937e-06, 1.375936e-06, 1.375931e-06, 1.375933e-06, 
    1.375918e-06, 1.375925e-06, 1.375906e-06, 1.375912e-06, 1.375947e-06, 
    1.375945e-06, 1.375939e-06, 1.375942e-06, 1.375934e-06, 1.375932e-06, 
    1.375931e-06, 1.375929e-06, 1.375929e-06, 1.375927e-06, 1.375929e-06, 
    1.375927e-06, 1.375935e-06, 1.375931e-06, 1.37594e-06, 1.375938e-06, 
    1.375939e-06, 1.37594e-06, 1.375937e-06, 1.375933e-06, 1.375933e-06, 
    1.375932e-06, 1.375929e-06, 1.375934e-06, 1.375917e-06, 1.375928e-06, 
    1.375943e-06, 1.37594e-06, 1.37594e-06, 1.375941e-06, 1.375932e-06, 
    1.375936e-06, 1.375927e-06, 1.37593e-06, 1.375926e-06, 1.375928e-06, 
    1.375928e-06, 1.37593e-06, 1.375932e-06, 1.375935e-06, 1.375938e-06, 
    1.375941e-06, 1.37594e-06, 1.375938e-06, 1.375933e-06, 1.375928e-06, 
    1.37593e-06, 1.375926e-06, 1.375935e-06, 1.375931e-06, 1.375933e-06, 
    1.375929e-06, 1.375937e-06, 1.37593e-06, 1.375939e-06, 1.375938e-06, 
    1.375936e-06, 1.375931e-06, 1.37593e-06, 1.375929e-06, 1.37593e-06, 
    1.375933e-06, 1.375933e-06, 1.375936e-06, 1.375936e-06, 1.375938e-06, 
    1.37594e-06, 1.375938e-06, 1.375937e-06, 1.375933e-06, 1.375929e-06, 
    1.375925e-06, 1.375924e-06, 1.37592e-06, 1.375923e-06, 1.375917e-06, 
    1.375923e-06, 1.375914e-06, 1.37593e-06, 1.375923e-06, 1.375936e-06, 
    1.375934e-06, 1.375932e-06, 1.375926e-06, 1.375929e-06, 1.375925e-06, 
    1.375933e-06, 1.375937e-06, 1.375939e-06, 1.375941e-06, 1.375938e-06, 
    1.375939e-06, 1.375937e-06, 1.375937e-06, 1.375933e-06, 1.375935e-06, 
    1.375928e-06, 1.375925e-06, 1.375918e-06, 1.375914e-06, 1.375909e-06, 
    1.375907e-06, 1.375906e-06, 1.375906e-06 ;

 TOTPFTC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTPFTN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TOTPRODC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTPRODN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 TOTSOMC =
  17.34481, 17.3448, 17.3448, 17.34479, 17.34479, 17.34479, 17.34481, 
    17.3448, 17.3448, 17.34481, 17.34477, 17.34479, 17.34475, 17.34476, 
    17.34473, 17.34475, 17.34472, 17.34473, 17.34471, 17.34472, 17.3447, 
    17.34471, 17.34469, 17.3447, 17.3447, 17.34471, 17.34478, 17.34477, 
    17.34478, 17.34478, 17.34478, 17.34479, 17.3448, 17.34481, 17.34481, 
    17.3448, 17.34478, 17.34479, 17.34477, 17.34477, 17.34476, 17.34476, 
    17.34473, 17.34474, 17.34472, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34473, 17.34472, 17.34473, 17.34476, 17.34475, 17.34478, 17.3448, 
    17.34481, 17.34481, 17.34481, 17.34481, 17.3448, 17.34479, 17.34478, 
    17.34478, 17.34477, 17.34476, 17.34475, 17.34473, 17.34473, 17.34473, 
    17.34472, 17.34472, 17.34472, 17.34471, 17.34473, 17.34472, 17.34474, 
    17.34473, 17.34477, 17.34479, 17.34479, 17.3448, 17.34481, 17.3448, 
    17.34481, 17.3448, 17.34479, 17.3448, 17.34478, 17.34478, 17.34475, 
    17.34476, 17.34472, 17.34473, 17.34472, 17.34473, 17.34472, 17.34473, 
    17.34471, 17.34471, 17.34471, 17.3447, 17.34473, 17.34472, 17.3448, 
    17.34479, 17.34479, 17.3448, 17.3448, 17.34481, 17.3448, 17.3448, 
    17.34479, 17.34479, 17.34478, 17.34477, 17.34476, 17.34475, 17.34473, 
    17.34473, 17.34473, 17.34473, 17.34473, 17.34473, 17.34471, 17.34472, 
    17.3447, 17.3447, 17.34471, 17.3447, 17.34479, 17.3448, 17.3448, 17.3448, 
    17.34481, 17.3448, 17.3448, 17.34478, 17.34478, 17.34478, 17.34477, 
    17.34476, 17.34475, 17.34474, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34473, 17.34472, 17.34472, 17.34472, 17.3447, 17.34471, 17.3447, 
    17.34471, 17.3448, 17.34479, 17.34479, 17.34479, 17.34479, 17.34478, 
    17.34477, 17.34476, 17.34476, 17.34475, 17.34476, 17.34476, 17.34475, 
    17.34476, 17.34474, 17.34475, 17.34472, 17.34474, 17.34472, 17.34472, 
    17.34472, 17.34471, 17.34471, 17.3447, 17.3447, 17.34469, 17.34478, 
    17.34478, 17.34478, 17.34477, 17.34477, 17.34476, 17.34474, 17.34475, 
    17.34474, 17.34474, 17.34475, 17.34474, 17.34477, 17.34477, 17.34477, 
    17.34478, 17.34475, 17.34477, 17.34473, 17.34474, 17.34472, 17.34473, 
    17.3447, 17.34469, 17.34468, 17.34466, 17.34478, 17.34478, 17.34477, 
    17.34476, 17.34476, 17.34474, 17.34474, 17.34474, 17.34473, 17.34473, 
    17.34474, 17.34473, 17.34477, 17.34475, 17.34478, 17.34477, 17.34476, 
    17.34477, 17.34475, 17.34475, 17.34473, 17.34474, 17.34469, 17.34471, 
    17.34465, 17.34467, 17.34478, 17.34478, 17.34476, 17.34477, 17.34474, 
    17.34474, 17.34473, 17.34472, 17.34472, 17.34472, 17.34473, 17.34472, 
    17.34474, 17.34473, 17.34476, 17.34475, 17.34476, 17.34476, 17.34475, 
    17.34474, 17.34474, 17.34473, 17.34472, 17.34474, 17.34469, 17.34472, 
    17.34477, 17.34476, 17.34476, 17.34476, 17.34474, 17.34475, 17.34472, 
    17.34473, 17.34472, 17.34472, 17.34472, 17.34473, 17.34473, 17.34475, 
    17.34476, 17.34476, 17.34476, 17.34475, 17.34474, 17.34472, 17.34473, 
    17.34472, 17.34474, 17.34473, 17.34474, 17.34472, 17.34475, 17.34473, 
    17.34476, 17.34475, 17.34475, 17.34473, 17.34473, 17.34472, 17.34473, 
    17.34474, 17.34474, 17.34475, 17.34475, 17.34475, 17.34476, 17.34475, 
    17.34475, 17.34474, 17.34473, 17.34471, 17.34471, 17.3447, 17.34471, 
    17.34469, 17.34471, 17.34468, 17.34473, 17.34471, 17.34475, 17.34474, 
    17.34473, 17.34472, 17.34472, 17.34471, 17.34474, 17.34475, 17.34476, 
    17.34476, 17.34476, 17.34476, 17.34475, 17.34475, 17.34474, 17.34475, 
    17.34472, 17.34471, 17.34469, 17.34468, 17.34466, 17.34466, 17.34465, 
    17.34465 ;

 TOTSOMC_1m =
  17.34481, 17.3448, 17.3448, 17.34479, 17.34479, 17.34479, 17.34481, 
    17.3448, 17.3448, 17.34481, 17.34477, 17.34479, 17.34475, 17.34476, 
    17.34473, 17.34475, 17.34472, 17.34473, 17.34471, 17.34472, 17.3447, 
    17.34471, 17.34469, 17.3447, 17.3447, 17.34471, 17.34478, 17.34477, 
    17.34478, 17.34478, 17.34478, 17.34479, 17.3448, 17.34481, 17.34481, 
    17.3448, 17.34478, 17.34479, 17.34477, 17.34477, 17.34476, 17.34476, 
    17.34473, 17.34474, 17.34472, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34473, 17.34472, 17.34473, 17.34476, 17.34475, 17.34478, 17.3448, 
    17.34481, 17.34481, 17.34481, 17.34481, 17.3448, 17.34479, 17.34478, 
    17.34478, 17.34477, 17.34476, 17.34475, 17.34473, 17.34473, 17.34473, 
    17.34472, 17.34472, 17.34472, 17.34471, 17.34473, 17.34472, 17.34474, 
    17.34473, 17.34477, 17.34479, 17.34479, 17.3448, 17.34481, 17.3448, 
    17.34481, 17.3448, 17.34479, 17.3448, 17.34478, 17.34478, 17.34475, 
    17.34476, 17.34472, 17.34473, 17.34472, 17.34473, 17.34472, 17.34473, 
    17.34471, 17.34471, 17.34471, 17.3447, 17.34473, 17.34472, 17.3448, 
    17.34479, 17.34479, 17.3448, 17.3448, 17.34481, 17.3448, 17.3448, 
    17.34479, 17.34479, 17.34478, 17.34477, 17.34476, 17.34475, 17.34473, 
    17.34473, 17.34473, 17.34473, 17.34473, 17.34473, 17.34471, 17.34472, 
    17.3447, 17.3447, 17.34471, 17.3447, 17.34479, 17.3448, 17.3448, 17.3448, 
    17.34481, 17.3448, 17.3448, 17.34478, 17.34478, 17.34478, 17.34477, 
    17.34476, 17.34475, 17.34474, 17.34472, 17.34472, 17.34472, 17.34472, 
    17.34473, 17.34472, 17.34472, 17.34472, 17.3447, 17.34471, 17.3447, 
    17.34471, 17.3448, 17.34479, 17.34479, 17.34479, 17.34479, 17.34478, 
    17.34477, 17.34476, 17.34476, 17.34475, 17.34476, 17.34476, 17.34475, 
    17.34476, 17.34474, 17.34475, 17.34472, 17.34474, 17.34472, 17.34472, 
    17.34472, 17.34471, 17.34471, 17.3447, 17.3447, 17.34469, 17.34478, 
    17.34478, 17.34478, 17.34477, 17.34477, 17.34476, 17.34474, 17.34475, 
    17.34474, 17.34474, 17.34475, 17.34474, 17.34477, 17.34477, 17.34477, 
    17.34478, 17.34475, 17.34477, 17.34473, 17.34474, 17.34472, 17.34473, 
    17.3447, 17.34469, 17.34468, 17.34466, 17.34478, 17.34478, 17.34477, 
    17.34476, 17.34476, 17.34474, 17.34474, 17.34474, 17.34473, 17.34473, 
    17.34474, 17.34473, 17.34477, 17.34475, 17.34478, 17.34477, 17.34476, 
    17.34477, 17.34475, 17.34475, 17.34473, 17.34474, 17.34469, 17.34471, 
    17.34465, 17.34467, 17.34478, 17.34478, 17.34476, 17.34477, 17.34474, 
    17.34474, 17.34473, 17.34472, 17.34472, 17.34472, 17.34473, 17.34472, 
    17.34474, 17.34473, 17.34476, 17.34475, 17.34476, 17.34476, 17.34475, 
    17.34474, 17.34474, 17.34473, 17.34472, 17.34474, 17.34469, 17.34472, 
    17.34477, 17.34476, 17.34476, 17.34476, 17.34474, 17.34475, 17.34472, 
    17.34473, 17.34472, 17.34472, 17.34472, 17.34473, 17.34473, 17.34475, 
    17.34476, 17.34476, 17.34476, 17.34475, 17.34474, 17.34472, 17.34473, 
    17.34472, 17.34474, 17.34473, 17.34474, 17.34472, 17.34475, 17.34473, 
    17.34476, 17.34475, 17.34475, 17.34473, 17.34473, 17.34472, 17.34473, 
    17.34474, 17.34474, 17.34475, 17.34475, 17.34475, 17.34476, 17.34475, 
    17.34475, 17.34474, 17.34473, 17.34471, 17.34471, 17.3447, 17.34471, 
    17.34469, 17.34471, 17.34468, 17.34473, 17.34471, 17.34475, 17.34474, 
    17.34473, 17.34472, 17.34472, 17.34471, 17.34474, 17.34475, 17.34476, 
    17.34476, 17.34476, 17.34476, 17.34475, 17.34475, 17.34474, 17.34475, 
    17.34472, 17.34471, 17.34469, 17.34468, 17.34466, 17.34466, 17.34465, 
    17.34465 ;

 TOTSOMN =
  1.773786, 1.773785, 1.773785, 1.773783, 1.773784, 1.773783, 1.773786, 
    1.773785, 1.773785, 1.773786, 1.773781, 1.773783, 1.773778, 1.773779, 
    1.773775, 1.773778, 1.773774, 1.773775, 1.773773, 1.773773, 1.773771, 
    1.773773, 1.773769, 1.773771, 1.773771, 1.773773, 1.773783, 1.773781, 
    1.773783, 1.773783, 1.773783, 1.773784, 1.773785, 1.773787, 1.773786, 
    1.773785, 1.773782, 1.773783, 1.773781, 1.773781, 1.773779, 1.77378, 
    1.773776, 1.773777, 1.773773, 1.773774, 1.773774, 1.773774, 1.773774, 
    1.773775, 1.773774, 1.773775, 1.77378, 1.773778, 1.773782, 1.773784, 
    1.773786, 1.773787, 1.773787, 1.773787, 1.773785, 1.773784, 1.773783, 
    1.773782, 1.773781, 1.773779, 1.773778, 1.773775, 1.773776, 1.773775, 
    1.773774, 1.773773, 1.773773, 1.773773, 1.773775, 1.773774, 1.773776, 
    1.773775, 1.773781, 1.773783, 1.773784, 1.773785, 1.773787, 1.773785, 
    1.773786, 1.773785, 1.773784, 1.773784, 1.773782, 1.773783, 1.773778, 
    1.77378, 1.773775, 1.773776, 1.773774, 1.773775, 1.773774, 1.773775, 
    1.773773, 1.773772, 1.773772, 1.773771, 1.773775, 1.773774, 1.773784, 
    1.773784, 1.773784, 1.773785, 1.773785, 1.773787, 1.773785, 1.773785, 
    1.773784, 1.773783, 1.773782, 1.773781, 1.77378, 1.773777, 1.773776, 
    1.773775, 1.773775, 1.773775, 1.773775, 1.773776, 1.773772, 1.773774, 
    1.773771, 1.773772, 1.773773, 1.773772, 1.773784, 1.773785, 1.773786, 
    1.773785, 1.773787, 1.773786, 1.773785, 1.773783, 1.773782, 1.773782, 
    1.773781, 1.77378, 1.773778, 1.773776, 1.773774, 1.773775, 1.773774, 
    1.773774, 1.773775, 1.773774, 1.773774, 1.773774, 1.773772, 1.773772, 
    1.773772, 1.773772, 1.773785, 1.773784, 1.773784, 1.773784, 1.773784, 
    1.773782, 1.773781, 1.773779, 1.77378, 1.773778, 1.77378, 1.773779, 
    1.773778, 1.77378, 1.773776, 1.773778, 1.773774, 1.773776, 1.773774, 
    1.773774, 1.773774, 1.773773, 1.773772, 1.773771, 1.773771, 1.77377, 
    1.773783, 1.773782, 1.773782, 1.773781, 1.773781, 1.773779, 1.773777, 
    1.773778, 1.773777, 1.773776, 1.773779, 1.773777, 1.773782, 1.773781, 
    1.773781, 1.773783, 1.773778, 1.77378, 1.773776, 1.773777, 1.773773, 
    1.773775, 1.773771, 1.773769, 1.773768, 1.773766, 1.773782, 1.773782, 
    1.773781, 1.77378, 1.773779, 1.773777, 1.773777, 1.773777, 1.773776, 
    1.773775, 1.773776, 1.773775, 1.773781, 1.773778, 1.773782, 1.773781, 
    1.77378, 1.77378, 1.773778, 1.773778, 1.773775, 1.773777, 1.77377, 
    1.773773, 1.773764, 1.773767, 1.773782, 1.773782, 1.773779, 1.77378, 
    1.773777, 1.773776, 1.773775, 1.773775, 1.773774, 1.773774, 1.773775, 
    1.773774, 1.773777, 1.773776, 1.773779, 1.773779, 1.773779, 1.773779, 
    1.773778, 1.773776, 1.773776, 1.773776, 1.773775, 1.773777, 1.773769, 
    1.773774, 1.773781, 1.77378, 1.773779, 1.77378, 1.773776, 1.773777, 
    1.773774, 1.773775, 1.773773, 1.773774, 1.773774, 1.773775, 1.773776, 
    1.773777, 1.773779, 1.77378, 1.77378, 1.773778, 1.773776, 1.773774, 
    1.773775, 1.773773, 1.773777, 1.773776, 1.773776, 1.773775, 1.773778, 
    1.773775, 1.773779, 1.773779, 1.773777, 1.773775, 1.773775, 1.773775, 
    1.773775, 1.773776, 1.773777, 1.773777, 1.773778, 1.773779, 1.773779, 
    1.773779, 1.773778, 1.773776, 1.773775, 1.773773, 1.773772, 1.77377, 
    1.773772, 1.773769, 1.773772, 1.773768, 1.773775, 1.773772, 1.773777, 
    1.773777, 1.773776, 1.773773, 1.773775, 1.773773, 1.773777, 1.773778, 
    1.773779, 1.77378, 1.773779, 1.773779, 1.773778, 1.773778, 1.773776, 
    1.773777, 1.773774, 1.773773, 1.77377, 1.773768, 1.773766, 1.773765, 
    1.773764, 1.773764 ;

 TOTSOMN_1m =
  1.773786, 1.773785, 1.773785, 1.773783, 1.773784, 1.773783, 1.773786, 
    1.773785, 1.773785, 1.773786, 1.773781, 1.773783, 1.773778, 1.773779, 
    1.773775, 1.773778, 1.773774, 1.773775, 1.773773, 1.773773, 1.773771, 
    1.773773, 1.773769, 1.773771, 1.773771, 1.773773, 1.773783, 1.773781, 
    1.773783, 1.773783, 1.773783, 1.773784, 1.773785, 1.773787, 1.773786, 
    1.773785, 1.773782, 1.773783, 1.773781, 1.773781, 1.773779, 1.77378, 
    1.773776, 1.773777, 1.773773, 1.773774, 1.773774, 1.773774, 1.773774, 
    1.773775, 1.773774, 1.773775, 1.77378, 1.773778, 1.773782, 1.773784, 
    1.773786, 1.773787, 1.773787, 1.773787, 1.773785, 1.773784, 1.773783, 
    1.773782, 1.773781, 1.773779, 1.773778, 1.773775, 1.773776, 1.773775, 
    1.773774, 1.773773, 1.773773, 1.773773, 1.773775, 1.773774, 1.773776, 
    1.773775, 1.773781, 1.773783, 1.773784, 1.773785, 1.773787, 1.773785, 
    1.773786, 1.773785, 1.773784, 1.773784, 1.773782, 1.773783, 1.773778, 
    1.77378, 1.773775, 1.773776, 1.773774, 1.773775, 1.773774, 1.773775, 
    1.773773, 1.773772, 1.773772, 1.773771, 1.773775, 1.773774, 1.773784, 
    1.773784, 1.773784, 1.773785, 1.773785, 1.773787, 1.773785, 1.773785, 
    1.773784, 1.773783, 1.773782, 1.773781, 1.77378, 1.773777, 1.773776, 
    1.773775, 1.773775, 1.773775, 1.773775, 1.773776, 1.773772, 1.773774, 
    1.773771, 1.773772, 1.773773, 1.773772, 1.773784, 1.773785, 1.773786, 
    1.773785, 1.773787, 1.773786, 1.773785, 1.773783, 1.773782, 1.773782, 
    1.773781, 1.77378, 1.773778, 1.773776, 1.773774, 1.773775, 1.773774, 
    1.773774, 1.773775, 1.773774, 1.773774, 1.773774, 1.773772, 1.773772, 
    1.773772, 1.773772, 1.773785, 1.773784, 1.773784, 1.773784, 1.773784, 
    1.773782, 1.773781, 1.773779, 1.77378, 1.773778, 1.77378, 1.773779, 
    1.773778, 1.77378, 1.773776, 1.773778, 1.773774, 1.773776, 1.773774, 
    1.773774, 1.773774, 1.773773, 1.773772, 1.773771, 1.773771, 1.77377, 
    1.773783, 1.773782, 1.773782, 1.773781, 1.773781, 1.773779, 1.773777, 
    1.773778, 1.773777, 1.773776, 1.773779, 1.773777, 1.773782, 1.773781, 
    1.773781, 1.773783, 1.773778, 1.77378, 1.773776, 1.773777, 1.773773, 
    1.773775, 1.773771, 1.773769, 1.773768, 1.773766, 1.773782, 1.773782, 
    1.773781, 1.77378, 1.773779, 1.773777, 1.773777, 1.773777, 1.773776, 
    1.773775, 1.773776, 1.773775, 1.773781, 1.773778, 1.773782, 1.773781, 
    1.77378, 1.77378, 1.773778, 1.773778, 1.773775, 1.773777, 1.77377, 
    1.773773, 1.773764, 1.773767, 1.773782, 1.773782, 1.773779, 1.77378, 
    1.773777, 1.773776, 1.773775, 1.773775, 1.773774, 1.773774, 1.773775, 
    1.773774, 1.773777, 1.773776, 1.773779, 1.773779, 1.773779, 1.773779, 
    1.773778, 1.773776, 1.773776, 1.773776, 1.773775, 1.773777, 1.773769, 
    1.773774, 1.773781, 1.77378, 1.773779, 1.77378, 1.773776, 1.773777, 
    1.773774, 1.773775, 1.773773, 1.773774, 1.773774, 1.773775, 1.773776, 
    1.773777, 1.773779, 1.77378, 1.77378, 1.773778, 1.773776, 1.773774, 
    1.773775, 1.773773, 1.773777, 1.773776, 1.773776, 1.773775, 1.773778, 
    1.773775, 1.773779, 1.773779, 1.773777, 1.773775, 1.773775, 1.773775, 
    1.773775, 1.773776, 1.773777, 1.773777, 1.773778, 1.773779, 1.773779, 
    1.773779, 1.773778, 1.773776, 1.773775, 1.773773, 1.773772, 1.77377, 
    1.773772, 1.773769, 1.773772, 1.773768, 1.773775, 1.773772, 1.773777, 
    1.773777, 1.773776, 1.773773, 1.773775, 1.773773, 1.773777, 1.773778, 
    1.773779, 1.77378, 1.773779, 1.773779, 1.773778, 1.773778, 1.773776, 
    1.773777, 1.773774, 1.773773, 1.77377, 1.773768, 1.773766, 1.773765, 
    1.773764, 1.773764 ;

 TOTVEGC =
  0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 0.8953198, 
    0.8953198, 0.8953198 ;

 TOTVEGN =
  0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 0.03250261, 
    0.03250261, 0.03250261 ;

 TREFMNAV =
  249.9695, 249.9697, 249.9697, 249.9699, 249.9698, 249.9699, 249.9695, 
    249.9697, 249.9696, 249.9695, 249.9703, 249.9699, 249.9707, 249.9704, 
    249.9711, 249.9706, 249.9711, 249.9711, 249.9714, 249.9713, 249.9716, 
    249.9714, 249.9718, 249.9716, 249.9716, 249.9714, 249.97, 249.9702, 
    249.9699, 249.97, 249.97, 249.9698, 249.9697, 249.9694, 249.9695, 
    249.9696, 249.97, 249.9699, 249.9702, 249.9702, 249.9705, 249.9704, 
    249.9709, 249.9708, 249.9713, 249.9711, 249.9713, 249.9712, 249.9713, 
    249.9711, 249.9712, 249.971, 249.9704, 249.9706, 249.97, 249.9697, 
    249.9695, 249.9694, 249.9694, 249.9694, 249.9696, 249.9698, 249.97, 
    249.9701, 249.9702, 249.9705, 249.9706, 249.971, 249.9709, 249.971, 
    249.9711, 249.9713, 249.9713, 249.9714, 249.971, 249.9713, 249.9709, 
    249.971, 249.9702, 249.9699, 249.9698, 249.9697, 249.9694, 249.9696, 
    249.9695, 249.9697, 249.9698, 249.9697, 249.9701, 249.97, 249.9706, 
    249.9703, 249.9711, 249.9709, 249.9712, 249.9711, 249.9713, 249.9711, 
    249.9714, 249.9715, 249.9714, 249.9716, 249.9711, 249.9713, 249.9697, 
    249.9698, 249.9698, 249.9696, 249.9696, 249.9694, 249.9696, 249.9696, 
    249.9698, 249.9699, 249.97, 249.9702, 249.9704, 249.9707, 249.9709, 
    249.9711, 249.971, 249.9711, 249.971, 249.971, 249.9714, 249.9712, 
    249.9716, 249.9715, 249.9714, 249.9715, 249.9698, 249.9697, 249.9695, 
    249.9697, 249.9694, 249.9696, 249.9696, 249.97, 249.97, 249.9701, 
    249.9702, 249.9704, 249.9707, 249.9709, 249.9711, 249.9711, 249.9711, 
    249.9712, 249.9711, 249.9712, 249.9712, 249.9712, 249.9715, 249.9714, 
    249.9715, 249.9715, 249.9697, 249.9698, 249.9698, 249.9698, 249.9698, 
    249.9701, 249.9701, 249.9705, 249.9704, 249.9706, 249.9704, 249.9704, 
    249.9706, 249.9704, 249.9709, 249.9706, 249.9712, 249.9708, 249.9712, 
    249.9711, 249.9713, 249.9713, 249.9715, 249.9717, 249.9716, 249.9718, 
    249.9699, 249.97, 249.97, 249.9702, 249.9702, 249.9704, 249.9707, 
    249.9706, 249.9708, 249.9709, 249.9706, 249.9707, 249.9701, 249.9702, 
    249.9702, 249.9699, 249.9706, 249.9703, 249.9709, 249.9708, 249.9713, 
    249.971, 249.9716, 249.9718, 249.9721, 249.9723, 249.9701, 249.97, 
    249.9702, 249.9704, 249.9705, 249.9708, 249.9708, 249.9708, 249.9709, 
    249.9711, 249.9708, 249.9711, 249.9702, 249.9707, 249.97, 249.9702, 
    249.9704, 249.9703, 249.9706, 249.9707, 249.971, 249.9708, 249.9718, 
    249.9714, 249.9725, 249.9722, 249.97, 249.9701, 249.9705, 249.9703, 
    249.9708, 249.9709, 249.971, 249.9711, 249.9711, 249.9712, 249.9711, 
    249.9712, 249.9708, 249.971, 249.9704, 249.9706, 249.9705, 249.9704, 
    249.9706, 249.9709, 249.9709, 249.9709, 249.9711, 249.9708, 249.9718, 
    249.9712, 249.9702, 249.9704, 249.9704, 249.9704, 249.9709, 249.9707, 
    249.9712, 249.9711, 249.9713, 249.9712, 249.9712, 249.971, 249.9709, 
    249.9707, 249.9705, 249.9704, 249.9704, 249.9706, 249.9709, 249.9711, 
    249.9711, 249.9713, 249.9707, 249.971, 249.9709, 249.9711, 249.9706, 
    249.971, 249.9705, 249.9706, 249.9707, 249.971, 249.9711, 249.9711, 
    249.9711, 249.9709, 249.9708, 249.9707, 249.9707, 249.9706, 249.9705, 
    249.9705, 249.9706, 249.9709, 249.9711, 249.9713, 249.9714, 249.9717, 
    249.9715, 249.9718, 249.9715, 249.9721, 249.9711, 249.9715, 249.9707, 
    249.9708, 249.9709, 249.9713, 249.9711, 249.9713, 249.9708, 249.9706, 
    249.9705, 249.9704, 249.9705, 249.9705, 249.9706, 249.9706, 249.9709, 
    249.9707, 249.9712, 249.9713, 249.9718, 249.9721, 249.9724, 249.9725, 
    249.9725, 249.9725 ;

 TREFMNAV_R =
  249.9695, 249.9697, 249.9697, 249.9699, 249.9698, 249.9699, 249.9695, 
    249.9697, 249.9696, 249.9695, 249.9703, 249.9699, 249.9707, 249.9704, 
    249.9711, 249.9706, 249.9711, 249.9711, 249.9714, 249.9713, 249.9716, 
    249.9714, 249.9718, 249.9716, 249.9716, 249.9714, 249.97, 249.9702, 
    249.9699, 249.97, 249.97, 249.9698, 249.9697, 249.9694, 249.9695, 
    249.9696, 249.97, 249.9699, 249.9702, 249.9702, 249.9705, 249.9704, 
    249.9709, 249.9708, 249.9713, 249.9711, 249.9713, 249.9712, 249.9713, 
    249.9711, 249.9712, 249.971, 249.9704, 249.9706, 249.97, 249.9697, 
    249.9695, 249.9694, 249.9694, 249.9694, 249.9696, 249.9698, 249.97, 
    249.9701, 249.9702, 249.9705, 249.9706, 249.971, 249.9709, 249.971, 
    249.9711, 249.9713, 249.9713, 249.9714, 249.971, 249.9713, 249.9709, 
    249.971, 249.9702, 249.9699, 249.9698, 249.9697, 249.9694, 249.9696, 
    249.9695, 249.9697, 249.9698, 249.9697, 249.9701, 249.97, 249.9706, 
    249.9703, 249.9711, 249.9709, 249.9712, 249.9711, 249.9713, 249.9711, 
    249.9714, 249.9715, 249.9714, 249.9716, 249.9711, 249.9713, 249.9697, 
    249.9698, 249.9698, 249.9696, 249.9696, 249.9694, 249.9696, 249.9696, 
    249.9698, 249.9699, 249.97, 249.9702, 249.9704, 249.9707, 249.9709, 
    249.9711, 249.971, 249.9711, 249.971, 249.971, 249.9714, 249.9712, 
    249.9716, 249.9715, 249.9714, 249.9715, 249.9698, 249.9697, 249.9695, 
    249.9697, 249.9694, 249.9696, 249.9696, 249.97, 249.97, 249.9701, 
    249.9702, 249.9704, 249.9707, 249.9709, 249.9711, 249.9711, 249.9711, 
    249.9712, 249.9711, 249.9712, 249.9712, 249.9712, 249.9715, 249.9714, 
    249.9715, 249.9715, 249.9697, 249.9698, 249.9698, 249.9698, 249.9698, 
    249.9701, 249.9701, 249.9705, 249.9704, 249.9706, 249.9704, 249.9704, 
    249.9706, 249.9704, 249.9709, 249.9706, 249.9712, 249.9708, 249.9712, 
    249.9711, 249.9713, 249.9713, 249.9715, 249.9717, 249.9716, 249.9718, 
    249.9699, 249.97, 249.97, 249.9702, 249.9702, 249.9704, 249.9707, 
    249.9706, 249.9708, 249.9709, 249.9706, 249.9707, 249.9701, 249.9702, 
    249.9702, 249.9699, 249.9706, 249.9703, 249.9709, 249.9708, 249.9713, 
    249.971, 249.9716, 249.9718, 249.9721, 249.9723, 249.9701, 249.97, 
    249.9702, 249.9704, 249.9705, 249.9708, 249.9708, 249.9708, 249.9709, 
    249.9711, 249.9708, 249.9711, 249.9702, 249.9707, 249.97, 249.9702, 
    249.9704, 249.9703, 249.9706, 249.9707, 249.971, 249.9708, 249.9718, 
    249.9714, 249.9725, 249.9722, 249.97, 249.9701, 249.9705, 249.9703, 
    249.9708, 249.9709, 249.971, 249.9711, 249.9711, 249.9712, 249.9711, 
    249.9712, 249.9708, 249.971, 249.9704, 249.9706, 249.9705, 249.9704, 
    249.9706, 249.9709, 249.9709, 249.9709, 249.9711, 249.9708, 249.9718, 
    249.9712, 249.9702, 249.9704, 249.9704, 249.9704, 249.9709, 249.9707, 
    249.9712, 249.9711, 249.9713, 249.9712, 249.9712, 249.971, 249.9709, 
    249.9707, 249.9705, 249.9704, 249.9704, 249.9706, 249.9709, 249.9711, 
    249.9711, 249.9713, 249.9707, 249.971, 249.9709, 249.9711, 249.9706, 
    249.971, 249.9705, 249.9706, 249.9707, 249.971, 249.9711, 249.9711, 
    249.9711, 249.9709, 249.9708, 249.9707, 249.9707, 249.9706, 249.9705, 
    249.9705, 249.9706, 249.9709, 249.9711, 249.9713, 249.9714, 249.9717, 
    249.9715, 249.9718, 249.9715, 249.9721, 249.9711, 249.9715, 249.9707, 
    249.9708, 249.9709, 249.9713, 249.9711, 249.9713, 249.9708, 249.9706, 
    249.9705, 249.9704, 249.9705, 249.9705, 249.9706, 249.9706, 249.9709, 
    249.9707, 249.9712, 249.9713, 249.9718, 249.9721, 249.9724, 249.9725, 
    249.9725, 249.9725 ;

 TREFMNAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TREFMXAV =
  258.516, 258.5164, 258.5163, 258.5167, 258.5165, 258.5167, 258.5161, 
    258.5164, 258.5162, 258.5161, 258.5173, 258.5167, 258.5179, 258.5175, 
    258.5185, 258.5179, 258.5187, 258.5185, 258.519, 258.5189, 258.5194, 
    258.519, 258.5197, 258.5193, 258.5194, 258.519, 258.5168, 258.5172, 
    258.5168, 258.5168, 258.5168, 258.5165, 258.5163, 258.516, 258.5161, 
    258.5163, 258.5168, 258.5167, 258.5172, 258.5172, 258.5177, 258.5175, 
    258.5184, 258.5181, 258.5189, 258.5187, 258.5189, 258.5188, 258.5189, 
    258.5186, 258.5187, 258.5184, 258.5175, 258.5178, 258.5169, 258.5164, 
    258.5161, 258.5159, 258.5159, 258.516, 258.5163, 258.5166, 258.5168, 
    258.517, 258.5172, 258.5176, 258.5179, 258.5184, 258.5183, 258.5185, 
    258.5186, 258.5189, 258.5189, 258.519, 258.5185, 258.5188, 258.5182, 
    258.5184, 258.5172, 258.5167, 258.5165, 258.5164, 258.5159, 258.5162, 
    258.5161, 258.5164, 258.5165, 258.5165, 258.517, 258.5168, 258.5179, 
    258.5174, 258.5186, 258.5183, 258.5187, 258.5185, 258.5188, 258.5186, 
    258.519, 258.5191, 258.5191, 258.5193, 258.5185, 258.5189, 258.5165, 
    258.5165, 258.5165, 258.5163, 258.5162, 258.516, 258.5162, 258.5163, 
    258.5166, 258.5167, 258.5168, 258.5172, 258.5175, 258.518, 258.5184, 
    258.5186, 258.5185, 258.5186, 258.5184, 258.5184, 258.5191, 258.5187, 
    258.5193, 258.5193, 258.519, 258.5193, 258.5165, 258.5164, 258.5161, 
    258.5164, 258.516, 258.5162, 258.5163, 258.5168, 258.5169, 258.517, 
    258.5172, 258.5175, 258.5179, 258.5183, 258.5186, 258.5186, 258.5186, 
    258.5187, 258.5185, 258.5188, 258.5188, 258.5187, 258.5193, 258.5191, 
    258.5193, 258.5192, 258.5164, 258.5166, 258.5165, 258.5166, 258.5165, 
    258.517, 258.5171, 258.5177, 258.5175, 258.5179, 258.5175, 258.5175, 
    258.5179, 258.5175, 258.5183, 258.5178, 258.5187, 258.5182, 258.5188, 
    258.5186, 258.5188, 258.519, 258.5192, 258.5195, 258.5194, 258.5197, 
    258.5168, 258.5169, 258.5169, 258.5171, 258.5172, 258.5175, 258.518, 
    258.5179, 258.5182, 258.5182, 258.5177, 258.518, 258.5171, 258.5172, 
    258.5171, 258.5168, 258.5179, 258.5173, 258.5184, 258.5181, 258.519, 
    258.5185, 258.5194, 258.5197, 258.5201, 258.5205, 258.517, 258.5169, 
    258.5172, 258.5174, 258.5177, 258.5181, 258.5181, 258.5182, 258.5184, 
    258.5185, 258.5182, 258.5186, 258.5172, 258.5179, 258.5169, 258.5172, 
    258.5174, 258.5173, 258.5178, 258.5179, 258.5184, 258.5182, 258.5197, 
    258.519, 258.5208, 258.5203, 258.5169, 258.5171, 258.5176, 258.5173, 
    258.5181, 258.5183, 258.5184, 258.5186, 258.5186, 258.5188, 258.5186, 
    258.5188, 258.5181, 258.5184, 258.5175, 258.5177, 258.5176, 258.5175, 
    258.5179, 258.5182, 258.5182, 258.5183, 258.5186, 258.5181, 258.5197, 
    258.5187, 258.5172, 258.5175, 258.5176, 258.5175, 258.5183, 258.518, 
    258.5188, 258.5186, 258.5189, 258.5187, 258.5187, 258.5185, 258.5183, 
    258.518, 258.5177, 258.5175, 258.5175, 258.5178, 258.5182, 258.5186, 
    258.5186, 258.5189, 258.518, 258.5184, 258.5182, 258.5186, 258.5179, 
    258.5185, 258.5177, 258.5177, 258.518, 258.5184, 258.5185, 258.5186, 
    258.5186, 258.5182, 258.5182, 258.518, 258.5179, 258.5177, 258.5176, 
    258.5177, 258.5179, 258.5182, 258.5186, 258.519, 258.5191, 258.5195, 
    258.5191, 258.5197, 258.5192, 258.5201, 258.5185, 258.5192, 258.518, 
    258.5181, 258.5183, 258.5189, 258.5186, 258.519, 258.5182, 258.5178, 
    258.5177, 258.5175, 258.5177, 258.5177, 258.5179, 258.5178, 258.5182, 
    258.518, 258.5187, 258.519, 258.5197, 258.5201, 258.5206, 258.5208, 
    258.5208, 258.5209 ;

 TREFMXAV_R =
  258.516, 258.5164, 258.5163, 258.5167, 258.5165, 258.5167, 258.5161, 
    258.5164, 258.5162, 258.5161, 258.5173, 258.5167, 258.5179, 258.5175, 
    258.5185, 258.5179, 258.5187, 258.5185, 258.519, 258.5189, 258.5194, 
    258.519, 258.5197, 258.5193, 258.5194, 258.519, 258.5168, 258.5172, 
    258.5168, 258.5168, 258.5168, 258.5165, 258.5163, 258.516, 258.5161, 
    258.5163, 258.5168, 258.5167, 258.5172, 258.5172, 258.5177, 258.5175, 
    258.5184, 258.5181, 258.5189, 258.5187, 258.5189, 258.5188, 258.5189, 
    258.5186, 258.5187, 258.5184, 258.5175, 258.5178, 258.5169, 258.5164, 
    258.5161, 258.5159, 258.5159, 258.516, 258.5163, 258.5166, 258.5168, 
    258.517, 258.5172, 258.5176, 258.5179, 258.5184, 258.5183, 258.5185, 
    258.5186, 258.5189, 258.5189, 258.519, 258.5185, 258.5188, 258.5182, 
    258.5184, 258.5172, 258.5167, 258.5165, 258.5164, 258.5159, 258.5162, 
    258.5161, 258.5164, 258.5165, 258.5165, 258.517, 258.5168, 258.5179, 
    258.5174, 258.5186, 258.5183, 258.5187, 258.5185, 258.5188, 258.5186, 
    258.519, 258.5191, 258.5191, 258.5193, 258.5185, 258.5189, 258.5165, 
    258.5165, 258.5165, 258.5163, 258.5162, 258.516, 258.5162, 258.5163, 
    258.5166, 258.5167, 258.5168, 258.5172, 258.5175, 258.518, 258.5184, 
    258.5186, 258.5185, 258.5186, 258.5184, 258.5184, 258.5191, 258.5187, 
    258.5193, 258.5193, 258.519, 258.5193, 258.5165, 258.5164, 258.5161, 
    258.5164, 258.516, 258.5162, 258.5163, 258.5168, 258.5169, 258.517, 
    258.5172, 258.5175, 258.5179, 258.5183, 258.5186, 258.5186, 258.5186, 
    258.5187, 258.5185, 258.5188, 258.5188, 258.5187, 258.5193, 258.5191, 
    258.5193, 258.5192, 258.5164, 258.5166, 258.5165, 258.5166, 258.5165, 
    258.517, 258.5171, 258.5177, 258.5175, 258.5179, 258.5175, 258.5175, 
    258.5179, 258.5175, 258.5183, 258.5178, 258.5187, 258.5182, 258.5188, 
    258.5186, 258.5188, 258.519, 258.5192, 258.5195, 258.5194, 258.5197, 
    258.5168, 258.5169, 258.5169, 258.5171, 258.5172, 258.5175, 258.518, 
    258.5179, 258.5182, 258.5182, 258.5177, 258.518, 258.5171, 258.5172, 
    258.5171, 258.5168, 258.5179, 258.5173, 258.5184, 258.5181, 258.519, 
    258.5185, 258.5194, 258.5197, 258.5201, 258.5205, 258.517, 258.5169, 
    258.5172, 258.5174, 258.5177, 258.5181, 258.5181, 258.5182, 258.5184, 
    258.5185, 258.5182, 258.5186, 258.5172, 258.5179, 258.5169, 258.5172, 
    258.5174, 258.5173, 258.5178, 258.5179, 258.5184, 258.5182, 258.5197, 
    258.519, 258.5208, 258.5203, 258.5169, 258.5171, 258.5176, 258.5173, 
    258.5181, 258.5183, 258.5184, 258.5186, 258.5186, 258.5188, 258.5186, 
    258.5188, 258.5181, 258.5184, 258.5175, 258.5177, 258.5176, 258.5175, 
    258.5179, 258.5182, 258.5182, 258.5183, 258.5186, 258.5181, 258.5197, 
    258.5187, 258.5172, 258.5175, 258.5176, 258.5175, 258.5183, 258.518, 
    258.5188, 258.5186, 258.5189, 258.5187, 258.5187, 258.5185, 258.5183, 
    258.518, 258.5177, 258.5175, 258.5175, 258.5178, 258.5182, 258.5186, 
    258.5186, 258.5189, 258.518, 258.5184, 258.5182, 258.5186, 258.5179, 
    258.5185, 258.5177, 258.5177, 258.518, 258.5184, 258.5185, 258.5186, 
    258.5186, 258.5182, 258.5182, 258.518, 258.5179, 258.5177, 258.5176, 
    258.5177, 258.5179, 258.5182, 258.5186, 258.519, 258.5191, 258.5195, 
    258.5191, 258.5197, 258.5192, 258.5201, 258.5185, 258.5192, 258.518, 
    258.5181, 258.5183, 258.5189, 258.5186, 258.519, 258.5182, 258.5178, 
    258.5177, 258.5175, 258.5177, 258.5177, 258.5179, 258.5178, 258.5182, 
    258.518, 258.5187, 258.519, 258.5197, 258.5201, 258.5206, 258.5208, 
    258.5208, 258.5209 ;

 TREFMXAV_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSA =
  253.9562, 253.9564, 253.9563, 253.9565, 253.9564, 253.9565, 253.9562, 
    253.9564, 253.9563, 253.9562, 253.9567, 253.9565, 253.957, 253.9568, 
    253.9573, 253.957, 253.9573, 253.9573, 253.9575, 253.9574, 253.9577, 
    253.9575, 253.9578, 253.9576, 253.9577, 253.9575, 253.9565, 253.9567, 
    253.9565, 253.9565, 253.9565, 253.9564, 253.9563, 253.9562, 253.9562, 
    253.9563, 253.9566, 253.9565, 253.9567, 253.9567, 253.9569, 253.9568, 
    253.9572, 253.9571, 253.9574, 253.9573, 253.9574, 253.9574, 253.9574, 
    253.9573, 253.9574, 253.9572, 253.9568, 253.957, 253.9566, 253.9564, 
    253.9562, 253.9561, 253.9561, 253.9562, 253.9563, 253.9565, 253.9566, 
    253.9566, 253.9567, 253.9569, 253.957, 253.9572, 253.9572, 253.9573, 
    253.9573, 253.9574, 253.9574, 253.9575, 253.9573, 253.9574, 253.9572, 
    253.9572, 253.9567, 253.9565, 253.9564, 253.9563, 253.9562, 253.9563, 
    253.9562, 253.9564, 253.9564, 253.9564, 253.9566, 253.9565, 253.957, 
    253.9568, 253.9573, 253.9572, 253.9574, 253.9573, 253.9574, 253.9573, 
    253.9575, 253.9576, 253.9575, 253.9576, 253.9573, 253.9574, 253.9564, 
    253.9564, 253.9564, 253.9563, 253.9563, 253.9562, 253.9563, 253.9563, 
    253.9564, 253.9565, 253.9566, 253.9567, 253.9568, 253.957, 253.9572, 
    253.9573, 253.9572, 253.9573, 253.9572, 253.9572, 253.9575, 253.9574, 
    253.9576, 253.9576, 253.9575, 253.9576, 253.9564, 253.9564, 253.9563, 
    253.9563, 253.9562, 253.9563, 253.9563, 253.9565, 253.9566, 253.9566, 
    253.9567, 253.9568, 253.957, 253.9572, 253.9573, 253.9573, 253.9573, 
    253.9574, 253.9573, 253.9574, 253.9574, 253.9574, 253.9576, 253.9575, 
    253.9576, 253.9576, 253.9564, 253.9564, 253.9564, 253.9565, 253.9564, 
    253.9566, 253.9567, 253.9569, 253.9568, 253.957, 253.9568, 253.9569, 
    253.957, 253.9568, 253.9572, 253.9569, 253.9574, 253.9571, 253.9574, 
    253.9573, 253.9574, 253.9575, 253.9576, 253.9577, 253.9577, 253.9578, 
    253.9565, 253.9566, 253.9566, 253.9567, 253.9567, 253.9569, 253.9571, 
    253.957, 253.9571, 253.9572, 253.9569, 253.9571, 253.9566, 253.9567, 
    253.9567, 253.9565, 253.957, 253.9568, 253.9572, 253.9571, 253.9575, 
    253.9573, 253.9576, 253.9578, 253.958, 253.9581, 253.9566, 253.9566, 
    253.9567, 253.9568, 253.9569, 253.9571, 253.9571, 253.9571, 253.9572, 
    253.9573, 253.9571, 253.9573, 253.9567, 253.957, 253.9566, 253.9567, 
    253.9568, 253.9568, 253.957, 253.957, 253.9572, 253.9571, 253.9578, 
    253.9575, 253.9583, 253.958, 253.9566, 253.9566, 253.9569, 253.9568, 
    253.9571, 253.9572, 253.9572, 253.9573, 253.9573, 253.9574, 253.9573, 
    253.9574, 253.9571, 253.9572, 253.9568, 253.9569, 253.9569, 253.9569, 
    253.957, 253.9571, 253.9571, 253.9572, 253.9573, 253.9571, 253.9578, 
    253.9574, 253.9567, 253.9568, 253.9569, 253.9568, 253.9572, 253.957, 
    253.9574, 253.9573, 253.9574, 253.9574, 253.9574, 253.9573, 253.9572, 
    253.957, 253.9569, 253.9568, 253.9568, 253.957, 253.9572, 253.9573, 
    253.9573, 253.9574, 253.9571, 253.9572, 253.9572, 253.9573, 253.957, 
    253.9573, 253.9569, 253.9569, 253.957, 253.9572, 253.9573, 253.9573, 
    253.9573, 253.9572, 253.9571, 253.957, 253.957, 253.9569, 253.9569, 
    253.9569, 253.957, 253.9572, 253.9573, 253.9575, 253.9575, 253.9577, 
    253.9575, 253.9578, 253.9576, 253.958, 253.9573, 253.9576, 253.957, 
    253.9571, 253.9572, 253.9574, 253.9573, 253.9575, 253.9571, 253.957, 
    253.9569, 253.9568, 253.9569, 253.9569, 253.957, 253.957, 253.9572, 
    253.9571, 253.9574, 253.9575, 253.9578, 253.958, 253.9582, 253.9583, 
    253.9583, 253.9583 ;

 TSAI =
  0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 0.4233107, 
    0.4233107, 0.4233107 ;

 TSA_R =
  253.9562, 253.9564, 253.9563, 253.9565, 253.9564, 253.9565, 253.9562, 
    253.9564, 253.9563, 253.9562, 253.9567, 253.9565, 253.957, 253.9568, 
    253.9573, 253.957, 253.9573, 253.9573, 253.9575, 253.9574, 253.9577, 
    253.9575, 253.9578, 253.9576, 253.9577, 253.9575, 253.9565, 253.9567, 
    253.9565, 253.9565, 253.9565, 253.9564, 253.9563, 253.9562, 253.9562, 
    253.9563, 253.9566, 253.9565, 253.9567, 253.9567, 253.9569, 253.9568, 
    253.9572, 253.9571, 253.9574, 253.9573, 253.9574, 253.9574, 253.9574, 
    253.9573, 253.9574, 253.9572, 253.9568, 253.957, 253.9566, 253.9564, 
    253.9562, 253.9561, 253.9561, 253.9562, 253.9563, 253.9565, 253.9566, 
    253.9566, 253.9567, 253.9569, 253.957, 253.9572, 253.9572, 253.9573, 
    253.9573, 253.9574, 253.9574, 253.9575, 253.9573, 253.9574, 253.9572, 
    253.9572, 253.9567, 253.9565, 253.9564, 253.9563, 253.9562, 253.9563, 
    253.9562, 253.9564, 253.9564, 253.9564, 253.9566, 253.9565, 253.957, 
    253.9568, 253.9573, 253.9572, 253.9574, 253.9573, 253.9574, 253.9573, 
    253.9575, 253.9576, 253.9575, 253.9576, 253.9573, 253.9574, 253.9564, 
    253.9564, 253.9564, 253.9563, 253.9563, 253.9562, 253.9563, 253.9563, 
    253.9564, 253.9565, 253.9566, 253.9567, 253.9568, 253.957, 253.9572, 
    253.9573, 253.9572, 253.9573, 253.9572, 253.9572, 253.9575, 253.9574, 
    253.9576, 253.9576, 253.9575, 253.9576, 253.9564, 253.9564, 253.9563, 
    253.9563, 253.9562, 253.9563, 253.9563, 253.9565, 253.9566, 253.9566, 
    253.9567, 253.9568, 253.957, 253.9572, 253.9573, 253.9573, 253.9573, 
    253.9574, 253.9573, 253.9574, 253.9574, 253.9574, 253.9576, 253.9575, 
    253.9576, 253.9576, 253.9564, 253.9564, 253.9564, 253.9565, 253.9564, 
    253.9566, 253.9567, 253.9569, 253.9568, 253.957, 253.9568, 253.9569, 
    253.957, 253.9568, 253.9572, 253.9569, 253.9574, 253.9571, 253.9574, 
    253.9573, 253.9574, 253.9575, 253.9576, 253.9577, 253.9577, 253.9578, 
    253.9565, 253.9566, 253.9566, 253.9567, 253.9567, 253.9569, 253.9571, 
    253.957, 253.9571, 253.9572, 253.9569, 253.9571, 253.9566, 253.9567, 
    253.9567, 253.9565, 253.957, 253.9568, 253.9572, 253.9571, 253.9575, 
    253.9573, 253.9576, 253.9578, 253.958, 253.9581, 253.9566, 253.9566, 
    253.9567, 253.9568, 253.9569, 253.9571, 253.9571, 253.9571, 253.9572, 
    253.9573, 253.9571, 253.9573, 253.9567, 253.957, 253.9566, 253.9567, 
    253.9568, 253.9568, 253.957, 253.957, 253.9572, 253.9571, 253.9578, 
    253.9575, 253.9583, 253.958, 253.9566, 253.9566, 253.9569, 253.9568, 
    253.9571, 253.9572, 253.9572, 253.9573, 253.9573, 253.9574, 253.9573, 
    253.9574, 253.9571, 253.9572, 253.9568, 253.9569, 253.9569, 253.9569, 
    253.957, 253.9571, 253.9571, 253.9572, 253.9573, 253.9571, 253.9578, 
    253.9574, 253.9567, 253.9568, 253.9569, 253.9568, 253.9572, 253.957, 
    253.9574, 253.9573, 253.9574, 253.9574, 253.9574, 253.9573, 253.9572, 
    253.957, 253.9569, 253.9568, 253.9568, 253.957, 253.9572, 253.9573, 
    253.9573, 253.9574, 253.9571, 253.9572, 253.9572, 253.9573, 253.957, 
    253.9573, 253.9569, 253.9569, 253.957, 253.9572, 253.9573, 253.9573, 
    253.9573, 253.9572, 253.9571, 253.957, 253.957, 253.9569, 253.9569, 
    253.9569, 253.957, 253.9572, 253.9573, 253.9575, 253.9575, 253.9577, 
    253.9575, 253.9578, 253.9576, 253.958, 253.9573, 253.9576, 253.957, 
    253.9571, 253.9572, 253.9574, 253.9573, 253.9575, 253.9571, 253.957, 
    253.9569, 253.9568, 253.9569, 253.9569, 253.957, 253.957, 253.9572, 
    253.9571, 253.9574, 253.9575, 253.9578, 253.958, 253.9582, 253.9583, 
    253.9583, 253.9583 ;

 TSA_U =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TSOI =
  254.3909, 254.3923, 254.3921, 254.3932, 254.3926, 254.3933, 254.3912, 
    254.3924, 254.3916, 254.391, 254.3954, 254.3932, 254.3977, 254.3963, 
    254.3999, 254.3975, 254.4004, 254.3998, 254.4015, 254.401, 254.4031, 
    254.4017, 254.4042, 254.4028, 254.403, 254.4017, 254.3937, 254.3951, 
    254.3936, 254.3938, 254.3937, 254.3926, 254.392, 254.3908, 254.391, 
    254.3919, 254.3939, 254.3932, 254.395, 254.3949, 254.3969, 254.396, 
    254.3993, 254.3983, 254.401, 254.4004, 254.401, 254.4008, 254.401, 254.4, 
    254.4004, 254.3996, 254.3962, 254.3972, 254.3942, 254.3924, 254.3913, 
    254.3904, 254.3905, 254.3907, 254.3919, 254.393, 254.3938, 254.3944, 
    254.3949, 254.3965, 254.3974, 254.3994, 254.3991, 254.3997, 254.4003, 
    254.4013, 254.4011, 254.4015, 254.3997, 254.4009, 254.3989, 254.3994, 
    254.395, 254.3934, 254.3927, 254.3921, 254.3906, 254.3916, 254.3912, 
    254.3922, 254.3928, 254.3925, 254.3944, 254.3937, 254.3975, 254.3958, 
    254.4002, 254.3992, 254.4005, 254.3998, 254.4009, 254.3999, 254.4017, 
    254.4021, 254.4018, 254.4028, 254.3999, 254.401, 254.3925, 254.3926, 
    254.3928, 254.3918, 254.3917, 254.3908, 254.3916, 254.392, 254.3929, 
    254.3934, 254.3939, 254.395, 254.3962, 254.398, 254.3992, 254.4001, 
    254.3996, 254.4, 254.3995, 254.3993, 254.4019, 254.4004, 254.4027, 
    254.4026, 254.4015, 254.4026, 254.3926, 254.3923, 254.3913, 254.3921, 
    254.3907, 254.3915, 254.3919, 254.3937, 254.3941, 254.3944, 254.3951, 
    254.396, 254.3976, 254.399, 254.4003, 254.4002, 254.4003, 254.4005, 
    254.3998, 254.4007, 254.4008, 254.4004, 254.4025, 254.4019, 254.4026, 
    254.4022, 254.3924, 254.3929, 254.3926, 254.3931, 254.3928, 254.3943, 
    254.3947, 254.3969, 254.396, 254.3974, 254.3962, 254.3964, 254.3974, 
    254.3963, 254.3989, 254.3971, 254.4006, 254.3987, 254.4007, 254.4003, 
    254.4009, 254.4014, 254.4021, 254.4033, 254.403, 254.4041, 254.3936, 
    254.3942, 254.3942, 254.3948, 254.3953, 254.3964, 254.398, 254.3974, 
    254.3986, 254.3988, 254.397, 254.3981, 254.3946, 254.3952, 254.3949, 
    254.3936, 254.3975, 254.3955, 254.3993, 254.3982, 254.4014, 254.3997, 
    254.4029, 254.4042, 254.4055, 254.407, 254.3946, 254.3941, 254.3949, 
    254.3959, 254.3969, 254.3982, 254.3984, 254.3986, 254.3993, 254.3998, 
    254.3987, 254.3999, 254.3953, 254.3977, 254.394, 254.3951, 254.3959, 
    254.3955, 254.3974, 254.3978, 254.3995, 254.3986, 254.4039, 254.4015, 
    254.4081, 254.4062, 254.394, 254.3946, 254.3965, 254.3956, 254.3983, 
    254.399, 254.3996, 254.4002, 254.4003, 254.4007, 254.4001, 254.4007, 
    254.3982, 254.3993, 254.3963, 254.3971, 254.3967, 254.3964, 254.3975, 
    254.3987, 254.3987, 254.3991, 254.4001, 254.3983, 254.4041, 254.4005, 
    254.3952, 254.3963, 254.3965, 254.396, 254.3989, 254.3979, 254.4007, 
    254.3999, 254.4012, 254.4006, 254.4005, 254.3997, 254.3992, 254.3979, 
    254.3969, 254.3961, 254.3963, 254.3972, 254.3988, 254.4003, 254.4, 
    254.4011, 254.3981, 254.3994, 254.3989, 254.4002, 254.3974, 254.3997, 
    254.3968, 254.3971, 254.3979, 254.3994, 254.3998, 254.4002, 254.4, 
    254.3988, 254.3986, 254.3978, 254.3976, 254.397, 254.3965, 254.397, 
    254.3974, 254.3988, 254.4001, 254.4014, 254.4018, 254.4033, 254.402, 
    254.4041, 254.4023, 254.4055, 254.3998, 254.4023, 254.3979, 254.3984, 
    254.3992, 254.4012, 254.4001, 254.4014, 254.3986, 254.3972, 254.3968, 
    254.3961, 254.3969, 254.3968, 254.3975, 254.3972, 254.3989, 254.398, 
    254.4005, 254.4014, 254.404, 254.4055, 254.4072, 254.4079, 254.4081, 
    254.4082,
  255.5028, 255.5043, 255.504, 255.5052, 255.5045, 255.5053, 255.5031, 
    255.5043, 255.5036, 255.503, 255.5075, 255.5052, 255.5099, 255.5085, 
    255.5121, 255.5096, 255.5126, 255.5121, 255.5138, 255.5133, 255.5154, 
    255.514, 255.5166, 255.5151, 255.5153, 255.514, 255.5057, 255.5072, 
    255.5056, 255.5058, 255.5058, 255.5046, 255.5039, 255.5027, 255.5029, 
    255.5038, 255.5059, 255.5052, 255.507, 255.507, 255.509, 255.5081, 
    255.5115, 255.5105, 255.5133, 255.5126, 255.5133, 255.5131, 255.5133, 
    255.5122, 255.5127, 255.5118, 255.5083, 255.5093, 255.5062, 255.5043, 
    255.5032, 255.5023, 255.5025, 255.5027, 255.5039, 255.505, 255.5059, 
    255.5064, 255.507, 255.5087, 255.5096, 255.5117, 255.5113, 255.5119, 
    255.5125, 255.5135, 255.5134, 255.5138, 255.5119, 255.5132, 255.5111, 
    255.5117, 255.507, 255.5054, 255.5047, 255.5041, 255.5025, 255.5036, 
    255.5032, 255.5042, 255.5048, 255.5045, 255.5064, 255.5057, 255.5096, 
    255.5079, 255.5125, 255.5114, 255.5127, 255.512, 255.5132, 255.5122, 
    255.514, 255.5144, 255.5141, 255.5152, 255.5121, 255.5133, 255.5045, 
    255.5045, 255.5048, 255.5037, 255.5037, 255.5027, 255.5036, 255.5039, 
    255.5049, 255.5054, 255.5059, 255.5071, 255.5083, 255.5101, 255.5114, 
    255.5123, 255.5118, 255.5123, 255.5117, 255.5115, 255.5142, 255.5127, 
    255.515, 255.5149, 255.5138, 255.5149, 255.5046, 255.5043, 255.5033, 
    255.5041, 255.5026, 255.5034, 255.5039, 255.5057, 255.5061, 255.5065, 
    255.5072, 255.5081, 255.5098, 255.5112, 255.5126, 255.5125, 255.5125, 
    255.5128, 255.5121, 255.5129, 255.5131, 255.5127, 255.5149, 255.5143, 
    255.5149, 255.5145, 255.5044, 255.5049, 255.5046, 255.5051, 255.5047, 
    255.5063, 255.5068, 255.509, 255.5081, 255.5096, 255.5083, 255.5085, 
    255.5096, 255.5083, 255.5111, 255.5092, 255.5128, 255.5108, 255.5129, 
    255.5126, 255.5132, 255.5137, 255.5144, 255.5157, 255.5154, 255.5165, 
    255.5056, 255.5062, 255.5062, 255.5069, 255.5074, 255.5085, 255.5102, 
    255.5096, 255.5108, 255.511, 255.5092, 255.5103, 255.5067, 255.5072, 
    255.5069, 255.5057, 255.5097, 255.5076, 255.5115, 255.5103, 255.5136, 
    255.512, 255.5152, 255.5166, 255.518, 255.5195, 255.5066, 255.5062, 
    255.507, 255.508, 255.509, 255.5104, 255.5105, 255.5108, 255.5115, 
    255.512, 255.5109, 255.5122, 255.5073, 255.5099, 255.506, 255.5071, 
    255.508, 255.5076, 255.5095, 255.5099, 255.5117, 255.5108, 255.5163, 
    255.5138, 255.5207, 255.5187, 255.506, 255.5066, 255.5087, 255.5077, 
    255.5105, 255.5112, 255.5118, 255.5125, 255.5126, 255.513, 255.5123, 
    255.513, 255.5104, 255.5116, 255.5084, 255.5092, 255.5089, 255.5085, 
    255.5096, 255.5109, 255.5109, 255.5113, 255.5124, 255.5105, 255.5165, 
    255.5127, 255.5073, 255.5084, 255.5085, 255.5081, 255.5111, 255.51, 
    255.513, 255.5122, 255.5135, 255.5128, 255.5127, 255.5119, 255.5114, 
    255.5101, 255.509, 255.5082, 255.5084, 255.5093, 255.511, 255.5126, 
    255.5122, 255.5134, 255.5103, 255.5116, 255.5111, 255.5124, 255.5095, 
    255.5119, 255.5089, 255.5092, 255.51, 255.5116, 255.5121, 255.5124, 
    255.5122, 255.511, 255.5108, 255.51, 255.5098, 255.5091, 255.5086, 
    255.5091, 255.5096, 255.511, 255.5123, 255.5137, 255.5141, 255.5157, 
    255.5143, 255.5165, 255.5146, 255.518, 255.5121, 255.5146, 255.5101, 
    255.5105, 255.5114, 255.5135, 255.5124, 255.5137, 255.5108, 255.5093, 
    255.5089, 255.5082, 255.509, 255.5089, 255.5096, 255.5094, 255.5111, 
    255.5102, 255.5127, 255.5137, 255.5164, 255.518, 255.5197, 255.5205, 
    255.5207, 255.5208,
  257.1093, 257.1106, 257.1103, 257.1114, 257.1108, 257.1115, 257.1095, 
    257.1106, 257.1099, 257.1094, 257.1135, 257.1115, 257.1157, 257.1144, 
    257.1177, 257.1155, 257.1182, 257.1177, 257.1193, 257.1188, 257.1208, 
    257.1195, 257.1219, 257.1205, 257.1207, 257.1194, 257.1119, 257.1132, 
    257.1118, 257.112, 257.1119, 257.1108, 257.1103, 257.1092, 257.1094, 
    257.1102, 257.1121, 257.1115, 257.1131, 257.113, 257.1149, 257.114, 
    257.1171, 257.1163, 257.1188, 257.1182, 257.1188, 257.1186, 257.1188, 
    257.1179, 257.1183, 257.1174, 257.1142, 257.1151, 257.1123, 257.1106, 
    257.1096, 257.1088, 257.1089, 257.1091, 257.1102, 257.1112, 257.112, 
    257.1125, 257.113, 257.1146, 257.1154, 257.1173, 257.117, 257.1176, 
    257.1181, 257.119, 257.1189, 257.1193, 257.1176, 257.1187, 257.1168, 
    257.1173, 257.1131, 257.1116, 257.1109, 257.1104, 257.109, 257.11, 
    257.1096, 257.1105, 257.1111, 257.1108, 257.1125, 257.1118, 257.1154, 
    257.1139, 257.118, 257.1171, 257.1183, 257.1177, 257.1187, 257.1178, 
    257.1194, 257.1198, 257.1196, 257.1205, 257.1177, 257.1188, 257.1107, 
    257.1108, 257.111, 257.11, 257.11, 257.1092, 257.1099, 257.1102, 
    257.1111, 257.1116, 257.1121, 257.1131, 257.1143, 257.1159, 257.1171, 
    257.1179, 257.1174, 257.1179, 257.1174, 257.1172, 257.1197, 257.1183, 
    257.1204, 257.1203, 257.1193, 257.1203, 257.1108, 257.1106, 257.1096, 
    257.1104, 257.1091, 257.1098, 257.1102, 257.1118, 257.1122, 257.1125, 
    257.1132, 257.1141, 257.1156, 257.1169, 257.1182, 257.1181, 257.1181, 
    257.1183, 257.1177, 257.1185, 257.1186, 257.1183, 257.1203, 257.1197, 
    257.1203, 257.1199, 257.1107, 257.1111, 257.1109, 257.1113, 257.111, 
    257.1124, 257.1129, 257.1149, 257.1141, 257.1154, 257.1142, 257.1144, 
    257.1154, 257.1143, 257.1168, 257.1151, 257.1184, 257.1165, 257.1185, 
    257.1181, 257.1187, 257.1192, 257.1199, 257.121, 257.1208, 257.1218, 
    257.1118, 257.1124, 257.1123, 257.1129, 257.1134, 257.1144, 257.116, 
    257.1154, 257.1165, 257.1167, 257.115, 257.116, 257.1128, 257.1133, 
    257.113, 257.1118, 257.1155, 257.1136, 257.1171, 257.1161, 257.1191, 
    257.1176, 257.1206, 257.1219, 257.1231, 257.1245, 257.1127, 257.1123, 
    257.113, 257.114, 257.1149, 257.1161, 257.1163, 257.1165, 257.1171, 
    257.1176, 257.1166, 257.1178, 257.1133, 257.1157, 257.1121, 257.1132, 
    257.1139, 257.1136, 257.1153, 257.1157, 257.1173, 257.1165, 257.1216, 
    257.1193, 257.1257, 257.1239, 257.1122, 257.1127, 257.1146, 257.1137, 
    257.1162, 257.1169, 257.1174, 257.1181, 257.1181, 257.1185, 257.1179, 
    257.1185, 257.1161, 257.1172, 257.1143, 257.1151, 257.1147, 257.1144, 
    257.1154, 257.1166, 257.1166, 257.117, 257.118, 257.1163, 257.1218, 
    257.1183, 257.1133, 257.1143, 257.1145, 257.1141, 257.1168, 257.1158, 
    257.1185, 257.1178, 257.119, 257.1184, 257.1183, 257.1176, 257.1171, 
    257.1158, 257.1149, 257.1141, 257.1143, 257.1151, 257.1167, 257.1181, 
    257.1178, 257.1189, 257.1161, 257.1172, 257.1168, 257.118, 257.1154, 
    257.1175, 257.1148, 257.1151, 257.1158, 257.1173, 257.1177, 257.118, 
    257.1178, 257.1167, 257.1165, 257.1158, 257.1156, 257.115, 257.1145, 
    257.1149, 257.1154, 257.1167, 257.1179, 257.1192, 257.1195, 257.121, 
    257.1198, 257.1218, 257.1201, 257.1231, 257.1177, 257.12, 257.1158, 
    257.1163, 257.1171, 257.119, 257.118, 257.1192, 257.1165, 257.1151, 
    257.1148, 257.1142, 257.1148, 257.1148, 257.1154, 257.1152, 257.1168, 
    257.1159, 257.1183, 257.1192, 257.1216, 257.1232, 257.1248, 257.1255, 
    257.1257, 257.1258,
  259.2228, 259.2238, 259.2236, 259.2244, 259.224, 259.2245, 259.223, 
    259.2238, 259.2233, 259.2229, 259.2259, 259.2244, 259.2275, 259.2266, 
    259.229, 259.2274, 259.2294, 259.229, 259.2302, 259.2298, 259.2313, 
    259.2303, 259.2321, 259.2311, 259.2312, 259.2303, 259.2247, 259.2257, 
    259.2247, 259.2248, 259.2248, 259.224, 259.2236, 259.2228, 259.2229, 
    259.2235, 259.2249, 259.2244, 259.2256, 259.2256, 259.2269, 259.2263, 
    259.2286, 259.2279, 259.2298, 259.2293, 259.2298, 259.2297, 259.2298, 
    259.2291, 259.2294, 259.2288, 259.2264, 259.2271, 259.2251, 259.2238, 
    259.2231, 259.2225, 259.2226, 259.2227, 259.2235, 259.2242, 259.2248, 
    259.2252, 259.2256, 259.2267, 259.2273, 259.2287, 259.2285, 259.2289, 
    259.2293, 259.23, 259.2299, 259.2302, 259.2289, 259.2297, 259.2283, 
    259.2287, 259.2256, 259.2245, 259.224, 259.2237, 259.2227, 259.2233, 
    259.2231, 259.2237, 259.2242, 259.2239, 259.2252, 259.2247, 259.2274, 
    259.2262, 259.2292, 259.2285, 259.2294, 259.229, 259.2298, 259.2291, 
    259.2303, 259.2306, 259.2304, 259.2311, 259.229, 259.2298, 259.2239, 
    259.224, 259.2241, 259.2234, 259.2234, 259.2228, 259.2233, 259.2235, 
    259.2242, 259.2245, 259.2249, 259.2256, 259.2265, 259.2277, 259.2286, 
    259.2292, 259.2288, 259.2291, 259.2288, 259.2286, 259.2305, 259.2294, 
    259.231, 259.2309, 259.2302, 259.2309, 259.224, 259.2238, 259.2231, 
    259.2236, 259.2227, 259.2232, 259.2235, 259.2247, 259.225, 259.2252, 
    259.2257, 259.2263, 259.2274, 259.2284, 259.2293, 259.2293, 259.2293, 
    259.2295, 259.229, 259.2296, 259.2297, 259.2294, 259.2309, 259.2305, 
    259.2309, 259.2307, 259.2238, 259.2242, 259.224, 259.2243, 259.2241, 
    259.2251, 259.2254, 259.2269, 259.2263, 259.2273, 259.2264, 259.2266, 
    259.2273, 259.2265, 259.2284, 259.2271, 259.2295, 259.2281, 259.2296, 
    259.2293, 259.2297, 259.2301, 259.2306, 259.2315, 259.2313, 259.232, 
    259.2247, 259.2251, 259.2251, 259.2255, 259.2258, 259.2266, 259.2277, 
    259.2273, 259.2281, 259.2283, 259.227, 259.2278, 259.2254, 259.2257, 
    259.2255, 259.2247, 259.2274, 259.226, 259.2286, 259.2278, 259.2301, 
    259.2289, 259.2312, 259.2321, 259.2331, 259.2341, 259.2253, 259.225, 
    259.2256, 259.2263, 259.227, 259.2279, 259.228, 259.2281, 259.2286, 
    259.2289, 259.2282, 259.229, 259.2258, 259.2275, 259.2249, 259.2257, 
    259.2262, 259.226, 259.2272, 259.2275, 259.2287, 259.2281, 259.2319, 
    259.2302, 259.235, 259.2336, 259.2249, 259.2253, 259.2267, 259.226, 
    259.2279, 259.2284, 259.2288, 259.2293, 259.2293, 259.2296, 259.2292, 
    259.2296, 259.2279, 259.2286, 259.2265, 259.2271, 259.2268, 259.2266, 
    259.2274, 259.2282, 259.2282, 259.2285, 259.2292, 259.2279, 259.2321, 
    259.2295, 259.2257, 259.2265, 259.2266, 259.2263, 259.2283, 259.2276, 
    259.2296, 259.2291, 259.2299, 259.2295, 259.2295, 259.2289, 259.2285, 
    259.2276, 259.2269, 259.2264, 259.2265, 259.2271, 259.2282, 259.2293, 
    259.2291, 259.2299, 259.2278, 259.2287, 259.2283, 259.2292, 259.2273, 
    259.2289, 259.2269, 259.2271, 259.2276, 259.2287, 259.229, 259.2292, 
    259.2291, 259.2283, 259.2281, 259.2276, 259.2274, 259.227, 259.2267, 
    259.227, 259.2273, 259.2283, 259.2292, 259.2301, 259.2304, 259.2315, 
    259.2306, 259.2321, 259.2307, 259.2331, 259.229, 259.2307, 259.2276, 
    259.228, 259.2285, 259.2299, 259.2292, 259.2301, 259.2281, 259.2271, 
    259.2269, 259.2264, 259.2269, 259.2269, 259.2273, 259.2272, 259.2283, 
    259.2277, 259.2294, 259.2301, 259.2319, 259.2331, 259.2343, 259.2348, 
    259.235, 259.235,
  261.4069, 261.4073, 261.4072, 261.4076, 261.4074, 261.4076, 261.407, 
    261.4073, 261.4071, 261.4069, 261.4083, 261.4076, 261.4091, 261.4086, 
    261.4098, 261.409, 261.41, 261.4098, 261.4104, 261.4102, 261.4109, 
    261.4104, 261.4113, 261.4108, 261.4109, 261.4104, 261.4077, 261.4082, 
    261.4077, 261.4078, 261.4077, 261.4074, 261.4072, 261.4068, 261.4069, 
    261.4072, 261.4078, 261.4076, 261.4081, 261.4081, 261.4088, 261.4085, 
    261.4096, 261.4093, 261.4102, 261.41, 261.4102, 261.4101, 261.4102, 
    261.4099, 261.41, 261.4097, 261.4085, 261.4089, 261.4079, 261.4073, 
    261.407, 261.4067, 261.4067, 261.4068, 261.4072, 261.4075, 261.4078, 
    261.408, 261.4081, 261.4087, 261.409, 261.4096, 261.4095, 261.4097, 
    261.4099, 261.4103, 261.4102, 261.4104, 261.4097, 261.4102, 261.4095, 
    261.4096, 261.4081, 261.4077, 261.4074, 261.4072, 261.4068, 261.4071, 
    261.407, 261.4073, 261.4074, 261.4073, 261.408, 261.4077, 261.409, 
    261.4084, 261.4099, 261.4095, 261.41, 261.4098, 261.4102, 261.4098, 
    261.4104, 261.4106, 261.4105, 261.4108, 261.4098, 261.4102, 261.4073, 
    261.4074, 261.4074, 261.4071, 261.4071, 261.4068, 261.4071, 261.4072, 
    261.4075, 261.4076, 261.4078, 261.4081, 261.4086, 261.4091, 261.4096, 
    261.4099, 261.4097, 261.4099, 261.4097, 261.4096, 261.4105, 261.41, 
    261.4108, 261.4107, 261.4104, 261.4107, 261.4074, 261.4073, 261.407, 
    261.4072, 261.4068, 261.407, 261.4072, 261.4077, 261.4079, 261.408, 
    261.4082, 261.4085, 261.409, 261.4095, 261.4099, 261.4099, 261.4099, 
    261.41, 261.4098, 261.4101, 261.4101, 261.41, 261.4107, 261.4105, 
    261.4107, 261.4106, 261.4073, 261.4075, 261.4074, 261.4075, 261.4074, 
    261.4079, 261.4081, 261.4088, 261.4085, 261.409, 261.4085, 261.4086, 
    261.409, 261.4086, 261.4095, 261.4088, 261.41, 261.4094, 261.4101, 
    261.4099, 261.4102, 261.4103, 261.4106, 261.411, 261.4109, 261.4113, 
    261.4077, 261.4079, 261.4079, 261.4081, 261.4083, 261.4086, 261.4092, 
    261.409, 261.4094, 261.4094, 261.4088, 261.4092, 261.4081, 261.4082, 
    261.4081, 261.4077, 261.409, 261.4083, 261.4096, 261.4092, 261.4103, 
    261.4098, 261.4109, 261.4113, 261.4118, 261.4124, 261.408, 261.4079, 
    261.4081, 261.4084, 261.4088, 261.4092, 261.4093, 261.4094, 261.4096, 
    261.4098, 261.4094, 261.4098, 261.4082, 261.4091, 261.4078, 261.4082, 
    261.4084, 261.4083, 261.4089, 261.4091, 261.4097, 261.4094, 261.4112, 
    261.4104, 261.4128, 261.4121, 261.4078, 261.408, 261.4087, 261.4084, 
    261.4093, 261.4095, 261.4097, 261.4099, 261.4099, 261.4101, 261.4099, 
    261.4101, 261.4092, 261.4096, 261.4086, 261.4088, 261.4087, 261.4086, 
    261.409, 261.4094, 261.4094, 261.4095, 261.4099, 261.4093, 261.4113, 
    261.41, 261.4082, 261.4086, 261.4086, 261.4085, 261.4095, 261.4091, 
    261.4101, 261.4098, 261.4103, 261.41, 261.41, 261.4097, 261.4095, 
    261.4091, 261.4088, 261.4085, 261.4086, 261.4089, 261.4094, 261.4099, 
    261.4098, 261.4102, 261.4092, 261.4096, 261.4095, 261.4099, 261.4089, 
    261.4097, 261.4088, 261.4088, 261.4091, 261.4096, 261.4098, 261.4099, 
    261.4098, 261.4094, 261.4094, 261.4091, 261.409, 261.4088, 261.4087, 
    261.4088, 261.409, 261.4094, 261.4099, 261.4103, 261.4105, 261.411, 
    261.4106, 261.4113, 261.4106, 261.4118, 261.4098, 261.4106, 261.4091, 
    261.4093, 261.4096, 261.4102, 261.4099, 261.4103, 261.4094, 261.4089, 
    261.4088, 261.4085, 261.4088, 261.4088, 261.409, 261.4089, 261.4095, 
    261.4091, 261.41, 261.4103, 261.4113, 261.4118, 261.4124, 261.4127, 
    261.4128, 261.4128,
  262.7627, 262.7628, 262.7628, 262.7629, 262.7628, 262.7629, 262.7627, 
    262.7628, 262.7628, 262.7627, 262.763, 262.7629, 262.7632, 262.7631, 
    262.7634, 262.7632, 262.7635, 262.7634, 262.7635, 262.7635, 262.7637, 
    262.7636, 262.7638, 262.7637, 262.7637, 262.7635, 262.7629, 262.763, 
    262.7629, 262.7629, 262.7629, 262.7628, 262.7628, 262.7627, 262.7627, 
    262.7628, 262.7629, 262.7629, 262.763, 262.763, 262.7632, 262.7631, 
    262.7634, 262.7633, 262.7635, 262.7635, 262.7635, 262.7635, 262.7635, 
    262.7634, 262.7635, 262.7634, 262.7631, 262.7632, 262.7629, 262.7628, 
    262.7628, 262.7627, 262.7627, 262.7627, 262.7628, 262.7629, 262.7629, 
    262.763, 262.763, 262.7631, 262.7632, 262.7634, 262.7633, 262.7634, 
    262.7635, 262.7635, 262.7635, 262.7635, 262.7634, 262.7635, 262.7633, 
    262.7634, 262.763, 262.7629, 262.7628, 262.7628, 262.7627, 262.7628, 
    262.7628, 262.7628, 262.7628, 262.7628, 262.763, 262.7629, 262.7632, 
    262.7631, 262.7634, 262.7633, 262.7635, 262.7634, 262.7635, 262.7634, 
    262.7636, 262.7636, 262.7636, 262.7637, 262.7634, 262.7635, 262.7628, 
    262.7628, 262.7628, 262.7628, 262.7628, 262.7627, 262.7628, 262.7628, 
    262.7628, 262.7629, 262.7629, 262.763, 262.7631, 262.7632, 262.7634, 
    262.7634, 262.7634, 262.7634, 262.7634, 262.7634, 262.7636, 262.7635, 
    262.7636, 262.7636, 262.7635, 262.7636, 262.7628, 262.7628, 262.7628, 
    262.7628, 262.7627, 262.7628, 262.7628, 262.7629, 262.7629, 262.763, 
    262.763, 262.7631, 262.7632, 262.7633, 262.7635, 262.7634, 262.7634, 
    262.7635, 262.7634, 262.7635, 262.7635, 262.7635, 262.7636, 262.7636, 
    262.7636, 262.7636, 262.7628, 262.7628, 262.7628, 262.7629, 262.7628, 
    262.763, 262.763, 262.7632, 262.7631, 262.7632, 262.7631, 262.7631, 
    262.7632, 262.7631, 262.7633, 262.7632, 262.7635, 262.7633, 262.7635, 
    262.7635, 262.7635, 262.7635, 262.7636, 262.7637, 262.7637, 262.7638, 
    262.7629, 262.763, 262.7629, 262.763, 262.763, 262.7631, 262.7632, 
    262.7632, 262.7633, 262.7633, 262.7632, 262.7633, 262.763, 262.763, 
    262.763, 262.7629, 262.7632, 262.7631, 262.7634, 262.7633, 262.7635, 
    262.7634, 262.7637, 262.7638, 262.7639, 262.7641, 262.763, 262.7629, 
    262.763, 262.7631, 262.7632, 262.7633, 262.7633, 262.7633, 262.7634, 
    262.7634, 262.7633, 262.7634, 262.763, 262.7632, 262.7629, 262.763, 
    262.7631, 262.7631, 262.7632, 262.7632, 262.7634, 262.7633, 262.7638, 
    262.7635, 262.7642, 262.764, 262.7629, 262.763, 262.7631, 262.7631, 
    262.7633, 262.7633, 262.7634, 262.7634, 262.7635, 262.7635, 262.7634, 
    262.7635, 262.7633, 262.7634, 262.7631, 262.7632, 262.7632, 262.7631, 
    262.7632, 262.7633, 262.7633, 262.7633, 262.7634, 262.7633, 262.7638, 
    262.7635, 262.763, 262.7631, 262.7631, 262.7631, 262.7633, 262.7632, 
    262.7635, 262.7634, 262.7635, 262.7635, 262.7635, 262.7634, 262.7633, 
    262.7632, 262.7632, 262.7631, 262.7631, 262.7632, 262.7633, 262.7635, 
    262.7634, 262.7635, 262.7633, 262.7634, 262.7633, 262.7634, 262.7632, 
    262.7634, 262.7632, 262.7632, 262.7632, 262.7634, 262.7634, 262.7634, 
    262.7634, 262.7633, 262.7633, 262.7632, 262.7632, 262.7632, 262.7631, 
    262.7632, 262.7632, 262.7633, 262.7634, 262.7635, 262.7636, 262.7637, 
    262.7636, 262.7638, 262.7636, 262.7639, 262.7634, 262.7636, 262.7632, 
    262.7633, 262.7634, 262.7635, 262.7634, 262.7635, 262.7633, 262.7632, 
    262.7632, 262.7631, 262.7632, 262.7632, 262.7632, 262.7632, 262.7633, 
    262.7632, 262.7635, 262.7635, 262.7638, 262.7639, 262.7641, 262.7642, 
    262.7642, 262.7642,
  263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1178, 263.1177, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1179, 263.1178, 263.1178, 263.1178, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1177, 263.1177, 263.1177, 263.1177, 263.1177, 
    263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1179, 
    263.1177, 263.1177, 263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 263.1178, 
    263.1177, 263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1179, 263.1179, 263.1179, 263.1177, 263.1177, 
    263.1177, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1177, 263.1177, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1179, 263.1179, 263.1177, 263.1177, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1179, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1179, 263.1178, 263.1179, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 263.1178, 
    263.1178, 263.1178, 263.1178, 263.1179, 263.1179, 263.1179, 263.1179, 
    263.1179, 263.1179,
  263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 263.1491, 
    263.1491, 263.1491,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15,
  263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 263.15, 
    263.15, 263.15, 263.15, 263.15, 263.15 ;

 TSOI_10CM =
  262.919, 262.9334, 262.9306, 262.9423, 262.9358, 262.9434, 262.9219, 
    262.934, 262.9263, 262.9203, 262.9647, 262.9428, 262.9875, 262.9735, 
    263.0085, 262.9853, 263.0132, 263.0079, 263.024, 263.0194, 263.0399, 
    263.0261, 263.0505, 263.0366, 263.0388, 263.0257, 262.9472, 262.9619, 
    262.9463, 262.9484, 262.9475, 262.9359, 262.9301, 262.9179, 262.9201, 
    262.9291, 262.9494, 262.9425, 262.9598, 262.9594, 262.9787, 262.97, 
    263.0023, 262.9931, 263.0196, 263.0129, 263.0193, 263.0174, 263.0193, 
    263.0096, 263.0137, 263.0052, 262.9716, 262.9815, 262.9521, 262.9343, 
    262.9225, 262.914, 262.9152, 262.9175, 262.9291, 262.9401, 262.9484, 
    262.9539, 262.9594, 262.9759, 262.9846, 263.0042, 263.0006, 263.0066, 
    263.0123, 263.0218, 263.0203, 263.0244, 263.0064, 263.0184, 262.9986, 
    263.0041, 262.9608, 262.9444, 262.9373, 262.9312, 262.9161, 262.9265, 
    262.9224, 262.9322, 262.9383, 262.9353, 262.9541, 262.9468, 262.9851, 
    262.9686, 263.0116, 263.0014, 263.0141, 263.0076, 263.0187, 263.0087, 
    263.026, 263.0298, 263.0272, 263.0371, 263.0081, 263.0193, 262.9352, 
    262.9357, 262.938, 262.9278, 262.9272, 262.9178, 262.9261, 262.9297, 
    262.9387, 262.944, 262.949, 262.9601, 262.9724, 262.9897, 263.002, 
    263.0103, 263.0052, 263.0097, 263.0047, 263.0023, 263.0284, 263.0138, 
    263.0357, 263.0345, 263.0245, 263.0346, 262.9361, 262.9332, 262.9232, 
    262.931, 262.9168, 262.9247, 262.9293, 262.9469, 262.9508, 262.9543, 
    262.9614, 262.9705, 262.9863, 263.0001, 263.0126, 263.0117, 263.012, 
    263.0148, 263.0079, 263.016, 263.0173, 263.0138, 263.0343, 263.0284, 
    263.0345, 263.0306, 262.9341, 262.9389, 262.9363, 262.9412, 262.9378, 
    262.9531, 262.9576, 262.979, 262.9703, 262.9843, 262.9717, 262.9739, 
    262.9846, 262.9724, 262.9993, 262.981, 263.0149, 262.9967, 263.0161, 
    263.0126, 263.0184, 263.0236, 263.0301, 263.0421, 263.0393, 263.0494, 
    262.9461, 262.9523, 262.9518, 262.9583, 262.9631, 262.9735, 262.9902, 
    262.984, 262.9955, 262.9978, 262.9803, 262.991, 262.9565, 262.9621, 
    262.9588, 262.9466, 262.9854, 262.9655, 263.0022, 262.9915, 263.0228, 
    263.0072, 263.0378, 263.0508, 263.063, 263.0772, 262.9557, 262.9515, 
    262.9591, 262.9695, 262.9792, 262.9921, 262.9934, 262.9958, 263.0021, 
    263.0074, 262.9966, 263.0087, 262.9633, 262.9871, 262.9499, 262.9611, 
    262.9689, 262.9655, 262.9832, 262.9874, 263.0044, 262.9956, 263.0476, 
    263.0246, 263.088, 263.0704, 262.95, 262.9557, 262.9755, 262.9661, 
    262.993, 262.9996, 263.005, 263.0118, 263.0125, 263.0166, 263.01, 
    263.0164, 262.9922, 263.003, 262.9733, 262.9805, 262.9772, 262.9735, 
    262.9848, 262.9968, 262.997, 263.0009, 263.0116, 262.9931, 263.0505, 
    263.0151, 262.9619, 262.9728, 262.9744, 262.9702, 262.9989, 262.9885, 
    263.0165, 263.009, 263.0213, 263.0152, 263.0143, 263.0064, 263.0015, 
    262.989, 262.9789, 262.9708, 262.9727, 262.9815, 262.9975, 263.0126, 
    263.0093, 263.0204, 262.9911, 263.0034, 262.9986, 263.011, 262.9838, 
    263.0069, 262.9779, 262.9804, 262.9883, 263.0042, 263.0077, 263.0114, 
    263.0092, 262.9979, 262.9961, 262.9881, 262.9859, 262.9799, 262.9749, 
    262.9794, 262.9843, 262.9979, 263.0102, 263.0236, 263.0269, 263.0425, 
    263.0298, 263.0507, 263.0329, 263.0637, 263.0083, 263.0324, 262.9887, 
    262.9934, 263.0019, 263.0215, 263.011, 263.0233, 262.996, 262.9818, 
    262.9782, 262.9713, 262.9783, 262.9778, 262.9845, 262.9823, 262.9984, 
    262.9897, 263.0143, 263.0232, 263.0483, 263.0636, 263.0792, 263.086, 
    263.0881, 263.089 ;

 TSOI_ICE =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 TV =
  253.9048, 253.9056, 253.9054, 253.9061, 253.9057, 253.9062, 253.9049, 
    253.9056, 253.9052, 253.9048, 253.9074, 253.9061, 253.9088, 253.908, 
    253.91, 253.9086, 253.9103, 253.91, 253.911, 253.9107, 253.9119, 
    253.9111, 253.9126, 253.9117, 253.9118, 253.9111, 253.9064, 253.9072, 
    253.9064, 253.9065, 253.9064, 253.9057, 253.9054, 253.9047, 253.9048, 
    253.9053, 253.9065, 253.9061, 253.9072, 253.9072, 253.9083, 253.9078, 
    253.9097, 253.9091, 253.9107, 253.9103, 253.9107, 253.9106, 253.9107, 
    253.9101, 253.9104, 253.9099, 253.9079, 253.9084, 253.9067, 253.9056, 
    253.905, 253.9045, 253.9045, 253.9047, 253.9053, 253.906, 253.9065, 
    253.9068, 253.9071, 253.9081, 253.9086, 253.9098, 253.9096, 253.9099, 
    253.9103, 253.9108, 253.9108, 253.911, 253.9099, 253.9106, 253.9095, 
    253.9098, 253.9072, 253.9062, 253.9058, 253.9055, 253.9046, 253.9052, 
    253.905, 253.9055, 253.9059, 253.9057, 253.9068, 253.9064, 253.9086, 
    253.9077, 253.9102, 253.9096, 253.9104, 253.91, 253.9107, 253.9101, 
    253.9111, 253.9113, 253.9112, 253.9118, 253.91, 253.9107, 253.9057, 
    253.9057, 253.9059, 253.9053, 253.9052, 253.9047, 253.9052, 253.9054, 
    253.9059, 253.9062, 253.9065, 253.9072, 253.9079, 253.9089, 253.9097, 
    253.9102, 253.9099, 253.9101, 253.9098, 253.9097, 253.9112, 253.9104, 
    253.9117, 253.9116, 253.911, 253.9116, 253.9058, 253.9056, 253.905, 
    253.9055, 253.9046, 253.9051, 253.9053, 253.9064, 253.9066, 253.9068, 
    253.9073, 253.9078, 253.9087, 253.9095, 253.9103, 253.9102, 253.9103, 
    253.9104, 253.91, 253.9105, 253.9106, 253.9104, 253.9116, 253.9113, 
    253.9116, 253.9114, 253.9057, 253.9059, 253.9058, 253.9061, 253.9059, 
    253.9068, 253.907, 253.9083, 253.9078, 253.9086, 253.9079, 253.908, 
    253.9086, 253.9079, 253.9095, 253.9084, 253.9104, 253.9093, 253.9105, 
    253.9103, 253.9106, 253.9109, 253.9113, 253.9121, 253.9119, 253.9125, 
    253.9064, 253.9067, 253.9067, 253.9071, 253.9073, 253.908, 253.909, 
    253.9086, 253.9093, 253.9094, 253.9084, 253.909, 253.907, 253.9073, 
    253.9071, 253.9064, 253.9087, 253.9075, 253.9097, 253.909, 253.9109, 
    253.91, 253.9118, 253.9126, 253.9133, 253.9142, 253.9069, 253.9067, 
    253.9071, 253.9077, 253.9083, 253.9091, 253.9092, 253.9093, 253.9097, 
    253.91, 253.9093, 253.9101, 253.9073, 253.9088, 253.9066, 253.9072, 
    253.9077, 253.9075, 253.9086, 253.9088, 253.9098, 253.9093, 253.9124, 
    253.911, 253.9149, 253.9138, 253.9066, 253.9069, 253.9081, 253.9075, 
    253.9091, 253.9095, 253.9099, 253.9102, 253.9103, 253.9105, 253.9101, 
    253.9105, 253.9091, 253.9097, 253.908, 253.9084, 253.9082, 253.908, 
    253.9086, 253.9093, 253.9094, 253.9096, 253.9102, 253.9091, 253.9125, 
    253.9104, 253.9073, 253.9079, 253.908, 253.9078, 253.9095, 253.9089, 
    253.9105, 253.9101, 253.9108, 253.9104, 253.9104, 253.9099, 253.9096, 
    253.9089, 253.9083, 253.9078, 253.9079, 253.9084, 253.9094, 253.9103, 
    253.9101, 253.9108, 253.909, 253.9097, 253.9095, 253.9102, 253.9086, 
    253.9099, 253.9082, 253.9084, 253.9088, 253.9098, 253.91, 253.9102, 
    253.9101, 253.9094, 253.9093, 253.9088, 253.9087, 253.9084, 253.9081, 
    253.9083, 253.9086, 253.9094, 253.9102, 253.9109, 253.9112, 253.912, 
    253.9113, 253.9125, 253.9115, 253.9133, 253.91, 253.9115, 253.9089, 
    253.9091, 253.9097, 253.9108, 253.9102, 253.9109, 253.9093, 253.9084, 
    253.9082, 253.9078, 253.9083, 253.9082, 253.9086, 253.9085, 253.9095, 
    253.9089, 253.9104, 253.9109, 253.9124, 253.9134, 253.9143, 253.9147, 
    253.9149, 253.9149 ;

 TWS =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 T_SCALAR =
  0.1399993, 0.1400072, 0.1400057, 0.1400119, 0.1400085, 0.1400126, 0.140001, 
    0.1400074, 0.1400033, 0.1400001, 0.1400239, 0.1400122, 0.1400368, 
    0.1400292, 0.1400485, 0.1400355, 0.1400512, 0.1400483, 0.1400574, 
    0.1400548, 0.1400661, 0.1400586, 0.1400722, 0.1400644, 0.1400655, 
    0.1400583, 0.1400147, 0.1400224, 0.1400142, 0.1400153, 0.1400149, 
    0.1400085, 0.1400052, 0.1399988, 0.14, 0.1400048, 0.1400158, 0.1400122, 
    0.1400217, 0.1400215, 0.140032, 0.1400273, 0.1400452, 0.1400401, 
    0.1400549, 0.1400511, 0.1400547, 0.1400536, 0.1400547, 0.1400492, 
    0.1400516, 0.1400468, 0.1400281, 0.1400335, 0.1400173, 0.1400074, 
    0.1400012, 0.1399967, 0.1399973, 0.1399985, 0.1400048, 0.1400108, 
    0.1400154, 0.1400184, 0.1400215, 0.1400302, 0.1400352, 0.1400461, 
    0.1400443, 0.1400475, 0.1400508, 0.1400561, 0.1400553, 0.1400576, 
    0.1400475, 0.1400541, 0.1400432, 0.1400462, 0.1400217, 0.1400132, 
    0.1400091, 0.1400059, 0.1399978, 0.1400034, 0.1400012, 0.1400065, 
    0.1400099, 0.1400083, 0.1400185, 0.1400145, 0.1400355, 0.1400264, 
    0.1400504, 0.1400447, 0.1400518, 0.1400482, 0.1400543, 0.1400488, 
    0.1400585, 0.1400605, 0.1400591, 0.1400647, 0.1400485, 0.1400546, 
    0.1400082, 0.1400084, 0.1400097, 0.1400041, 0.1400038, 0.1399987, 
    0.1400032, 0.1400051, 0.1400101, 0.140013, 0.1400157, 0.1400218, 
    0.1400285, 0.1400381, 0.140045, 0.1400497, 0.1400469, 0.1400494, 
    0.1400466, 0.1400453, 0.1400597, 0.1400515, 0.1400639, 0.1400633, 
    0.1400576, 0.1400633, 0.1400086, 0.1400071, 0.1400016, 0.1400059, 
    0.1399982, 0.1400025, 0.1400049, 0.1400145, 0.1400167, 0.1400186, 
    0.1400225, 0.1400275, 0.1400362, 0.1400439, 0.140051, 0.1400505, 
    0.1400506, 0.1400522, 0.1400483, 0.1400528, 0.1400535, 0.1400516, 
    0.1400632, 0.1400599, 0.1400632, 0.1400611, 0.1400076, 0.1400102, 
    0.1400088, 0.1400114, 0.1400095, 0.1400178, 0.1400203, 0.1400321, 
    0.1400274, 0.140035, 0.1400282, 0.1400294, 0.1400351, 0.1400286, 
    0.1400433, 0.1400331, 0.1400522, 0.1400418, 0.1400529, 0.140051, 
    0.1400542, 0.1400571, 0.1400608, 0.1400675, 0.1400659, 0.1400716, 
    0.1400141, 0.1400175, 0.1400173, 0.1400208, 0.1400234, 0.1400292, 
    0.1400384, 0.140035, 0.1400414, 0.1400427, 0.140033, 0.1400388, 
    0.1400198, 0.1400227, 0.1400211, 0.1400144, 0.1400357, 0.1400246, 
    0.1400451, 0.1400391, 0.1400567, 0.1400478, 0.1400651, 0.1400722, 
    0.1400794, 0.1400873, 0.1400194, 0.1400171, 0.1400213, 0.1400269, 
    0.1400324, 0.1400395, 0.1400403, 0.1400416, 0.1400451, 0.140048, 
    0.1400419, 0.1400488, 0.1400232, 0.1400367, 0.1400162, 0.1400222, 
    0.1400266, 0.1400248, 0.1400346, 0.1400369, 0.1400463, 0.1400415, 
    0.1400703, 0.1400575, 0.1400937, 0.1400835, 0.1400163, 0.1400194, 
    0.1400302, 0.1400251, 0.14004, 0.1400437, 0.1400467, 0.1400505, 
    0.1400509, 0.1400532, 0.1400495, 0.1400531, 0.1400395, 0.1400456, 
    0.1400291, 0.1400331, 0.1400313, 0.1400293, 0.1400355, 0.140042, 
    0.1400423, 0.1400443, 0.1400498, 0.1400401, 0.1400717, 0.1400518, 
    0.1400228, 0.1400287, 0.1400297, 0.1400274, 0.1400433, 0.1400375, 
    0.1400531, 0.1400489, 0.1400559, 0.1400524, 0.1400519, 0.1400475, 
    0.1400447, 0.1400377, 0.1400321, 0.1400278, 0.1400288, 0.1400336, 
    0.1400424, 0.1400509, 0.140049, 0.1400553, 0.1400389, 0.1400457, 
    0.140043, 0.1400501, 0.1400349, 0.1400473, 0.1400317, 0.1400331, 
    0.1400374, 0.1400461, 0.1400482, 0.1400502, 0.140049, 0.1400427, 
    0.1400417, 0.1400373, 0.140036, 0.1400328, 0.14003, 0.1400325, 0.1400351, 
    0.1400427, 0.1400496, 0.1400571, 0.140059, 0.1400674, 0.1400603, 
    0.1400718, 0.1400617, 0.1400794, 0.1400483, 0.1400617, 0.1400376, 
    0.1400403, 0.1400449, 0.1400557, 0.14005, 0.1400568, 0.1400417, 
    0.1400337, 0.1400318, 0.140028, 0.1400319, 0.1400316, 0.1400353, 
    0.1400341, 0.140043, 0.1400382, 0.1400518, 0.1400568, 0.140071, 
    0.1400796, 0.1400887, 0.1400926, 0.1400939, 0.1400944,
  0.1463936, 0.1464023, 0.1464007, 0.1464076, 0.1464038, 0.1464083, 
    0.1463954, 0.1464026, 0.1463981, 0.1463945, 0.146421, 0.1464079, 
    0.1464353, 0.1464268, 0.1464484, 0.1464339, 0.1464514, 0.1464481, 
    0.1464583, 0.1464554, 0.146468, 0.1464596, 0.1464749, 0.1464661, 
    0.1464674, 0.1464593, 0.1464107, 0.1464193, 0.1464102, 0.1464114, 
    0.1464109, 0.1464038, 0.1464002, 0.146393, 0.1463944, 0.1463997, 
    0.146412, 0.1464079, 0.1464185, 0.1464183, 0.14643, 0.1464247, 0.1464446, 
    0.146439, 0.1464555, 0.1464513, 0.1464553, 0.1464541, 0.1464553, 
    0.1464491, 0.1464518, 0.1464464, 0.1464256, 0.1464317, 0.1464136, 
    0.1464026, 0.1463957, 0.1463907, 0.1463914, 0.1463927, 0.1463997, 
    0.1464064, 0.1464115, 0.1464149, 0.1464182, 0.146428, 0.1464335, 
    0.1464457, 0.1464436, 0.1464472, 0.1464509, 0.1464568, 0.1464559, 
    0.1464585, 0.1464472, 0.1464546, 0.1464424, 0.1464457, 0.1464186, 
    0.146409, 0.1464045, 0.146401, 0.146392, 0.1463981, 0.1463957, 0.1464016, 
    0.1464054, 0.1464035, 0.146415, 0.1464105, 0.1464338, 0.1464238, 
    0.1464505, 0.1464441, 0.146452, 0.146448, 0.1464549, 0.1464487, 
    0.1464595, 0.1464618, 0.1464602, 0.1464665, 0.1464483, 0.1464552, 
    0.1464035, 0.1464037, 0.1464052, 0.1463989, 0.1463985, 0.146393, 
    0.146398, 0.1464001, 0.1464056, 0.1464088, 0.1464119, 0.1464186, 
    0.1464261, 0.1464367, 0.1464445, 0.1464497, 0.1464465, 0.1464493, 
    0.1464462, 0.1464447, 0.1464609, 0.1464518, 0.1464656, 0.1464648, 
    0.1464585, 0.1464649, 0.146404, 0.1464023, 0.1463962, 0.1464009, 
    0.1463924, 0.1463971, 0.1463998, 0.1464105, 0.1464129, 0.1464151, 
    0.1464194, 0.1464249, 0.1464346, 0.1464432, 0.1464511, 0.1464505, 
    0.1464507, 0.1464525, 0.1464481, 0.1464532, 0.146454, 0.1464518, 
    0.1464647, 0.146461, 0.1464648, 0.1464624, 0.1464028, 0.1464057, 
    0.1464041, 0.1464071, 0.146405, 0.1464142, 0.1464169, 0.1464301, 
    0.1464248, 0.1464334, 0.1464257, 0.146427, 0.1464334, 0.1464262, 
    0.1464426, 0.1464313, 0.1464525, 0.1464409, 0.1464532, 0.1464511, 
    0.1464547, 0.1464579, 0.1464621, 0.1464695, 0.1464678, 0.1464742, 
    0.1464101, 0.1464138, 0.1464136, 0.1464175, 0.1464204, 0.1464269, 
    0.1464371, 0.1464333, 0.1464404, 0.1464418, 0.1464311, 0.1464376, 
    0.1464164, 0.1464197, 0.1464178, 0.1464103, 0.146434, 0.1464218, 
    0.1464446, 0.1464379, 0.1464574, 0.1464476, 0.1464669, 0.1464749, 
    0.1464829, 0.1464918, 0.1464159, 0.1464134, 0.146418, 0.1464242, 
    0.1464303, 0.1464383, 0.1464392, 0.1464406, 0.1464446, 0.1464478, 
    0.146441, 0.1464486, 0.1464202, 0.1464352, 0.1464123, 0.146419, 
    0.1464239, 0.1464219, 0.1464329, 0.1464355, 0.1464459, 0.1464405, 
    0.1464728, 0.1464584, 0.146499, 0.1464875, 0.1464125, 0.146416, 0.146428, 
    0.1464223, 0.1464389, 0.1464429, 0.1464463, 0.1464505, 0.1464511, 
    0.1464536, 0.1464495, 0.1464534, 0.1464383, 0.1464451, 0.1464267, 
    0.1464311, 0.1464291, 0.1464269, 0.1464338, 0.1464411, 0.1464414, 
    0.1464437, 0.1464499, 0.146439, 0.1464743, 0.1464521, 0.1464198, 
    0.1464263, 0.1464274, 0.1464248, 0.1464425, 0.1464361, 0.1464535, 
    0.1464488, 0.1464566, 0.1464527, 0.1464521, 0.1464472, 0.1464441, 
    0.1464363, 0.1464301, 0.1464252, 0.1464264, 0.1464317, 0.1464416, 
    0.146451, 0.1464489, 0.146456, 0.1464377, 0.1464452, 0.1464423, 
    0.1464501, 0.1464332, 0.146447, 0.1464296, 0.1464311, 0.146436, 
    0.1464456, 0.146448, 0.1464503, 0.1464489, 0.1464418, 0.1464408, 
    0.1464359, 0.1464345, 0.1464308, 0.1464277, 0.1464305, 0.1464334, 
    0.1464419, 0.1464495, 0.1464579, 0.1464601, 0.1464695, 0.1464616, 
    0.1464744, 0.1464632, 0.1464829, 0.1464481, 0.1464632, 0.1464362, 
    0.1464392, 0.1464443, 0.1464564, 0.14645, 0.1464576, 0.1464407, 
    0.1464318, 0.1464297, 0.1464255, 0.1464298, 0.1464295, 0.1464336, 
    0.1464323, 0.1464422, 0.1464369, 0.1464521, 0.1464576, 0.1464735, 
    0.1464832, 0.1464933, 0.1464978, 0.1464991, 0.1464997,
  0.1561804, 0.1561888, 0.1561872, 0.156194, 0.1561903, 0.1561947, 0.1561822, 
    0.1561891, 0.1561847, 0.1561813, 0.156207, 0.1561943, 0.1562209, 
    0.1562126, 0.1562337, 0.1562195, 0.1562366, 0.1562334, 0.1562433, 
    0.1562405, 0.1562529, 0.1562447, 0.1562597, 0.156251, 0.1562523, 
    0.1562444, 0.156197, 0.1562053, 0.1561965, 0.1561977, 0.1561971, 
    0.1561903, 0.1561868, 0.1561799, 0.1561812, 0.1561863, 0.1561982, 
    0.1561942, 0.1562045, 0.1562043, 0.1562157, 0.1562105, 0.15623, 
    0.1562245, 0.1562406, 0.1562365, 0.1562404, 0.1562392, 0.1562404, 
    0.1562344, 0.156237, 0.1562318, 0.1562115, 0.1562174, 0.1561998, 
    0.1561891, 0.1561825, 0.1561776, 0.1561783, 0.1561796, 0.1561863, 
    0.1561928, 0.1561977, 0.156201, 0.1562043, 0.1562138, 0.1562192, 
    0.156231, 0.156229, 0.1562326, 0.1562361, 0.156242, 0.156241, 0.1562436, 
    0.1562326, 0.1562398, 0.1562278, 0.1562311, 0.1562046, 0.1561953, 
    0.156191, 0.1561875, 0.1561788, 0.1561848, 0.1561824, 0.1561882, 
    0.1561918, 0.15619, 0.1562011, 0.1561968, 0.1562195, 0.1562096, 
    0.1562357, 0.1562294, 0.1562372, 0.1562333, 0.15624, 0.156234, 0.1562445, 
    0.1562468, 0.1562453, 0.1562514, 0.1562336, 0.1562404, 0.1561899, 
    0.1561902, 0.1561916, 0.1561856, 0.1561852, 0.1561798, 0.1561847, 
    0.1561867, 0.156192, 0.1561951, 0.1561981, 0.1562046, 0.1562119, 
    0.1562223, 0.1562298, 0.1562349, 0.1562318, 0.1562346, 0.1562315, 
    0.1562301, 0.1562459, 0.156237, 0.1562505, 0.1562498, 0.1562436, 
    0.1562499, 0.1561904, 0.1561888, 0.1561829, 0.1561875, 0.1561792, 
    0.1561838, 0.1561864, 0.1561967, 0.1561991, 0.1562012, 0.1562054, 
    0.1562108, 0.1562203, 0.1562286, 0.1562364, 0.1562358, 0.156236, 
    0.1562377, 0.1562334, 0.1562384, 0.1562392, 0.156237, 0.1562497, 
    0.1562461, 0.1562498, 0.1562474, 0.1561893, 0.1561921, 0.1561906, 
    0.1561935, 0.1561914, 0.1562003, 0.156203, 0.1562158, 0.1562107, 
    0.156219, 0.1562116, 0.1562128, 0.156219, 0.156212, 0.156228, 0.1562169, 
    0.1562377, 0.1562264, 0.1562384, 0.1562363, 0.1562399, 0.156243, 
    0.1562471, 0.1562544, 0.1562528, 0.156259, 0.1561964, 0.1562, 0.1561997, 
    0.1562036, 0.1562064, 0.1562127, 0.1562227, 0.1562189, 0.1562259, 
    0.1562273, 0.1562167, 0.1562231, 0.1562025, 0.1562057, 0.1562038, 
    0.1561966, 0.1562197, 0.1562077, 0.1562299, 0.1562234, 0.1562425, 
    0.1562329, 0.1562518, 0.1562597, 0.1562676, 0.1562764, 0.156202, 
    0.1561996, 0.1562041, 0.1562101, 0.1562161, 0.1562238, 0.1562247, 
    0.1562261, 0.1562299, 0.1562331, 0.1562265, 0.1562339, 0.1562062, 
    0.1562207, 0.1561986, 0.1562051, 0.1562098, 0.1562078, 0.1562185, 
    0.156221, 0.1562312, 0.156226, 0.1562577, 0.1562435, 0.1562835, 
    0.1562722, 0.1561987, 0.1562021, 0.1562137, 0.1562082, 0.1562244, 
    0.1562283, 0.1562317, 0.1562358, 0.1562363, 0.1562387, 0.1562347, 
    0.1562386, 0.1562238, 0.1562304, 0.1562125, 0.1562168, 0.1562149, 
    0.1562127, 0.1562194, 0.1562265, 0.1562268, 0.1562291, 0.1562352, 
    0.1562245, 0.1562592, 0.1562374, 0.1562058, 0.1562121, 0.1562132, 
    0.1562107, 0.1562279, 0.1562217, 0.1562387, 0.1562341, 0.1562417, 
    0.1562379, 0.1562373, 0.1562325, 0.1562295, 0.1562219, 0.1562158, 
    0.1562111, 0.1562122, 0.1562174, 0.156227, 0.1562363, 0.1562342, 
    0.1562411, 0.1562232, 0.1562306, 0.1562277, 0.1562353, 0.1562188, 
    0.1562324, 0.1562153, 0.1562168, 0.1562215, 0.156231, 0.1562333, 
    0.1562355, 0.1562342, 0.1562273, 0.1562262, 0.1562214, 0.1562201, 
    0.1562165, 0.1562135, 0.1562162, 0.156219, 0.1562274, 0.1562348, 
    0.156243, 0.1562451, 0.1562544, 0.1562466, 0.1562593, 0.1562482, 
    0.1562676, 0.1562334, 0.1562482, 0.1562218, 0.1562247, 0.1562297, 
    0.1562416, 0.1562353, 0.1562427, 0.1562262, 0.1562175, 0.1562155, 
    0.1562113, 0.1562155, 0.1562152, 0.1562192, 0.156218, 0.1562276, 
    0.1562224, 0.1562373, 0.1562427, 0.1562583, 0.1562679, 0.1562779, 
    0.1562823, 0.1562837, 0.1562842,
  0.1699228, 0.1699293, 0.1699281, 0.1699333, 0.1699304, 0.1699338, 
    0.1699242, 0.1699295, 0.1699261, 0.1699235, 0.1699434, 0.1699335, 
    0.1699543, 0.1699478, 0.1699644, 0.1699532, 0.1699667, 0.1699642, 
    0.1699721, 0.1699698, 0.1699798, 0.1699731, 0.1699851, 0.1699782, 
    0.1699793, 0.1699729, 0.1699356, 0.1699421, 0.1699352, 0.1699362, 
    0.1699357, 0.1699305, 0.1699277, 0.1699224, 0.1699234, 0.1699273, 
    0.1699366, 0.1699335, 0.1699415, 0.1699413, 0.1699502, 0.1699462, 
    0.1699615, 0.1699571, 0.1699699, 0.1699667, 0.1699698, 0.1699688, 
    0.1699698, 0.169965, 0.169967, 0.1699629, 0.1699469, 0.1699515, 
    0.1699378, 0.1699295, 0.1699244, 0.1699207, 0.1699212, 0.1699222, 
    0.1699274, 0.1699324, 0.1699362, 0.1699387, 0.1699413, 0.1699487, 
    0.169953, 0.1699623, 0.1699607, 0.1699635, 0.1699664, 0.169971, 
    0.1699702, 0.1699723, 0.1699635, 0.1699693, 0.1699598, 0.1699624, 
    0.1699416, 0.1699343, 0.1699309, 0.1699283, 0.1699216, 0.1699262, 
    0.1699244, 0.1699288, 0.1699316, 0.1699302, 0.1699388, 0.1699354, 
    0.1699532, 0.1699455, 0.169966, 0.1699611, 0.1699672, 0.1699641, 
    0.1699694, 0.1699646, 0.169973, 0.1699748, 0.1699736, 0.1699785, 
    0.1699644, 0.1699697, 0.1699302, 0.1699304, 0.1699315, 0.1699268, 
    0.1699265, 0.1699224, 0.1699261, 0.1699276, 0.1699318, 0.1699342, 
    0.1699365, 0.1699416, 0.1699473, 0.1699554, 0.1699614, 0.1699654, 
    0.169963, 0.1699651, 0.1699627, 0.1699616, 0.1699741, 0.169967, 
    0.1699778, 0.1699772, 0.1699723, 0.1699773, 0.1699305, 0.1699293, 
    0.1699248, 0.1699283, 0.1699219, 0.1699254, 0.1699274, 0.1699354, 
    0.1699373, 0.1699389, 0.1699422, 0.1699464, 0.1699538, 0.1699604, 
    0.1699665, 0.1699661, 0.1699662, 0.1699676, 0.1699642, 0.1699681, 
    0.1699688, 0.1699671, 0.1699771, 0.1699743, 0.1699772, 0.1699753, 
    0.1699297, 0.1699319, 0.1699307, 0.1699329, 0.1699313, 0.1699382, 
    0.1699403, 0.1699503, 0.1699463, 0.1699528, 0.169947, 0.169948, 
    0.1699529, 0.1699473, 0.16996, 0.1699512, 0.1699676, 0.1699587, 
    0.1699682, 0.1699665, 0.1699693, 0.1699718, 0.1699751, 0.1699809, 
    0.1699796, 0.1699846, 0.1699351, 0.1699379, 0.1699378, 0.1699408, 
    0.169943, 0.1699479, 0.1699557, 0.1699528, 0.1699583, 0.1699594, 
    0.1699511, 0.1699561, 0.1699399, 0.1699424, 0.1699409, 0.1699353, 
    0.1699533, 0.169944, 0.1699615, 0.1699563, 0.1699715, 0.1699638, 
    0.1699788, 0.1699852, 0.1699915, 0.1699986, 0.1699395, 0.1699376, 
    0.1699411, 0.1699459, 0.1699505, 0.1699566, 0.1699573, 0.1699584, 
    0.1699615, 0.169964, 0.1699587, 0.1699646, 0.1699428, 0.1699542, 
    0.1699369, 0.1699419, 0.1699456, 0.1699441, 0.1699525, 0.1699544, 
    0.1699625, 0.1699583, 0.1699835, 0.1699723, 0.1700043, 0.1699952, 
    0.169937, 0.1699396, 0.1699487, 0.1699444, 0.1699571, 0.1699602, 
    0.1699628, 0.1699661, 0.1699665, 0.1699684, 0.1699652, 0.1699683, 
    0.1699566, 0.1699619, 0.1699478, 0.1699511, 0.1699496, 0.1699479, 
    0.1699532, 0.1699588, 0.169959, 0.1699608, 0.1699656, 0.1699571, 
    0.1699848, 0.1699674, 0.1699425, 0.1699474, 0.1699483, 0.1699463, 
    0.1699599, 0.1699549, 0.1699684, 0.1699648, 0.1699708, 0.1699678, 
    0.1699673, 0.1699635, 0.1699611, 0.1699551, 0.1699503, 0.1699466, 
    0.1699475, 0.1699516, 0.1699591, 0.1699665, 0.1699648, 0.1699703, 
    0.1699561, 0.169962, 0.1699597, 0.1699657, 0.1699527, 0.1699634, 
    0.1699499, 0.1699511, 0.1699548, 0.1699623, 0.1699641, 0.1699659, 
    0.1699648, 0.1699594, 0.1699585, 0.1699548, 0.1699537, 0.1699509, 
    0.1699485, 0.1699506, 0.1699529, 0.1699594, 0.1699653, 0.1699718, 
    0.1699735, 0.1699809, 0.1699747, 0.1699848, 0.169976, 0.1699915, 
    0.1699642, 0.169976, 0.169955, 0.1699573, 0.1699612, 0.1699707, 
    0.1699657, 0.1699716, 0.1699585, 0.1699517, 0.1699501, 0.1699468, 
    0.1699501, 0.1699499, 0.169953, 0.169952, 0.1699596, 0.1699555, 
    0.1699673, 0.1699716, 0.169984, 0.1699917, 0.1699998, 0.1700034, 
    0.1700045, 0.1700049,
  0.185219, 0.1852223, 0.1852217, 0.1852244, 0.1852229, 0.1852246, 0.1852197, 
    0.1852224, 0.1852207, 0.1852194, 0.1852295, 0.1852245, 0.1852352, 
    0.1852318, 0.1852406, 0.1852347, 0.1852418, 0.1852405, 0.1852447, 
    0.1852435, 0.1852488, 0.1852452, 0.1852517, 0.185248, 0.1852486, 
    0.1852451, 0.1852255, 0.1852289, 0.1852253, 0.1852258, 0.1852256, 
    0.1852229, 0.1852215, 0.1852188, 0.1852193, 0.1852213, 0.185226, 
    0.1852245, 0.1852286, 0.1852285, 0.1852331, 0.185231, 0.185239, 
    0.1852367, 0.1852435, 0.1852418, 0.1852434, 0.185243, 0.1852434, 
    0.1852409, 0.185242, 0.1852398, 0.1852314, 0.1852338, 0.1852267, 
    0.1852224, 0.1852198, 0.185218, 0.1852182, 0.1852187, 0.1852213, 
    0.1852239, 0.1852258, 0.1852272, 0.1852285, 0.1852323, 0.1852345, 
    0.1852395, 0.1852386, 0.1852401, 0.1852416, 0.1852441, 0.1852437, 
    0.1852448, 0.1852401, 0.1852432, 0.1852381, 0.1852395, 0.1852286, 
    0.1852249, 0.1852232, 0.1852218, 0.1852184, 0.1852207, 0.1852198, 
    0.1852221, 0.1852235, 0.1852228, 0.1852272, 0.1852255, 0.1852347, 
    0.1852306, 0.1852414, 0.1852388, 0.1852421, 0.1852404, 0.1852433, 
    0.1852407, 0.1852452, 0.1852462, 0.1852455, 0.1852482, 0.1852406, 
    0.1852434, 0.1852228, 0.1852229, 0.1852234, 0.185221, 0.1852209, 
    0.1852188, 0.1852207, 0.1852215, 0.1852236, 0.1852248, 0.185226, 
    0.1852286, 0.1852316, 0.1852358, 0.185239, 0.1852411, 0.1852398, 
    0.185241, 0.1852397, 0.1852391, 0.1852458, 0.185242, 0.1852478, 
    0.1852475, 0.1852448, 0.1852475, 0.185223, 0.1852223, 0.18522, 0.1852218, 
    0.1852186, 0.1852204, 0.1852214, 0.1852254, 0.1852264, 0.1852272, 
    0.1852289, 0.1852311, 0.185235, 0.1852385, 0.1852417, 0.1852415, 
    0.1852416, 0.1852423, 0.1852405, 0.1852426, 0.1852429, 0.185242, 
    0.1852474, 0.1852459, 0.1852475, 0.1852464, 0.1852225, 0.1852236, 
    0.185223, 0.1852241, 0.1852233, 0.1852269, 0.185228, 0.1852331, 
    0.1852311, 0.1852345, 0.1852314, 0.1852319, 0.1852345, 0.1852316, 
    0.1852382, 0.1852336, 0.1852423, 0.1852375, 0.1852426, 0.1852417, 
    0.1852432, 0.1852445, 0.1852463, 0.1852495, 0.1852487, 0.1852515, 
    0.1852253, 0.1852267, 0.1852266, 0.1852282, 0.1852293, 0.1852319, 
    0.185236, 0.1852344, 0.1852373, 0.1852379, 0.1852335, 0.1852362, 
    0.1852277, 0.185229, 0.1852283, 0.1852254, 0.1852347, 0.1852299, 
    0.185239, 0.1852363, 0.1852444, 0.1852403, 0.1852483, 0.1852518, 
    0.1852552, 0.1852592, 0.1852276, 0.1852266, 0.1852284, 0.1852308, 
    0.1852333, 0.1852365, 0.1852368, 0.1852374, 0.185239, 0.1852404, 
    0.1852376, 0.1852407, 0.1852293, 0.1852352, 0.1852262, 0.1852288, 
    0.1852307, 0.1852299, 0.1852343, 0.1852353, 0.1852396, 0.1852374, 
    0.1852509, 0.1852448, 0.1852623, 0.1852573, 0.1852262, 0.1852276, 
    0.1852323, 0.1852301, 0.1852367, 0.1852384, 0.1852397, 0.1852415, 
    0.1852417, 0.1852427, 0.185241, 0.1852427, 0.1852365, 0.1852392, 
    0.1852318, 0.1852336, 0.1852328, 0.1852319, 0.1852347, 0.1852376, 
    0.1852377, 0.1852387, 0.1852412, 0.1852367, 0.1852515, 0.1852422, 
    0.1852291, 0.1852316, 0.1852321, 0.1852311, 0.1852382, 0.1852356, 
    0.1852427, 0.1852408, 0.185244, 0.1852424, 0.1852421, 0.1852401, 
    0.1852388, 0.1852357, 0.1852332, 0.1852312, 0.1852317, 0.1852338, 
    0.1852378, 0.1852417, 0.1852408, 0.1852437, 0.1852362, 0.1852393, 
    0.1852381, 0.1852413, 0.1852344, 0.18524, 0.185233, 0.1852336, 0.1852355, 
    0.1852395, 0.1852404, 0.1852414, 0.1852408, 0.1852379, 0.1852375, 
    0.1852355, 0.1852349, 0.1852334, 0.1852322, 0.1852333, 0.1852345, 
    0.1852379, 0.1852411, 0.1852446, 0.1852455, 0.1852495, 0.1852461, 
    0.1852516, 0.1852468, 0.1852552, 0.1852405, 0.1852468, 0.1852356, 
    0.1852368, 0.1852389, 0.1852439, 0.1852413, 0.1852444, 0.1852375, 
    0.1852339, 0.185233, 0.1852313, 0.1852331, 0.1852329, 0.1852346, 
    0.185234, 0.185238, 0.1852359, 0.1852421, 0.1852444, 0.1852511, 
    0.1852553, 0.1852598, 0.1852618, 0.1852624, 0.1852626,
  0.1954509, 0.1954517, 0.1954516, 0.1954522, 0.1954519, 0.1954523, 
    0.1954511, 0.1954518, 0.1954513, 0.195451, 0.1954535, 0.1954523, 
    0.195455, 0.1954541, 0.1954563, 0.1954548, 0.1954567, 0.1954563, 
    0.1954574, 0.1954571, 0.1954586, 0.1954576, 0.1954594, 0.1954583, 
    0.1954585, 0.1954576, 0.1954525, 0.1954533, 0.1954525, 0.1954526, 
    0.1954525, 0.1954519, 0.1954515, 0.1954509, 0.195451, 0.1954515, 
    0.1954526, 0.1954522, 0.1954533, 0.1954532, 0.1954544, 0.1954539, 
    0.1954559, 0.1954553, 0.1954571, 0.1954567, 0.1954571, 0.195457, 
    0.1954571, 0.1954564, 0.1954567, 0.1954561, 0.195454, 0.1954546, 
    0.1954528, 0.1954518, 0.1954511, 0.1954507, 0.1954508, 0.1954509, 
    0.1954515, 0.1954521, 0.1954526, 0.1954529, 0.1954532, 0.1954542, 
    0.1954548, 0.1954561, 0.1954558, 0.1954562, 0.1954566, 0.1954573, 
    0.1954572, 0.1954575, 0.1954562, 0.195457, 0.1954557, 0.1954561, 
    0.1954533, 0.1954523, 0.1954519, 0.1954516, 0.1954508, 0.1954513, 
    0.1954511, 0.1954517, 0.195452, 0.1954518, 0.1954529, 0.1954525, 
    0.1954548, 0.1954538, 0.1954566, 0.1954559, 0.1954567, 0.1954563, 
    0.1954571, 0.1954564, 0.1954576, 0.1954578, 0.1954577, 0.1954584, 
    0.1954563, 0.1954571, 0.1954518, 0.1954519, 0.195452, 0.1954514, 
    0.1954514, 0.1954509, 0.1954513, 0.1954515, 0.195452, 0.1954523, 
    0.1954526, 0.1954533, 0.195454, 0.1954551, 0.1954559, 0.1954565, 
    0.1954561, 0.1954564, 0.1954561, 0.195456, 0.1954577, 0.1954567, 
    0.1954583, 0.1954582, 0.1954575, 0.1954582, 0.1954519, 0.1954517, 
    0.1954512, 0.1954516, 0.1954508, 0.1954513, 0.1954515, 0.1954525, 
    0.1954527, 0.1954529, 0.1954534, 0.1954539, 0.1954549, 0.1954558, 
    0.1954567, 0.1954566, 0.1954566, 0.1954568, 0.1954563, 0.1954569, 
    0.195457, 0.1954567, 0.1954582, 0.1954578, 0.1954582, 0.1954579, 
    0.1954518, 0.195452, 0.1954519, 0.1954522, 0.195452, 0.1954528, 
    0.1954531, 0.1954544, 0.1954539, 0.1954547, 0.195454, 0.1954541, 
    0.1954548, 0.195454, 0.1954557, 0.1954545, 0.1954568, 0.1954556, 
    0.1954569, 0.1954566, 0.195457, 0.1954574, 0.1954579, 0.1954587, 
    0.1954585, 0.1954593, 0.1954525, 0.1954528, 0.1954528, 0.1954532, 
    0.1954535, 0.1954541, 0.1954551, 0.1954547, 0.1954555, 0.1954556, 
    0.1954545, 0.1954552, 0.195453, 0.1954534, 0.1954532, 0.1954525, 
    0.1954548, 0.1954536, 0.1954559, 0.1954552, 0.1954574, 0.1954563, 
    0.1954584, 0.1954594, 0.1954603, 0.1954614, 0.195453, 0.1954528, 
    0.1954532, 0.1954538, 0.1954544, 0.1954553, 0.1954554, 0.1954555, 
    0.1954559, 0.1954563, 0.1954556, 0.1954564, 0.1954534, 0.1954549, 
    0.1954527, 0.1954533, 0.1954538, 0.1954536, 0.1954547, 0.195455, 
    0.1954561, 0.1954555, 0.1954591, 0.1954575, 0.1954623, 0.1954609, 
    0.1954527, 0.195453, 0.1954542, 0.1954536, 0.1954553, 0.1954558, 
    0.1954561, 0.1954566, 0.1954566, 0.1954569, 0.1954565, 0.1954569, 
    0.1954553, 0.195456, 0.1954541, 0.1954545, 0.1954543, 0.1954541, 
    0.1954548, 0.1954556, 0.1954556, 0.1954558, 0.1954565, 0.1954553, 
    0.1954593, 0.1954568, 0.1954534, 0.195454, 0.1954542, 0.1954539, 
    0.1954557, 0.195455, 0.1954569, 0.1954564, 0.1954572, 0.1954568, 
    0.1954568, 0.1954562, 0.1954559, 0.1954551, 0.1954544, 0.1954539, 
    0.195454, 0.1954546, 0.1954556, 0.1954566, 0.1954564, 0.1954572, 
    0.1954552, 0.195456, 0.1954557, 0.1954565, 0.1954547, 0.1954562, 
    0.1954544, 0.1954545, 0.195455, 0.1954561, 0.1954563, 0.1954566, 
    0.1954564, 0.1954556, 0.1954555, 0.195455, 0.1954549, 0.1954545, 
    0.1954542, 0.1954545, 0.1954548, 0.1954557, 0.1954565, 0.1954574, 
    0.1954577, 0.1954587, 0.1954578, 0.1954593, 0.195458, 0.1954603, 
    0.1954563, 0.195458, 0.1954551, 0.1954554, 0.1954559, 0.1954572, 
    0.1954565, 0.1954574, 0.1954555, 0.1954546, 0.1954544, 0.195454, 
    0.1954544, 0.1954544, 0.1954548, 0.1954546, 0.1954557, 0.1954551, 
    0.1954568, 0.1954574, 0.1954592, 0.1954604, 0.1954616, 0.1954622, 
    0.1954623, 0.1954624,
  0.1982629, 0.198263, 0.198263, 0.1982631, 0.198263, 0.1982631, 0.1982629, 
    0.198263, 0.198263, 0.1982629, 0.1982632, 0.1982631, 0.1982634, 
    0.1982633, 0.1982636, 0.1982634, 0.1982636, 0.1982636, 0.1982637, 
    0.1982637, 0.1982639, 0.1982637, 0.198264, 0.1982638, 0.1982639, 
    0.1982637, 0.1982631, 0.1982632, 0.1982631, 0.1982631, 0.1982631, 
    0.198263, 0.198263, 0.1982629, 0.1982629, 0.198263, 0.1982631, 0.1982631, 
    0.1982632, 0.1982632, 0.1982633, 0.1982633, 0.1982635, 0.1982634, 
    0.1982637, 0.1982636, 0.1982637, 0.1982636, 0.1982637, 0.1982636, 
    0.1982636, 0.1982635, 0.1982633, 0.1982633, 0.1982631, 0.198263, 
    0.1982629, 0.1982629, 0.1982629, 0.1982629, 0.198263, 0.198263, 
    0.1982631, 0.1982631, 0.1982632, 0.1982633, 0.1982634, 0.1982635, 
    0.1982635, 0.1982636, 0.1982636, 0.1982637, 0.1982637, 0.1982637, 
    0.1982636, 0.1982637, 0.1982635, 0.1982635, 0.1982632, 0.1982631, 
    0.198263, 0.198263, 0.1982629, 0.198263, 0.1982629, 0.198263, 0.198263, 
    0.198263, 0.1982631, 0.1982631, 0.1982634, 0.1982632, 0.1982636, 
    0.1982635, 0.1982636, 0.1982636, 0.1982637, 0.1982636, 0.1982637, 
    0.1982638, 0.1982637, 0.1982638, 0.1982636, 0.1982637, 0.198263, 
    0.198263, 0.198263, 0.198263, 0.198263, 0.1982629, 0.198263, 0.198263, 
    0.198263, 0.1982631, 0.1982631, 0.1982632, 0.1982633, 0.1982634, 
    0.1982635, 0.1982636, 0.1982635, 0.1982636, 0.1982635, 0.1982635, 
    0.1982637, 0.1982636, 0.1982638, 0.1982638, 0.1982637, 0.1982638, 
    0.198263, 0.198263, 0.1982629, 0.198263, 0.1982629, 0.1982629, 0.198263, 
    0.1982631, 0.1982631, 0.1982632, 0.1982632, 0.1982633, 0.1982634, 
    0.1982635, 0.1982636, 0.1982636, 0.1982636, 0.1982636, 0.1982636, 
    0.1982636, 0.1982636, 0.1982636, 0.1982638, 0.1982637, 0.1982638, 
    0.1982638, 0.198263, 0.198263, 0.198263, 0.198263, 0.198263, 0.1982631, 
    0.1982632, 0.1982633, 0.1982633, 0.1982634, 0.1982633, 0.1982633, 
    0.1982634, 0.1982633, 0.1982635, 0.1982633, 0.1982636, 0.1982635, 
    0.1982636, 0.1982636, 0.1982637, 0.1982637, 0.1982638, 0.1982639, 
    0.1982639, 0.198264, 0.1982631, 0.1982631, 0.1982631, 0.1982632, 
    0.1982632, 0.1982633, 0.1982634, 0.1982634, 0.1982635, 0.1982635, 
    0.1982633, 0.1982634, 0.1982632, 0.1982632, 0.1982632, 0.1982631, 
    0.1982634, 0.1982632, 0.1982635, 0.1982634, 0.1982637, 0.1982636, 
    0.1982638, 0.198264, 0.1982641, 0.1982642, 0.1982632, 0.1982631, 
    0.1982632, 0.1982633, 0.1982633, 0.1982634, 0.1982635, 0.1982635, 
    0.1982635, 0.1982636, 0.1982635, 0.1982636, 0.1982632, 0.1982634, 
    0.1982631, 0.1982632, 0.1982633, 0.1982632, 0.1982634, 0.1982634, 
    0.1982635, 0.1982635, 0.1982639, 0.1982637, 0.1982644, 0.1982642, 
    0.1982631, 0.1982632, 0.1982633, 0.1982632, 0.1982634, 0.1982635, 
    0.1982635, 0.1982636, 0.1982636, 0.1982636, 0.1982636, 0.1982636, 
    0.1982634, 0.1982635, 0.1982633, 0.1982633, 0.1982633, 0.1982633, 
    0.1982634, 0.1982635, 0.1982635, 0.1982635, 0.1982636, 0.1982634, 
    0.198264, 0.1982636, 0.1982632, 0.1982633, 0.1982633, 0.1982633, 
    0.1982635, 0.1982634, 0.1982636, 0.1982636, 0.1982637, 0.1982636, 
    0.1982636, 0.1982636, 0.1982635, 0.1982634, 0.1982633, 0.1982633, 
    0.1982633, 0.1982633, 0.1982635, 0.1982636, 0.1982636, 0.1982637, 
    0.1982634, 0.1982635, 0.1982635, 0.1982636, 0.1982634, 0.1982636, 
    0.1982633, 0.1982633, 0.1982634, 0.1982635, 0.1982636, 0.1982636, 
    0.1982636, 0.1982635, 0.1982635, 0.1982634, 0.1982634, 0.1982633, 
    0.1982633, 0.1982633, 0.1982634, 0.1982635, 0.1982636, 0.1982637, 
    0.1982637, 0.1982639, 0.1982638, 0.198264, 0.1982638, 0.1982641, 
    0.1982636, 0.1982638, 0.1982634, 0.1982635, 0.1982635, 0.1982637, 
    0.1982636, 0.1982637, 0.1982635, 0.1982633, 0.1982633, 0.1982633, 
    0.1982633, 0.1982633, 0.1982634, 0.1982634, 0.1982635, 0.1982634, 
    0.1982636, 0.1982637, 0.1982639, 0.1982641, 0.1982643, 0.1982643, 
    0.1982644, 0.1982644,
  0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985154, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985154, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985154, 0.1985154, 0.1985154, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985154, 0.1985153, 0.1985154, 0.1985154, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985154, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985154, 0.1985153, 0.1985154, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 0.1985153, 
    0.1985153, 0.1985153, 0.1985154, 0.1985154, 0.1985154, 0.1985154, 
    0.1985154, 0.1985154,
  0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 0.1985223, 
    0.1985223, 0.1985223,
  0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 0.1985224, 
    0.1985224, 0.1985224,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 U10 =
  8.601478, 8.601529, 8.60152, 8.60156, 8.601538, 8.601564, 8.601489, 
    8.60153, 8.601504, 8.601483, 8.601637, 8.601562, 8.60172, 8.601671, 
    8.601795, 8.601712, 8.601812, 8.601794, 8.601852, 8.601835, 8.601908, 
    8.60186, 8.601947, 8.601896, 8.601904, 8.601858, 8.601578, 8.601627, 
    8.601575, 8.601582, 8.601579, 8.601538, 8.601517, 8.601475, 8.601482, 
    8.601514, 8.601585, 8.601562, 8.601624, 8.601622, 8.601689, 8.601659, 
    8.601774, 8.601742, 8.601836, 8.601812, 8.601835, 8.601828, 8.601835, 
    8.6018, 8.601815, 8.601784, 8.601665, 8.601699, 8.601595, 8.60153, 
    8.60149, 8.601461, 8.601465, 8.601473, 8.601514, 8.601553, 8.601583, 
    8.601602, 8.601622, 8.601678, 8.601709, 8.60178, 8.601768, 8.601789, 
    8.60181, 8.601844, 8.601838, 8.601853, 8.601789, 8.601831, 8.601761, 
    8.60178, 8.601624, 8.601568, 8.601542, 8.601521, 8.601468, 8.601504, 
    8.60149, 8.601525, 8.601546, 8.601536, 8.601603, 8.601577, 8.601711, 
    8.601653, 8.601808, 8.60177, 8.601816, 8.601793, 8.601832, 8.601797, 
    8.601859, 8.601872, 8.601863, 8.601899, 8.601795, 8.601834, 8.601536, 
    8.601538, 8.601545, 8.601509, 8.601507, 8.601475, 8.601503, 8.601516, 
    8.601548, 8.601566, 8.601584, 8.601624, 8.601666, 8.601728, 8.601773, 
    8.601803, 8.601785, 8.601801, 8.601783, 8.601774, 8.601867, 8.601814, 
    8.601893, 8.60189, 8.601853, 8.60189, 8.601539, 8.601529, 8.601493, 
    8.601521, 8.601471, 8.601499, 8.601514, 8.601576, 8.601591, 8.601604, 
    8.601628, 8.601661, 8.601716, 8.601766, 8.601811, 8.601808, 8.60181, 
    8.601819, 8.601794, 8.601823, 8.601828, 8.601815, 8.601889, 8.601868, 
    8.60189, 8.601875, 8.601532, 8.601549, 8.60154, 8.601557, 8.601544, 
    8.601598, 8.601614, 8.60169, 8.60166, 8.601709, 8.601665, 8.601672, 
    8.601709, 8.601667, 8.601762, 8.601697, 8.601819, 8.601752, 8.601824, 
    8.601811, 8.601831, 8.601851, 8.601873, 8.601916, 8.601907, 8.601943, 
    8.601574, 8.601596, 8.601595, 8.601618, 8.601634, 8.601671, 8.60173, 
    8.601708, 8.60175, 8.601758, 8.601696, 8.601733, 8.60161, 8.601629, 
    8.601619, 8.601576, 8.601713, 8.601642, 8.601773, 8.601735, 8.601848, 
    8.60179, 8.601901, 8.601947, 8.601993, 8.602042, 8.601608, 8.601593, 
    8.601621, 8.601656, 8.601691, 8.601737, 8.601743, 8.601751, 8.601773, 
    8.601792, 8.601753, 8.601797, 8.601633, 8.601719, 8.601587, 8.601626, 
    8.601654, 8.601643, 8.601707, 8.601721, 8.601781, 8.60175, 8.601934, 
    8.601853, 8.602083, 8.602018, 8.601588, 8.601608, 8.601678, 8.601645, 
    8.601741, 8.601765, 8.601784, 8.601808, 8.60181, 8.601825, 8.601802, 
    8.601825, 8.601738, 8.601776, 8.601671, 8.601696, 8.601685, 8.601671, 
    8.601712, 8.601753, 8.601755, 8.601768, 8.601804, 8.601742, 8.601943, 
    8.601816, 8.60163, 8.601668, 8.601675, 8.60166, 8.601762, 8.601725, 
    8.601825, 8.601798, 8.601842, 8.60182, 8.601817, 8.601789, 8.601771, 
    8.601727, 8.60169, 8.601662, 8.601668, 8.6017, 8.601756, 8.60181, 
    8.601799, 8.601839, 8.601734, 8.601777, 8.60176, 8.601805, 8.601707, 
    8.601788, 8.601687, 8.601696, 8.601724, 8.60178, 8.601793, 8.601807, 
    8.601799, 8.601758, 8.601751, 8.601724, 8.601715, 8.601694, 8.601676, 
    8.601692, 8.601709, 8.601758, 8.601802, 8.601851, 8.601862, 8.601916, 
    8.601871, 8.601944, 8.601879, 8.601992, 8.601793, 8.60188, 8.601726, 
    8.601743, 8.601771, 8.601841, 8.601805, 8.601849, 8.601751, 8.6017, 
    8.601688, 8.601664, 8.601688, 8.601686, 8.60171, 8.601703, 8.60176, 
    8.601729, 8.601816, 8.601848, 8.601938, 8.601994, 8.602052, 8.602077, 
    8.602084, 8.602087 ;

 URBAN_AC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 URBAN_HEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 VOCFLXT =
  3.95534e-15, 3.955743e-15, 3.955667e-15, 3.955989e-15, 3.955813e-15, 
    3.956022e-15, 3.955425e-15, 3.955757e-15, 3.955547e-15, 3.955381e-15, 
    3.956604e-15, 3.956004e-15, 3.957262e-15, 3.956873e-15, 3.957862e-15, 
    3.957197e-15, 3.957998e-15, 3.957851e-15, 3.958313e-15, 3.958181e-15, 
    3.958757e-15, 3.958374e-15, 3.959069e-15, 3.95867e-15, 3.958729e-15, 
    3.958361e-15, 3.956132e-15, 3.956527e-15, 3.956107e-15, 3.956164e-15, 
    3.95614e-15, 3.955814e-15, 3.955645e-15, 3.955314e-15, 3.955376e-15, 
    3.955621e-15, 3.956189e-15, 3.956002e-15, 3.95649e-15, 3.956479e-15, 
    3.957019e-15, 3.956776e-15, 3.957691e-15, 3.957432e-15, 3.958187e-15, 
    3.957996e-15, 3.958176e-15, 3.958123e-15, 3.958177e-15, 3.957897e-15, 
    3.958017e-15, 3.957773e-15, 3.95682e-15, 3.957097e-15, 3.956267e-15, 
    3.955757e-15, 3.955438e-15, 3.955206e-15, 3.955239e-15, 3.9553e-15, 
    3.955623e-15, 3.955933e-15, 3.956167e-15, 3.956323e-15, 3.956478e-15, 
    3.956926e-15, 3.957181e-15, 3.957739e-15, 3.957645e-15, 3.95781e-15, 
    3.957977e-15, 3.958249e-15, 3.958205e-15, 3.958323e-15, 3.957811e-15, 
    3.958149e-15, 3.95759e-15, 3.957742e-15, 3.956493e-15, 3.956053e-15, 
    3.955844e-15, 3.955681e-15, 3.955264e-15, 3.95555e-15, 3.955436e-15, 
    3.955712e-15, 3.955884e-15, 3.9558e-15, 3.956327e-15, 3.956122e-15, 
    3.957196e-15, 3.956733e-15, 3.957958e-15, 3.957665e-15, 3.958029e-15, 
    3.957844e-15, 3.958158e-15, 3.957876e-15, 3.95837e-15, 3.958474e-15, 
    3.958402e-15, 3.958688e-15, 3.957859e-15, 3.958174e-15, 3.955797e-15, 
    3.95581e-15, 3.955876e-15, 3.955585e-15, 3.955569e-15, 3.955311e-15, 
    3.955543e-15, 3.95564e-15, 3.955896e-15, 3.956043e-15, 3.956184e-15, 
    3.956495e-15, 3.956839e-15, 3.957327e-15, 3.957684e-15, 3.957922e-15, 
    3.957778e-15, 3.957904e-15, 3.957761e-15, 3.957695e-15, 3.958433e-15, 
    3.958016e-15, 3.958647e-15, 3.958613e-15, 3.958325e-15, 3.958617e-15, 
    3.95582e-15, 3.955742e-15, 3.95546e-15, 3.95568e-15, 3.955283e-15, 
    3.955502e-15, 3.955626e-15, 3.95612e-15, 3.956235e-15, 3.956333e-15, 
    3.956534e-15, 3.956788e-15, 3.957233e-15, 3.957625e-15, 3.957988e-15, 
    3.957962e-15, 3.957971e-15, 3.958049e-15, 3.957852e-15, 3.958082e-15, 
    3.958118e-15, 3.958019e-15, 3.958608e-15, 3.95844e-15, 3.958612e-15, 
    3.958503e-15, 3.955768e-15, 3.955901e-15, 3.955829e-15, 3.955964e-15, 
    3.955866e-15, 3.956291e-15, 3.956418e-15, 3.957023e-15, 3.956781e-15, 
    3.957174e-15, 3.956823e-15, 3.956884e-15, 3.957175e-15, 3.956844e-15, 
    3.957598e-15, 3.957077e-15, 3.958052e-15, 3.957519e-15, 3.958085e-15, 
    3.957986e-15, 3.958152e-15, 3.958298e-15, 3.958487e-15, 3.958827e-15, 
    3.95875e-15, 3.959039e-15, 3.956103e-15, 3.956274e-15, 3.956263e-15, 
    3.956446e-15, 3.95658e-15, 3.956876e-15, 3.957347e-15, 3.957171e-15, 
    3.9575e-15, 3.957564e-15, 3.957069e-15, 3.957368e-15, 3.956392e-15, 
    3.956544e-15, 3.956457e-15, 3.956113e-15, 3.957205e-15, 3.956641e-15, 
    3.957689e-15, 3.957383e-15, 3.958277e-15, 3.957827e-15, 3.958705e-15, 
    3.959069e-15, 3.959436e-15, 3.959837e-15, 3.956372e-15, 3.956255e-15, 
    3.956469e-15, 3.956755e-15, 3.957036e-15, 3.957401e-15, 3.957441e-15, 
    3.957508e-15, 3.957688e-15, 3.957837e-15, 3.957524e-15, 3.957875e-15, 
    3.956569e-15, 3.957257e-15, 3.956207e-15, 3.956515e-15, 3.956741e-15, 
    3.956647e-15, 3.957153e-15, 3.957271e-15, 3.957747e-15, 3.957504e-15, 
    3.958975e-15, 3.958322e-15, 3.96016e-15, 3.959641e-15, 3.956213e-15, 
    3.956374e-15, 3.956927e-15, 3.956665e-15, 3.957428e-15, 3.957614e-15, 
    3.95777e-15, 3.957961e-15, 3.957985e-15, 3.958099e-15, 3.957912e-15, 
    3.958094e-15, 3.957402e-15, 3.957711e-15, 3.95687e-15, 3.957071e-15, 
    3.95698e-15, 3.956877e-15, 3.957196e-15, 3.957528e-15, 3.957543e-15, 
    3.957648e-15, 3.957931e-15, 3.957431e-15, 3.959044e-15, 3.958032e-15, 
    3.956549e-15, 3.956848e-15, 3.9569e-15, 3.956783e-15, 3.957595e-15, 
    3.957299e-15, 3.958098e-15, 3.957883e-15, 3.958237e-15, 3.95806e-15, 
    3.958034e-15, 3.95781e-15, 3.957668e-15, 3.957311e-15, 3.957024e-15, 
    3.956801e-15, 3.956853e-15, 3.957099e-15, 3.95755e-15, 3.957984e-15, 
    3.957888e-15, 3.95821e-15, 3.957372e-15, 3.957719e-15, 3.957582e-15, 
    3.95794e-15, 3.957165e-15, 3.9578e-15, 3.957e-15, 3.957072e-15, 
    3.957293e-15, 3.957737e-15, 3.957847e-15, 3.95795e-15, 3.957889e-15, 
    3.957563e-15, 3.957514e-15, 3.95729e-15, 3.957224e-15, 3.957057e-15, 
    3.956914e-15, 3.957043e-15, 3.957176e-15, 3.957567e-15, 3.957915e-15, 
    3.958299e-15, 3.958396e-15, 3.958825e-15, 3.958464e-15, 3.959048e-15, 
    3.958535e-15, 3.959433e-15, 3.957849e-15, 3.958536e-15, 3.957307e-15, 
    3.957441e-15, 3.957675e-15, 3.95823e-15, 3.957938e-15, 3.958284e-15, 
    3.957512e-15, 3.957103e-15, 3.957008e-15, 3.956813e-15, 3.957012e-15, 
    3.956997e-15, 3.957187e-15, 3.957126e-15, 3.95758e-15, 3.957336e-15, 
    3.958031e-15, 3.958283e-15, 3.959006e-15, 3.959445e-15, 3.959907e-15, 
    3.960106e-15, 3.960168e-15, 3.960193e-15 ;

 VOLR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WA =
  4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 4000, 
    4000, 4000 ;

 WASTEHEAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WF =
  9.833859, 9.881695, 9.872383, 9.911053, 9.889587, 9.914927, 9.843543, 
    9.883599, 9.858015, 9.838156, 9.986374, 9.912779, 10.06316, 10.01596, 
    10.13477, 10.05581, 10.15074, 10.13248, 10.18748, 10.1717, 10.24226, 
    10.19476, 10.27893, 10.2309, 10.23841, 10.1932, 9.927557, 9.977195, 
    9.924622, 9.931689, 9.928516, 9.890033, 9.870679, 9.830205, 9.837544, 
    9.867272, 9.934868, 9.911886, 9.969859, 9.968547, 10.03333, 10.00409, 
    10.11337, 10.08224, 10.17236, 10.14965, 10.1713, 10.16473, 10.17138, 
    10.13808, 10.15234, 10.12307, 10.00957, 10.04284, 9.943797, 9.884545, 
    9.845299, 9.817513, 9.821438, 9.828924, 9.867447, 9.903747, 9.931468, 
    9.95004, 9.968359, 10.02395, 10.05344, 10.11968, 10.1077, 10.12799, 
    10.14739, 10.18003, 10.17465, 10.18904, 10.12745, 10.16836, 10.10088, 
    10.11931, 9.973363, 9.918082, 9.89466, 9.874173, 9.824457, 9.858774, 
    9.845238, 9.877458, 9.897967, 9.887819, 9.950548, 9.926132, 10.05519, 
    9.999474, 10.14513, 10.11016, 10.15352, 10.13138, 10.16934, 10.13517, 
    10.1944, 10.20733, 10.19849, 10.23245, 10.13328, 10.1713, 9.887536, 
    9.889191, 9.896899, 9.863041, 9.86097, 9.830005, 9.857553, 9.869302, 
    9.899156, 9.916844, 9.933677, 9.970748, 10.01226, 10.07047, 10.11242, 
    10.1406, 10.12331, 10.13857, 10.12152, 10.11353, 10.20249, 10.15248, 
    10.22756, 10.2234, 10.18939, 10.22387, 9.890352, 9.880833, 9.847831, 
    9.873652, 9.826636, 9.852938, 9.868083, 9.926646, 9.939537, 9.951507, 
    9.975167, 10.00559, 10.05909, 10.10578, 10.14852, 10.14539, 10.14649, 
    10.15605, 10.13238, 10.15994, 10.16458, 10.15247, 10.22284, 10.20271, 
    10.22331, 10.2102, 9.883925, 9.89995, 9.89129, 9.90758, 9.896103, 
    9.947206, 9.962561, 10.0346, 10.00499, 10.05213, 10.00977, 10.01727, 
    10.05368, 10.01205, 10.10321, 10.04136, 10.15642, 10.09447, 10.16032, 
    10.14834, 10.16817, 10.18596, 10.20836, 10.24978, 10.24018, 10.27487, 
    9.923867, 9.944709, 9.942869, 9.964705, 9.980873, 10.01597, 10.07242, 
    10.05117, 10.0902, 10.09805, 10.03876, 10.07514, 9.95867, 9.977434, 
    9.966257, 9.925512, 10.05607, 9.988936, 10.11312, 10.07658, 10.18342, 
    10.13021, 10.2349, 10.27986, 10.3218, 10.37077, 9.956091, 9.941917, 
    9.967302, 10.0025, 10.03521, 10.07881, 10.08328, 10.09146, 10.11267, 
    10.13053, 10.09405, 10.13501, 9.981797, 10.06191, 9.936564, 9.974211, 
    10.00042, 9.988913, 10.04874, 10.06287, 10.12044, 10.09065, 10.26876, 
    10.18973, 10.40813, 10.34725, 9.936969, 9.95604, 10.0226, 9.990897, 
    10.08172, 10.10416, 10.12242, 10.14579, 10.14832, 10.16218, 10.13947, 
    10.16129, 10.0789, 10.11567, 10.01498, 10.03943, 10.02817, 10.01584, 
    10.05394, 10.09463, 10.09549, 10.10856, 10.14546, 10.08209, 10.27899, 
    10.15713, 9.976864, 10.01372, 10.01898, 10.00469, 10.10191, 10.06662, 
    10.16185, 10.13605, 10.17833, 10.15731, 10.15422, 10.12726, 10.1105, 
    10.06824, 10.03393, 10.00677, 10.01308, 10.04292, 10.09712, 10.14855, 
    10.13727, 10.17512, 10.07512, 10.11698, 10.10079, 10.14304, 10.05061, 
    10.1293, 10.03055, 10.03919, 10.06592, 10.11983, 10.13177, 10.14454, 
    10.13666, 10.0985, 10.09225, 10.06527, 10.05783, 10.03731, 10.02034, 
    10.03584, 10.05214, 10.09851, 10.14041, 10.18622, 10.19744, 10.25117, 
    10.20743, 10.27968, 10.21824, 10.32422, 10.13386, 10.21643, 10.06713, 
    10.08315, 10.11217, 10.1789, 10.14284, 10.18502, 10.092, 10.04396, 
    10.03154, 10.00842, 10.03207, 10.03015, 10.05281, 10.04552, 10.10005, 
    10.07074, 10.15414, 10.18469, 10.27124, 10.32401, 10.37759, 10.4013, 
    10.40852, 10.41154 ;

 WIND =
  8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 8.568267, 
    8.568267, 8.568267 ;

 WOODC =
  0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 0.03074508, 
    0.03074508, 0.03074508 ;

 WOODC_ALLOC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOODC_LOSS =
  1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 1.949842e-11, 
    1.949842e-11, 1.949842e-11, 1.949842e-11 ;

 WOOD_HARVESTC =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WOOD_HARVESTN =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 WTGQ =
  1.728758e-09, 1.708626e-09, 1.712501e-09, 1.696543e-09, 1.705356e-09, 
    1.694964e-09, 1.724636e-09, 1.707837e-09, 1.718521e-09, 1.726925e-09, 
    1.666452e-09, 1.695839e-09, 1.637036e-09, 1.654966e-09, 1.610681e-09, 
    1.639799e-09, 1.60494e-09, 1.611506e-09, 1.59191e-09, 1.597473e-09, 
    1.572943e-09, 1.589356e-09, 1.560532e-09, 1.576831e-09, 1.574258e-09, 
    1.589903e-09, 1.689837e-09, 1.670053e-09, 1.691025e-09, 1.68817e-09, 
    1.68945e-09, 1.705173e-09, 1.713215e-09, 1.730317e-09, 1.727186e-09, 
    1.714637e-09, 1.686889e-09, 1.696201e-09, 1.672935e-09, 1.673453e-09, 
    1.64831e-09, 1.659548e-09, 1.61845e-09, 1.629913e-09, 1.59724e-09, 
    1.605328e-09, 1.597618e-09, 1.599948e-09, 1.597588e-09, 1.609484e-09, 
    1.604365e-09, 1.614916e-09, 1.657431e-09, 1.644695e-09, 1.683302e-09, 
    1.707447e-09, 1.723892e-09, 1.735766e-09, 1.734077e-09, 1.730867e-09, 
    1.714564e-09, 1.699529e-09, 1.688257e-09, 1.680804e-09, 1.673528e-09, 
    1.651901e-09, 1.640689e-09, 1.616152e-09, 1.620523e-09, 1.613133e-09, 
    1.606137e-09, 1.594533e-09, 1.596431e-09, 1.591361e-09, 1.613327e-09, 
    1.598659e-09, 1.623024e-09, 1.616284e-09, 1.671562e-09, 1.693678e-09, 
    1.703267e-09, 1.711754e-09, 1.732781e-09, 1.718202e-09, 1.723918e-09, 
    1.710385e-09, 1.701902e-09, 1.706087e-09, 1.680601e-09, 1.690414e-09, 
    1.640029e-09, 1.661341e-09, 1.60695e-09, 1.619624e-09, 1.603942e-09, 
    1.611905e-09, 1.598312e-09, 1.610534e-09, 1.589483e-09, 1.584975e-09, 
    1.588053e-09, 1.576296e-09, 1.611218e-09, 1.597618e-09, 1.706204e-09, 
    1.70552e-09, 1.702341e-09, 1.71641e-09, 1.717279e-09, 1.730403e-09, 
    1.718715e-09, 1.713788e-09, 1.701413e-09, 1.694182e-09, 1.687367e-09, 
    1.672585e-09, 1.656394e-09, 1.634296e-09, 1.618796e-09, 1.608577e-09, 
    1.614827e-09, 1.609306e-09, 1.615481e-09, 1.618392e-09, 1.586661e-09, 
    1.604317e-09, 1.577976e-09, 1.57941e-09, 1.591241e-09, 1.579248e-09, 
    1.70504e-09, 1.708982e-09, 1.722819e-09, 1.71197e-09, 1.731846e-09, 
    1.720661e-09, 1.714299e-09, 1.690207e-09, 1.685009e-09, 1.68022e-09, 
    1.670843e-09, 1.658969e-09, 1.638561e-09, 1.621226e-09, 1.605732e-09, 
    1.606857e-09, 1.606461e-09, 1.603038e-09, 1.611544e-09, 1.601651e-09, 
    1.600003e-09, 1.604319e-09, 1.579602e-09, 1.586583e-09, 1.579441e-09, 
    1.583977e-09, 1.707699e-09, 1.701087e-09, 1.704653e-09, 1.697961e-09, 
    1.70267e-09, 1.681939e-09, 1.675826e-09, 1.647832e-09, 1.659201e-09, 
    1.641183e-09, 1.657352e-09, 1.654463e-09, 1.640602e-09, 1.65647e-09, 
    1.622172e-09, 1.64526e-09, 1.602905e-09, 1.625389e-09, 1.601518e-09, 
    1.605798e-09, 1.598724e-09, 1.592444e-09, 1.584614e-09, 1.570376e-09, 
    1.57365e-09, 1.561894e-09, 1.69133e-09, 1.682937e-09, 1.683672e-09, 
    1.674974e-09, 1.668601e-09, 1.654962e-09, 1.633567e-09, 1.641544e-09, 
    1.62696e-09, 1.624065e-09, 1.646246e-09, 1.632553e-09, 1.677368e-09, 
    1.669954e-09, 1.67436e-09, 1.690665e-09, 1.639698e-09, 1.665446e-09, 
    1.618543e-09, 1.632014e-09, 1.593336e-09, 1.61233e-09, 1.575458e-09, 
    1.560224e-09, 1.546161e-09, 1.530056e-09, 1.678393e-09, 1.684054e-09, 
    1.673946e-09, 1.660168e-09, 1.647595e-09, 1.631186e-09, 1.629526e-09, 
    1.626496e-09, 1.618703e-09, 1.61221e-09, 1.625541e-09, 1.610591e-09, 
    1.668244e-09, 1.637503e-09, 1.686205e-09, 1.671223e-09, 1.660974e-09, 
    1.665453e-09, 1.642461e-09, 1.637138e-09, 1.615874e-09, 1.626794e-09, 
    1.563955e-09, 1.591124e-09, 1.518023e-09, 1.537744e-09, 1.686042e-09, 
    1.678412e-09, 1.652415e-09, 1.664678e-09, 1.630102e-09, 1.621821e-09, 
    1.615152e-09, 1.606711e-09, 1.605805e-09, 1.600853e-09, 1.608985e-09, 
    1.601173e-09, 1.631151e-09, 1.617611e-09, 1.655344e-09, 1.645991e-09, 
    1.65028e-09, 1.655011e-09, 1.6405e-09, 1.625329e-09, 1.625008e-09, 
    1.620208e-09, 1.606838e-09, 1.629965e-09, 1.560518e-09, 1.602661e-09, 
    1.670175e-09, 1.65583e-09, 1.653802e-09, 1.659314e-09, 1.622647e-09, 
    1.635736e-09, 1.600973e-09, 1.610216e-09, 1.59513e-09, 1.602589e-09, 
    1.603693e-09, 1.613395e-09, 1.619497e-09, 1.635131e-09, 1.648086e-09, 
    1.658512e-09, 1.656075e-09, 1.644664e-09, 1.624411e-09, 1.605723e-09, 
    1.609779e-09, 1.596266e-09, 1.632559e-09, 1.617133e-09, 1.623059e-09, 
    1.607701e-09, 1.641757e-09, 1.612664e-09, 1.64937e-09, 1.646082e-09, 
    1.635998e-09, 1.616098e-09, 1.611763e-09, 1.607162e-09, 1.609998e-09, 
    1.623903e-09, 1.626205e-09, 1.636241e-09, 1.639035e-09, 1.646797e-09, 
    1.653282e-09, 1.647355e-09, 1.641178e-09, 1.623897e-09, 1.608646e-09, 
    1.592355e-09, 1.58842e-09, 1.569908e-09, 1.584943e-09, 1.56029e-09, 
    1.581199e-09, 1.545363e-09, 1.611011e-09, 1.581822e-09, 1.635542e-09, 
    1.629572e-09, 1.61889e-09, 1.594931e-09, 1.607773e-09, 1.592775e-09, 
    1.626296e-09, 1.644274e-09, 1.648993e-09, 1.657874e-09, 1.648791e-09, 
    1.649526e-09, 1.640923e-09, 1.643677e-09, 1.62333e-09, 1.634194e-09, 
    1.603721e-09, 1.592893e-09, 1.563118e-09, 1.545427e-09, 1.52784e-09, 
    1.520206e-09, 1.517897e-09, 1.516935e-09 ;

 W_SCALAR =
  0.6203898, 0.6220559, 0.6217321, 0.6230751, 0.6223302, 0.6232094, 
    0.6207277, 0.622122, 0.621232, 0.6205398, 0.6256785, 0.623135, 0.6283165, 
    0.6266972, 0.6307619, 0.6280646, 0.6313052, 0.6306841, 0.6325526, 
    0.6320176, 0.6344052, 0.6327995, 0.6356414, 0.6340219, 0.6342754, 
    0.6327465, 0.6236471, 0.625362, 0.6235455, 0.6237901, 0.6236804, 
    0.6223456, 0.6216727, 0.6202624, 0.6205184, 0.6215543, 0.6239001, 
    0.6231041, 0.6251095, 0.6250642, 0.6272941, 0.6262891, 0.6300327, 
    0.6289696, 0.6320398, 0.6312683, 0.6320036, 0.6317807, 0.6320065, 
    0.6308748, 0.6313598, 0.6303635, 0.6264774, 0.6276204, 0.6242091, 
    0.6221548, 0.6207889, 0.619819, 0.6199562, 0.6202176, 0.6215603, 
    0.6228218, 0.6237826, 0.624425, 0.6250577, 0.6269717, 0.6279837, 
    0.6302477, 0.6298392, 0.630531, 0.6311915, 0.6322998, 0.6321175, 
    0.6326056, 0.6305127, 0.6319039, 0.6296066, 0.6302353, 0.6252298, 
    0.6233189, 0.6225061, 0.6217943, 0.6200616, 0.6212584, 0.6207867, 
    0.6219087, 0.6226212, 0.6222688, 0.6244425, 0.6235978, 0.6280437, 
    0.62613, 0.6311145, 0.6299231, 0.6313999, 0.6306465, 0.6319372, 
    0.6307756, 0.6327872, 0.633225, 0.6329258, 0.6340744, 0.6307112, 
    0.6320037, 0.622259, 0.6223164, 0.6225842, 0.621407, 0.6213349, 
    0.6202554, 0.6212159, 0.6216249, 0.6226625, 0.623276, 0.623859, 
    0.6251401, 0.6265698, 0.628567, 0.6300004, 0.6309604, 0.6303717, 
    0.6308915, 0.6303105, 0.6300381, 0.6330609, 0.6313643, 0.6339093, 
    0.6337686, 0.6326172, 0.6337844, 0.6223568, 0.622026, 0.6208771, 
    0.6217763, 0.6201378, 0.6210551, 0.6215824, 0.6236154, 0.6240618, 
    0.6244756, 0.6252926, 0.6263405, 0.6281773, 0.6297739, 0.6312299, 
    0.6311232, 0.6311608, 0.6314859, 0.6306805, 0.6316181, 0.6317754, 
    0.6313641, 0.6337497, 0.6330685, 0.6337656, 0.6333221, 0.6221336, 
    0.62269, 0.6223893, 0.6229547, 0.6225564, 0.6243269, 0.6248574, 
    0.6273373, 0.6263199, 0.6279388, 0.6264845, 0.6267422, 0.6279917, 
    0.626563, 0.6296859, 0.6275694, 0.6314986, 0.6293874, 0.6316308, 
    0.6312236, 0.6318977, 0.6325011, 0.63326, 0.6346592, 0.6343353, 
    0.6355048, 0.6235194, 0.6242406, 0.624177, 0.6249315, 0.6254893, 
    0.6266976, 0.6286338, 0.627906, 0.6292419, 0.62951, 0.6274803, 0.6287268, 
    0.6247231, 0.6253706, 0.6249851, 0.6235763, 0.6280738, 0.6257671, 
    0.630024, 0.6287763, 0.6324151, 0.6306065, 0.634157, 0.6356725, 
    0.6370972, 0.6387606, 0.624634, 0.6241441, 0.6250212, 0.6262341, 
    0.6273586, 0.6288524, 0.6290051, 0.6292849, 0.6300091, 0.6306177, 
    0.6293733, 0.6307703, 0.6255208, 0.6282738, 0.6239589, 0.6252594, 
    0.6261626, 0.6257664, 0.6278228, 0.628307, 0.6302737, 0.6292573, 
    0.6352986, 0.6326286, 0.6400258, 0.6379623, 0.623973, 0.6246324, 
    0.6269255, 0.6258348, 0.6289521, 0.6297185, 0.6303413, 0.6311371, 
    0.631223, 0.6316943, 0.6309218, 0.6316637, 0.6288556, 0.6301111, 
    0.6266635, 0.6275033, 0.627117, 0.6266932, 0.6280009, 0.6293929, 
    0.6294226, 0.6298687, 0.6311253, 0.6289647, 0.6356429, 0.6315221, 
    0.6253511, 0.6266202, 0.6268013, 0.6263099, 0.6296417, 0.6284352, 
    0.6316828, 0.6308057, 0.6322424, 0.6315287, 0.6314236, 0.6305063, 
    0.629935, 0.6284906, 0.6273144, 0.6263812, 0.6265982, 0.6276232, 
    0.629478, 0.6312307, 0.630847, 0.6321333, 0.6287262, 0.6301558, 
    0.6296034, 0.6310433, 0.6278867, 0.6305752, 0.6271988, 0.6274951, 
    0.6284112, 0.6302527, 0.6306598, 0.6310944, 0.6308262, 0.6295251, 
    0.6293118, 0.628389, 0.6281341, 0.6274306, 0.6268478, 0.6273803, 
    0.6279392, 0.6295256, 0.6309539, 0.6325097, 0.6328902, 0.6347058, 
    0.6332281, 0.6356659, 0.6335937, 0.637179, 0.6307308, 0.6335325, 
    0.6284529, 0.6290009, 0.6299917, 0.6322616, 0.6310365, 0.6324692, 
    0.6293034, 0.6276586, 0.6272327, 0.6264379, 0.6272509, 0.6271847, 
    0.6279624, 0.6277125, 0.6295782, 0.6285763, 0.631421, 0.6324579, 
    0.6353823, 0.6371723, 0.6389922, 0.6397949, 0.6400391, 0.6401412,
  0.5451764, 0.547204, 0.5468099, 0.5484441, 0.5475377, 0.5486075, 0.5455876, 
    0.5472845, 0.5462013, 0.545359, 0.5516114, 0.5485169, 0.5548193, 
    0.5528501, 0.5577924, 0.5545131, 0.5584528, 0.5576977, 0.5599691, 
    0.5593187, 0.5622209, 0.5602691, 0.5637231, 0.5617549, 0.562063, 
    0.5602047, 0.5491399, 0.5512265, 0.5490162, 0.549314, 0.5491803, 
    0.5475565, 0.5467377, 0.5450212, 0.545333, 0.5465935, 0.5494478, 
    0.5484793, 0.5509188, 0.5508637, 0.553576, 0.5523536, 0.5569059, 
    0.5556132, 0.5593458, 0.5584079, 0.5593018, 0.5590308, 0.5593053, 
    0.5579295, 0.5585191, 0.557308, 0.5525827, 0.5539728, 0.5498236, 
    0.5473244, 0.5456621, 0.5444817, 0.5446486, 0.5449668, 0.5466009, 
    0.5481358, 0.5493047, 0.5500862, 0.5508559, 0.553184, 0.5544146, 
    0.5571672, 0.5566706, 0.5575117, 0.5583146, 0.5596619, 0.5594401, 
    0.5600335, 0.5574894, 0.5591807, 0.5563877, 0.5571521, 0.5510657, 
    0.5487406, 0.547752, 0.5468857, 0.544777, 0.5462335, 0.5456595, 
    0.5470247, 0.5478917, 0.5474629, 0.5501075, 0.5490799, 0.5544875, 
    0.5521603, 0.5582209, 0.5567725, 0.5585679, 0.5576519, 0.5592211, 
    0.5578089, 0.5602542, 0.5607863, 0.5604227, 0.5618187, 0.5577307, 
    0.5593019, 0.547451, 0.5475209, 0.5478467, 0.5464143, 0.5463266, 
    0.5450127, 0.5461818, 0.5466795, 0.5479419, 0.5486884, 0.5493977, 
    0.5509561, 0.5526952, 0.5551239, 0.5568665, 0.5580336, 0.557318, 
    0.5579498, 0.5572435, 0.5569124, 0.560587, 0.5585247, 0.561618, 
    0.5614469, 0.5600476, 0.5614662, 0.54757, 0.5471675, 0.5457695, 
    0.5468637, 0.5448696, 0.5459861, 0.5466279, 0.5491015, 0.5496444, 
    0.5501478, 0.5511416, 0.5524162, 0.55465, 0.5565912, 0.5583612, 
    0.5582316, 0.5582772, 0.5586725, 0.5576933, 0.5588332, 0.5590245, 
    0.5585244, 0.561424, 0.5605961, 0.5614433, 0.5609043, 0.5472983, 
    0.5479755, 0.5476096, 0.5482976, 0.547813, 0.549967, 0.5506123, 
    0.5536286, 0.5523912, 0.55436, 0.5525912, 0.5529048, 0.5544244, 
    0.5526868, 0.5564843, 0.5539109, 0.5586878, 0.5561215, 0.5588486, 
    0.5583535, 0.5591729, 0.5599065, 0.5608288, 0.5625295, 0.5621358, 
    0.563557, 0.5489845, 0.549862, 0.5497846, 0.5507024, 0.5513809, 
    0.5528505, 0.555205, 0.55432, 0.5559443, 0.5562703, 0.5538023, 0.5553181, 
    0.5504489, 0.5512366, 0.5507676, 0.5490538, 0.5545241, 0.5517189, 
    0.5568953, 0.5553782, 0.5598019, 0.5576035, 0.5619191, 0.5637609, 
    0.5654919, 0.5675131, 0.5503406, 0.5497445, 0.5508115, 0.5522869, 
    0.5536543, 0.5554708, 0.5556565, 0.5559966, 0.5568771, 0.5576171, 
    0.5561042, 0.5578025, 0.5514195, 0.5547674, 0.5495192, 0.5511014, 
    0.5521998, 0.5517179, 0.5542187, 0.5548077, 0.5571989, 0.5559631, 
    0.5633066, 0.5600616, 0.56905, 0.5665432, 0.5495363, 0.5503384, 
    0.5531277, 0.5518011, 0.5555919, 0.5565239, 0.557281, 0.5582485, 
    0.5583528, 0.5589257, 0.5579867, 0.5588886, 0.5554747, 0.5570011, 
    0.5528089, 0.5538303, 0.5533605, 0.5528451, 0.5544353, 0.5561281, 
    0.556164, 0.5567065, 0.5582346, 0.5556073, 0.5637254, 0.5587168, 
    0.5512128, 0.5527564, 0.5529765, 0.5523789, 0.5564305, 0.5549635, 
    0.5589117, 0.5578455, 0.5595921, 0.5587244, 0.5585967, 0.5574816, 
    0.556787, 0.5550308, 0.5536006, 0.5524656, 0.5527295, 0.5539761, 
    0.5562316, 0.5583623, 0.5578958, 0.5594594, 0.5553173, 0.5570555, 
    0.556384, 0.5581344, 0.5542965, 0.5575658, 0.5534599, 0.5538203, 
    0.5549344, 0.5571735, 0.5576681, 0.5581965, 0.5578705, 0.5562887, 
    0.5560293, 0.5549073, 0.5545974, 0.5537418, 0.5530331, 0.5536807, 
    0.5543604, 0.5562893, 0.5580258, 0.559917, 0.5603794, 0.5625862, 
    0.5607903, 0.5637532, 0.561235, 0.5655917, 0.5577548, 0.5611604, 
    0.554985, 0.5556513, 0.556856, 0.5596156, 0.5581262, 0.5598678, 
    0.5560192, 0.5540192, 0.5535012, 0.5525346, 0.5535232, 0.5534429, 
    0.5543885, 0.5540846, 0.5563533, 0.555135, 0.5585936, 0.559854, 
    0.5634081, 0.5655833, 0.5677942, 0.5687695, 0.5690662, 0.5691901,
  0.5138817, 0.5161299, 0.5156929, 0.5175053, 0.5165, 0.5176866, 0.5143375, 
    0.5162192, 0.515018, 0.514084, 0.5210195, 0.5175861, 0.5245802, 
    0.5223941, 0.5278819, 0.5242403, 0.5286155, 0.5277767, 0.5303, 0.5295774, 
    0.5328026, 0.5306334, 0.5344725, 0.5322846, 0.5326271, 0.5305619, 
    0.5182772, 0.5205923, 0.51814, 0.5184702, 0.518322, 0.5165209, 0.5156128, 
    0.5137096, 0.5140552, 0.5154529, 0.5186188, 0.5175443, 0.5202508, 
    0.5201897, 0.5231999, 0.5218431, 0.5268972, 0.5254616, 0.5296075, 
    0.5285655, 0.5295586, 0.5292575, 0.5295625, 0.5280342, 0.5286891, 
    0.5273438, 0.5220973, 0.5236403, 0.5190356, 0.5162635, 0.5144201, 
    0.5131115, 0.5132965, 0.5136493, 0.5154611, 0.5171633, 0.51846, 0.519327, 
    0.5201809, 0.5227649, 0.5241309, 0.5271875, 0.5266359, 0.5275701, 
    0.5284619, 0.5299587, 0.5297123, 0.5303717, 0.5275453, 0.5294241, 
    0.5263218, 0.5271707, 0.5204139, 0.5178342, 0.5167377, 0.5157769, 
    0.5134388, 0.5150537, 0.5144172, 0.5159311, 0.5168927, 0.5164171, 
    0.5193506, 0.5182106, 0.5242118, 0.5216285, 0.5283579, 0.5267491, 
    0.5287433, 0.5277259, 0.529469, 0.5279002, 0.5306169, 0.5312082, 
    0.5308042, 0.5323555, 0.5278133, 0.5295587, 0.5164038, 0.5164813, 
    0.5168427, 0.5152542, 0.5151569, 0.5137002, 0.5149963, 0.5155482, 
    0.5169483, 0.5177763, 0.5185631, 0.5202922, 0.5222222, 0.5249183, 
    0.5268534, 0.5281498, 0.5273549, 0.5280567, 0.5272722, 0.5269044, 
    0.5309867, 0.5286953, 0.5321324, 0.5319423, 0.5303873, 0.5319637, 
    0.5165358, 0.5160894, 0.5145392, 0.5157524, 0.5135415, 0.5147794, 
    0.515491, 0.5182346, 0.5188368, 0.5193954, 0.520498, 0.5219125, 
    0.5243922, 0.5265477, 0.5285137, 0.5283697, 0.5284204, 0.5288595, 
    0.5277718, 0.529038, 0.5292505, 0.5286949, 0.5319169, 0.5309968, 
    0.5319383, 0.5313392, 0.5162345, 0.5169855, 0.5165797, 0.5173428, 
    0.5168053, 0.5191947, 0.5199108, 0.5232583, 0.5218847, 0.5240702, 
    0.5221068, 0.5224548, 0.5241418, 0.5222129, 0.5264291, 0.5235716, 
    0.5288765, 0.5260261, 0.5290551, 0.5285052, 0.5294155, 0.5302305, 
    0.5312554, 0.5331456, 0.532708, 0.5342878, 0.5181047, 0.5190782, 
    0.5189924, 0.5200107, 0.5207636, 0.5223945, 0.5250084, 0.5240257, 
    0.5258294, 0.5261914, 0.523451, 0.525134, 0.5197294, 0.5206035, 0.520083, 
    0.5181816, 0.5242525, 0.5211387, 0.5268854, 0.5252007, 0.5301144, 
    0.5276721, 0.5324671, 0.5345145, 0.5364392, 0.5386873, 0.5196092, 
    0.5189479, 0.5201317, 0.521769, 0.5232868, 0.5253035, 0.5255097, 
    0.5258874, 0.5268652, 0.5276871, 0.5260069, 0.5278931, 0.5208065, 
    0.5245225, 0.518698, 0.5204534, 0.5216724, 0.5211376, 0.5239134, 
    0.5245672, 0.5272226, 0.5258502, 0.5340095, 0.5304029, 0.5403971, 
    0.5376084, 0.5187169, 0.5196068, 0.5227022, 0.5212299, 0.5254381, 
    0.5264729, 0.5273138, 0.5283884, 0.5285043, 0.5291408, 0.5280977, 
    0.5290995, 0.5253078, 0.5270029, 0.5223484, 0.5234821, 0.5229606, 
    0.5223885, 0.5241538, 0.5260334, 0.5260733, 0.5266758, 0.5283732, 
    0.5254551, 0.5344751, 0.5289088, 0.520577, 0.5222902, 0.5225345, 
    0.5218711, 0.5263692, 0.5247403, 0.5291253, 0.5279409, 0.5298811, 
    0.5289172, 0.5287753, 0.5275366, 0.5267652, 0.524815, 0.5232272, 
    0.5219673, 0.5222602, 0.5236441, 0.5261483, 0.5285149, 0.5279967, 
    0.5297337, 0.5251331, 0.5270634, 0.5263176, 0.5282617, 0.5239997, 
    0.5276303, 0.523071, 0.523471, 0.5247079, 0.5271944, 0.5277438, 
    0.5283308, 0.5279686, 0.5262118, 0.5259237, 0.5246778, 0.5243338, 
    0.5233839, 0.5225973, 0.523316, 0.5240707, 0.5262125, 0.5281411, 
    0.5302421, 0.530756, 0.5332087, 0.5312126, 0.5345061, 0.5317068, 
    0.5365502, 0.5278401, 0.531624, 0.5247641, 0.525504, 0.5268419, 
    0.5299073, 0.5282526, 0.5301875, 0.5259125, 0.523692, 0.5231168, 
    0.5220439, 0.5231413, 0.5230521, 0.5241018, 0.5237645, 0.5262835, 
    0.5249307, 0.5287718, 0.5301722, 0.5341223, 0.5365409, 0.539, 0.540085, 
    0.540415, 0.540553,
  0.5071226, 0.5095131, 0.5090484, 0.5109763, 0.5099068, 0.5111692, 
    0.5076072, 0.5096081, 0.5083308, 0.5073377, 0.5147167, 0.5110623, 
    0.5185099, 0.5161807, 0.5220302, 0.5181476, 0.5228127, 0.5219179, 
    0.5246101, 0.5238389, 0.5272819, 0.524966, 0.5290655, 0.5267287, 
    0.5270945, 0.5248896, 0.5117976, 0.5142619, 0.5116516, 0.5120031, 
    0.5118454, 0.509929, 0.5089633, 0.5069396, 0.5073071, 0.5087932, 
    0.5121611, 0.5110179, 0.5138983, 0.5138333, 0.5170391, 0.5155938, 
    0.5209799, 0.5194494, 0.5238711, 0.5227594, 0.523819, 0.5234976, 
    0.5238231, 0.5221926, 0.5228912, 0.5214562, 0.5158646, 0.5175084, 
    0.5126048, 0.5096553, 0.507695, 0.5063038, 0.5065005, 0.5068755, 
    0.5088019, 0.5106125, 0.5119921, 0.5129149, 0.5138239, 0.5165756, 
    0.5180311, 0.5212895, 0.5207013, 0.5216975, 0.5226488, 0.5242459, 
    0.523983, 0.5246866, 0.5216711, 0.5236754, 0.5203664, 0.5212716, 
    0.5140719, 0.5113263, 0.5101597, 0.5091377, 0.5066518, 0.5083687, 
    0.5076919, 0.5093017, 0.5103245, 0.5098186, 0.5129401, 0.5117267, 
    0.5181174, 0.5153653, 0.5225378, 0.520822, 0.522949, 0.5218637, 
    0.5237232, 0.5220497, 0.5249484, 0.5255795, 0.5251482, 0.5268044, 
    0.5219569, 0.523819, 0.5098045, 0.509887, 0.5102713, 0.5085819, 
    0.5084785, 0.5069296, 0.5083077, 0.5088946, 0.5103837, 0.5112646, 
    0.5121019, 0.5139424, 0.5159976, 0.5188703, 0.5209333, 0.5223159, 
    0.5214681, 0.5222166, 0.5213799, 0.5209876, 0.5253431, 0.5228978, 
    0.5265662, 0.5263633, 0.5247033, 0.5263861, 0.509945, 0.5094701, 
    0.5078216, 0.5091118, 0.506761, 0.508077, 0.5088337, 0.5117523, 
    0.5123932, 0.5129877, 0.5141615, 0.5156678, 0.5183096, 0.5206073, 
    0.5227041, 0.5225505, 0.5226045, 0.523073, 0.5219127, 0.5232635, 
    0.5234902, 0.5228974, 0.5263361, 0.5253538, 0.526359, 0.5257194, 
    0.5096244, 0.5104234, 0.5099916, 0.5108034, 0.5102316, 0.5127742, 
    0.5135363, 0.5171013, 0.5156382, 0.5179664, 0.5158747, 0.5162454, 
    0.5180427, 0.5159877, 0.5204808, 0.5174352, 0.5230912, 0.5200512, 
    0.5232816, 0.522695, 0.5236662, 0.524536, 0.5256299, 0.5276482, 
    0.5271809, 0.5288683, 0.5116141, 0.5126501, 0.5125588, 0.5136427, 
    0.5144443, 0.5161812, 0.5189664, 0.5179191, 0.5198414, 0.5202274, 
    0.5173067, 0.5191002, 0.5133433, 0.5142738, 0.5137197, 0.5116959, 
    0.5181606, 0.5148437, 0.5209674, 0.5191713, 0.524412, 0.5218064, 
    0.5269236, 0.5291106, 0.5311674, 0.5335712, 0.5132153, 0.5125114, 
    0.5137715, 0.5155149, 0.5171317, 0.5192809, 0.5195007, 0.5199033, 
    0.5209458, 0.5218223, 0.5200307, 0.522042, 0.5144899, 0.5184484, 
    0.5122454, 0.514114, 0.5154121, 0.5148425, 0.5177993, 0.5184961, 
    0.521327, 0.5198636, 0.528571, 0.5247199, 0.5354005, 0.5324174, 
    0.5122655, 0.5132128, 0.516509, 0.5149408, 0.5194243, 0.5205275, 
    0.5214242, 0.5225704, 0.5226941, 0.5233731, 0.5222604, 0.5233291, 
    0.5192855, 0.5210928, 0.5161321, 0.5173399, 0.5167842, 0.5161748, 
    0.5180555, 0.520059, 0.5201015, 0.5207438, 0.5225542, 0.5194424, 
    0.5290684, 0.5231256, 0.5142456, 0.51607, 0.5163302, 0.5156236, 0.520417, 
    0.5186806, 0.5233566, 0.522093, 0.5241631, 0.5231345, 0.5229832, 
    0.5216619, 0.5208392, 0.5187602, 0.5170682, 0.5157261, 0.5160382, 
    0.5175124, 0.5201815, 0.5227054, 0.5221526, 0.5240058, 0.5190993, 
    0.5211572, 0.520362, 0.5224353, 0.5178913, 0.5217618, 0.5169018, 
    0.517328, 0.5186461, 0.521297, 0.5218829, 0.522509, 0.5221226, 0.5202491, 
    0.519942, 0.518614, 0.5182474, 0.5172352, 0.5163971, 0.5171629, 0.517967, 
    0.5202498, 0.5223067, 0.5245484, 0.5250968, 0.5277157, 0.5255842, 
    0.5291016, 0.5261118, 0.5312861, 0.5219856, 0.5260233, 0.518706, 
    0.5194945, 0.520921, 0.524191, 0.5224255, 0.5244901, 0.51993, 0.5175634, 
    0.5169506, 0.5158077, 0.5169767, 0.5168816, 0.5180001, 0.5176407, 
    0.5203256, 0.5188835, 0.5229795, 0.5244737, 0.5286915, 0.5312761, 
    0.5339057, 0.5350664, 0.5354196, 0.5355673,
  0.5311409, 0.5336102, 0.5331299, 0.5351226, 0.534017, 0.5353221, 0.5316412, 
    0.5337083, 0.5323886, 0.531363, 0.5389929, 0.5352115, 0.5429235, 
    0.5405092, 0.5465765, 0.5425478, 0.5473893, 0.5464599, 0.549257, 
    0.5484555, 0.5520359, 0.549627, 0.5538929, 0.5514604, 0.5518409, 
    0.5495476, 0.5359719, 0.5385219, 0.535821, 0.5361845, 0.5360213, 0.53404, 
    0.533042, 0.530952, 0.5313313, 0.5328663, 0.5363479, 0.5351655, 
    0.5381456, 0.5380782, 0.5413987, 0.5399013, 0.5454862, 0.5438979, 
    0.5484889, 0.5473339, 0.5484347, 0.5481008, 0.5484391, 0.5467452, 
    0.5474709, 0.5459806, 0.5401817, 0.5418851, 0.536807, 0.5337571, 
    0.5317319, 0.5302957, 0.5304987, 0.5308858, 0.5328753, 0.5347465, 
    0.5361732, 0.5371278, 0.5380686, 0.5409184, 0.542427, 0.5458075, 
    0.545197, 0.5462311, 0.547219, 0.5488784, 0.5486052, 0.5493365, 
    0.5462037, 0.5482855, 0.5448493, 0.5457889, 0.5383253, 0.5354845, 
    0.5342784, 0.5332223, 0.5306548, 0.5324277, 0.5317287, 0.5333917, 
    0.5344488, 0.5339259, 0.5371539, 0.5358987, 0.5425165, 0.5396646, 
    0.5471038, 0.5453222, 0.5475308, 0.5464036, 0.5483353, 0.5465968, 
    0.5496086, 0.5502649, 0.5498164, 0.5515391, 0.5465004, 0.5484348, 
    0.5339113, 0.5339966, 0.5343938, 0.532648, 0.5325411, 0.5309417, 
    0.5323647, 0.532971, 0.53451, 0.5354208, 0.5362867, 0.5381913, 0.5403195, 
    0.5432972, 0.5454377, 0.5468733, 0.5459929, 0.5467702, 0.5459013, 
    0.5454941, 0.5500191, 0.5474777, 0.5512913, 0.5510802, 0.549354, 
    0.5511039, 0.5340564, 0.5335657, 0.5318627, 0.5331954, 0.5307675, 
    0.5321264, 0.5329081, 0.5359251, 0.536588, 0.5372031, 0.5384181, 
    0.5399778, 0.5427157, 0.5450993, 0.5472764, 0.5471168, 0.547173, 
    0.5476596, 0.5464545, 0.5478575, 0.5480931, 0.5474772, 0.5510519, 
    0.5500303, 0.5510756, 0.5504104, 0.5337252, 0.5345509, 0.5341047, 
    0.5349439, 0.5343527, 0.5369822, 0.5377709, 0.5414632, 0.5399472, 
    0.5423599, 0.5401922, 0.5405762, 0.542439, 0.5403092, 0.544968, 
    0.5418093, 0.5476785, 0.5445223, 0.5478764, 0.547267, 0.548276, 0.54918, 
    0.5503173, 0.5524172, 0.5519308, 0.5536874, 0.5357822, 0.5368538, 
    0.5367593, 0.537881, 0.5387108, 0.5405097, 0.5433968, 0.5423108, 
    0.5443046, 0.544705, 0.541676, 0.5435357, 0.5375711, 0.5385343, 
    0.5379606, 0.5358668, 0.5425613, 0.5391244, 0.5454732, 0.5436094, 
    0.5490511, 0.546344, 0.5516631, 0.5539398, 0.5560828, 0.5585898, 
    0.5374387, 0.5367104, 0.5380144, 0.5398195, 0.5414947, 0.5437231, 
    0.5439511, 0.5443688, 0.5454507, 0.5463607, 0.544501, 0.5465888, 
    0.5387581, 0.5428597, 0.5364352, 0.5383689, 0.539713, 0.5391232, 
    0.5421867, 0.5429091, 0.5458464, 0.5443276, 0.5533779, 0.5493712, 
    0.5604993, 0.5573862, 0.536456, 0.5374361, 0.5408493, 0.5392249, 
    0.5438718, 0.5450166, 0.5459473, 0.5471376, 0.547266, 0.5479715, 
    0.5468156, 0.5479257, 0.5437279, 0.5456032, 0.5404589, 0.5417104, 
    0.5411345, 0.5405031, 0.5424523, 0.5445303, 0.5445745, 0.5452411, 
    0.5471207, 0.5438907, 0.5538958, 0.5477143, 0.5385051, 0.5403945, 
    0.5406641, 0.5399321, 0.5449018, 0.5431004, 0.5479543, 0.5466418, 
    0.5487924, 0.5477236, 0.5475664, 0.5461941, 0.54534, 0.543183, 0.5414289, 
    0.5400383, 0.5403615, 0.5418893, 0.5446574, 0.5472778, 0.5467037, 
    0.5486289, 0.5435347, 0.5456702, 0.5448447, 0.5469972, 0.542282, 
    0.5462978, 0.5412564, 0.5416981, 0.5430647, 0.5458152, 0.5464236, 
    0.5470738, 0.5466725, 0.5447277, 0.544409, 0.5430314, 0.5426512, 
    0.5416019, 0.5407335, 0.541527, 0.5423605, 0.5447284, 0.5468636, 
    0.5491928, 0.549763, 0.5524874, 0.5502698, 0.5539303, 0.5508186, 
    0.5562065, 0.5465302, 0.5507265, 0.5431268, 0.5439447, 0.5454249, 
    0.5488214, 0.5469871, 0.5491322, 0.5443965, 0.5419421, 0.541307, 
    0.5401229, 0.541334, 0.5412355, 0.5423949, 0.5420222, 0.544807, 
    0.5433109, 0.5475625, 0.5491152, 0.5535034, 0.5561962, 0.5589388, 
    0.5601504, 0.5605193, 0.5606735,
  0.5352592, 0.5381025, 0.5375492, 0.5398464, 0.5385714, 0.5400766, 0.535835, 
    0.5382156, 0.5366953, 0.5355148, 0.5443175, 0.539949, 0.5488714, 
    0.5460728, 0.5531155, 0.5484356, 0.5540615, 0.5529799, 0.5562374, 
    0.5553032, 0.5594807, 0.5566688, 0.5616519, 0.5588083, 0.5592528, 
    0.5565763, 0.5408266, 0.5437729, 0.5406523, 0.5410719, 0.5408835, 
    0.5385979, 0.5374479, 0.535042, 0.5354784, 0.5372455, 0.5412607, 
    0.539896, 0.5433377, 0.5432599, 0.5471033, 0.5453688, 0.5518475, 
    0.5500024, 0.5553422, 0.553997, 0.555279, 0.5548901, 0.5552841, 
    0.5533118, 0.5541564, 0.5524224, 0.5456935, 0.5476671, 0.5417908, 
    0.5382718, 0.5359394, 0.5342872, 0.5345206, 0.5349658, 0.5372558, 
    0.5394126, 0.5410588, 0.5421613, 0.5432487, 0.5465468, 0.5482955, 
    0.5522211, 0.5515114, 0.5527138, 0.5538632, 0.555796, 0.5554776, 
    0.5563301, 0.5526819, 0.5551053, 0.5511074, 0.5521995, 0.5435454, 
    0.540264, 0.5388727, 0.5376555, 0.5347002, 0.5367404, 0.5359357, 
    0.5378507, 0.5390692, 0.5384664, 0.5421915, 0.540742, 0.5483992, 
    0.5450948, 0.5537291, 0.551657, 0.5542263, 0.5529145, 0.5551632, 
    0.5531392, 0.5566474, 0.5574129, 0.5568898, 0.5589003, 0.5530271, 
    0.5552791, 0.5384495, 0.5385479, 0.5390058, 0.536994, 0.536871, 
    0.5350301, 0.5366679, 0.537366, 0.5391398, 0.5401905, 0.5411899, 
    0.5433905, 0.5458531, 0.549305, 0.5517913, 0.5534609, 0.5524367, 
    0.5533409, 0.5523302, 0.5518568, 0.5571261, 0.5541644, 0.5586109, 
    0.5583644, 0.5563504, 0.5583922, 0.5386168, 0.5380512, 0.5360899, 
    0.5376245, 0.5348297, 0.5363935, 0.5372936, 0.5407724, 0.5415379, 
    0.5422484, 0.5436527, 0.5454575, 0.5486304, 0.5513979, 0.5539301, 
    0.5537444, 0.5538098, 0.5543762, 0.5529737, 0.5546067, 0.554881, 
    0.5541639, 0.5583314, 0.5571392, 0.5583591, 0.5575827, 0.5382351, 
    0.539187, 0.5386725, 0.5396402, 0.5389585, 0.5419931, 0.5429045, 
    0.547178, 0.545422, 0.5482177, 0.5457056, 0.5461504, 0.5483094, 
    0.5458412, 0.5512454, 0.5475791, 0.5543982, 0.5507275, 0.5546287, 
    0.5539191, 0.5550941, 0.5561476, 0.5574741, 0.5599262, 0.5593578, 
    0.5614114, 0.5406075, 0.5418449, 0.5417357, 0.5430318, 0.5439913, 
    0.5460733, 0.5494207, 0.5481607, 0.5504746, 0.5509398, 0.5474247, 
    0.5495818, 0.5426736, 0.5437872, 0.5431239, 0.5407051, 0.5484512, 
    0.5444697, 0.5518324, 0.5496675, 0.5559973, 0.5528452, 0.5590451, 
    0.5617067, 0.5642166, 0.5671582, 0.5425206, 0.5416791, 0.5431859, 
    0.5452742, 0.5472145, 0.5497994, 0.5500641, 0.5505492, 0.5518063, 
    0.5528646, 0.5507028, 0.5531299, 0.544046, 0.5487974, 0.5413614, 
    0.5435959, 0.5451509, 0.5444683, 0.5480168, 0.5488548, 0.5522664, 
    0.5505014, 0.5610493, 0.5563705, 0.5694026, 0.5657451, 0.5413854, 
    0.5425175, 0.5464667, 0.5445861, 0.5499721, 0.5513018, 0.5523837, 
    0.5537685, 0.553918, 0.5547394, 0.5533937, 0.5546861, 0.5498049, 
    0.5519837, 0.5460144, 0.5474645, 0.5467972, 0.5460657, 0.5483248, 
    0.5507368, 0.5507881, 0.5515627, 0.5537488, 0.5499939, 0.5616553, 
    0.5544398, 0.5437534, 0.54594, 0.5462523, 0.5454046, 0.5511684, 
    0.5490767, 0.5547193, 0.5531915, 0.5556958, 0.5544507, 0.5542676, 
    0.5526707, 0.5516776, 0.5491726, 0.5471383, 0.5455275, 0.5459018, 
    0.5476719, 0.5508845, 0.5539317, 0.5532635, 0.5555053, 0.5495807, 
    0.5520614, 0.5511021, 0.5536051, 0.5481274, 0.5527913, 0.5469384, 
    0.5474502, 0.5490352, 0.5522301, 0.5529377, 0.5536942, 0.5532272, 
    0.5509661, 0.5505959, 0.5489966, 0.5485556, 0.5473388, 0.5463325, 
    0.5472519, 0.5482184, 0.5509669, 0.5534497, 0.5561626, 0.5568274, 
    0.5600082, 0.5574186, 0.5616957, 0.558059, 0.5643616, 0.5530617, 
    0.5579516, 0.5491073, 0.5500568, 0.5517763, 0.5557296, 0.5535933, 
    0.556092, 0.5505814, 0.5477332, 0.546997, 0.5456254, 0.5470284, 
    0.5469142, 0.5482582, 0.5478261, 0.5510583, 0.5493209, 0.5542631, 
    0.5560721, 0.5611962, 0.5643494, 0.5675681, 0.5689924, 0.5694262, 
    0.5696076,
  0.5840976, 0.5875086, 0.5868437, 0.5896073, 0.5880724, 0.5898846, 
    0.5847872, 0.5876446, 0.5858188, 0.5844036, 0.5950114, 0.5897309, 
    0.6005509, 0.5971422, 0.6057471, 0.6000192, 0.6069097, 0.6055806, 
    0.6095905, 0.6084385, 0.613603, 0.610123, 0.6163005, 0.6127695, 
    0.6133204, 0.6100087, 0.5907891, 0.5943512, 0.5905789, 0.5910851, 
    0.5908578, 0.5881042, 0.5867221, 0.5838375, 0.58436, 0.5864791, 
    0.5913129, 0.589667, 0.5938241, 0.5937299, 0.5983957, 0.596287, 
    0.6041912, 0.6019324, 0.6084865, 0.6068304, 0.6084087, 0.6079295, 
    0.6084149, 0.6059882, 0.6070265, 0.6048962, 0.5966813, 0.5990824, 
    0.5919532, 0.5877121, 0.5849124, 0.5829344, 0.5832136, 0.5837463, 
    0.5864915, 0.5890847, 0.5910693, 0.5924011, 0.5937164, 0.5977185, 
    0.5998483, 0.6046493, 0.6037793, 0.6052538, 0.6066659, 0.609046, 
    0.6086534, 0.6097049, 0.6052146, 0.6081945, 0.6032844, 0.6046228, 
    0.5940757, 0.5901105, 0.5884349, 0.5869715, 0.5834284, 0.5858728, 
    0.5849079, 0.587206, 0.5886714, 0.5879461, 0.5924375, 0.590687, 
    0.5999748, 0.5959544, 0.606501, 0.6039577, 0.6071125, 0.6055002, 
    0.6082659, 0.6057761, 0.6100966, 0.6110424, 0.6103959, 0.6128834, 
    0.6056384, 0.6084088, 0.5879259, 0.588044, 0.5885951, 0.5861772, 
    0.5860295, 0.5838232, 0.5857859, 0.5866238, 0.5887564, 0.5900219, 
    0.5912276, 0.593888, 0.5968752, 0.6010803, 0.6041222, 0.6061714, 
    0.6049138, 0.6060239, 0.6047831, 0.6042026, 0.6106879, 0.6070363, 
    0.6125249, 0.6122196, 0.6097299, 0.612254, 0.5881271, 0.587447, 
    0.5850927, 0.5869343, 0.5835835, 0.5854568, 0.5865368, 0.5907238, 
    0.5916477, 0.5925063, 0.5942057, 0.5963947, 0.6002568, 0.6036403, 
    0.6067482, 0.6065198, 0.6066002, 0.6072969, 0.6055729, 0.6075805, 
    0.6079184, 0.6070357, 0.6121787, 0.6107041, 0.6122131, 0.6112524, 
    0.5876679, 0.5888132, 0.5881941, 0.5893589, 0.5885381, 0.5921977, 
    0.5932998, 0.5984868, 0.5963516, 0.5997534, 0.596696, 0.5972366, 
    0.5998653, 0.5968608, 0.6034534, 0.5989752, 0.6073241, 0.6028193, 
    0.6076077, 0.6067347, 0.6081808, 0.6094796, 0.6111181, 0.6141557, 
    0.6134506, 0.6160014, 0.5905248, 0.5920186, 0.5918867, 0.5934538, 
    0.5946159, 0.5971429, 0.6012216, 0.5996841, 0.60251, 0.6030792, 
    0.5987871, 0.6014184, 0.5930204, 0.5943686, 0.5935653, 0.5906426, 
    0.6000383, 0.5951958, 0.6041727, 0.601523, 0.6092943, 0.6054151, 
    0.613063, 0.6163687, 0.619499, 0.623184, 0.5928354, 0.5918184, 0.5936404, 
    0.5961721, 0.5985312, 0.6016843, 0.6020079, 0.6026012, 0.6041408, 
    0.6054389, 0.6027891, 0.6057648, 0.5946822, 0.6004606, 0.5914346, 
    0.5941368, 0.5960224, 0.5951942, 0.5995085, 0.6005306, 0.6047048, 
    0.6025427, 0.615551, 0.6097547, 0.6260078, 0.6214116, 0.5914636, 
    0.5928317, 0.5976212, 0.595337, 0.6018954, 0.6035225, 0.6048487, 
    0.6065495, 0.6067333, 0.607744, 0.6060889, 0.6076784, 0.6016911, 
    0.6043581, 0.5970713, 0.5988357, 0.5980232, 0.5971336, 0.5998841, 
    0.6028308, 0.6028935, 0.6038421, 0.6065252, 0.6019221, 0.6163048, 
    0.6073753, 0.5943276, 0.5969808, 0.5973604, 0.5963304, 0.6033591, 
    0.6008015, 0.6077192, 0.6058404, 0.6089224, 0.6073886, 0.6071634, 
    0.6052009, 0.603983, 0.6009186, 0.5984383, 0.5964796, 0.5969344, 
    0.5990883, 0.6030115, 0.6067501, 0.6059289, 0.6086875, 0.6014171, 
    0.6044534, 0.6032779, 0.6063486, 0.5996433, 0.6053489, 0.598195, 
    0.5988182, 0.6007509, 0.6046603, 0.6055287, 0.6064581, 0.6058843, 
    0.6031114, 0.6026583, 0.6007037, 0.6001655, 0.5986825, 0.5974579, 
    0.5985767, 0.5997543, 0.6031124, 0.6061576, 0.6094982, 0.6103189, 
    0.6142576, 0.6110495, 0.6163551, 0.6118417, 0.6196803, 0.6056809, 
    0.6117087, 0.6008388, 0.6019989, 0.604104, 0.6089641, 0.6063341, 
    0.609411, 0.6026406, 0.5991629, 0.5982664, 0.5965986, 0.5983046, 
    0.5981656, 0.5998029, 0.5992761, 0.6032243, 0.6010998, 0.6071578, 
    0.6093865, 0.6157336, 0.6196651, 0.623699, 0.6254908, 0.6260375, 0.6262662,
  0.6622251, 0.667787, 0.6666976, 0.6712429, 0.6687129, 0.6717016, 0.6633443, 
    0.6680101, 0.6650231, 0.6627214, 0.6802661, 0.6714472, 0.6897115, 
    0.6838751, 0.6987642, 0.6887959, 0.7008165, 0.6984711, 0.7055877, 
    0.7035307, 0.7128337, 0.7065421, 0.7177787, 0.711318, 0.7123192, 
    0.706337, 0.6732006, 0.679154, 0.6728517, 0.6736924, 0.6733148, 
    0.6687651, 0.6664985, 0.6618038, 0.6626507, 0.6661011, 0.6740712, 
    0.6713416, 0.6782681, 0.6781098, 0.6860123, 0.682423, 0.6960332, 
    0.6920996, 0.7036162, 0.7006762, 0.7034775, 0.7026251, 0.7034886, 
    0.6991889, 0.7010233, 0.6972684, 0.683092, 0.6871875, 0.6751375, 
    0.6681209, 0.6635476, 0.6603438, 0.6607947, 0.6616562, 0.6661214, 
    0.6703799, 0.6736662, 0.6758848, 0.6780871, 0.6848564, 0.688502, 
    0.6968355, 0.6953132, 0.6978964, 0.7003853, 0.7046142, 0.7039137, 
    0.7057924, 0.6978275, 0.7030964, 0.6944497, 0.696789, 0.6786907, 
    0.6720755, 0.669309, 0.6669068, 0.6611419, 0.6651114, 0.6635405, 
    0.6672908, 0.6696985, 0.6685052, 0.6759457, 0.6730312, 0.6887196, 
    0.6818596, 0.7000939, 0.6956249, 0.7011755, 0.6983296, 0.7032234, 
    0.6988153, 0.7064946, 0.7081949, 0.707032, 0.7115249, 0.6985729, 
    0.7034777, 0.6684719, 0.6686662, 0.6695728, 0.665608, 0.665367, 
    0.6617807, 0.6649695, 0.6663378, 0.6698384, 0.6719288, 0.6739292, 
    0.6783753, 0.6834213, 0.6906251, 0.6959125, 0.6995119, 0.6972994, 
    0.6992519, 0.6970701, 0.6960531, 0.7075568, 0.7010406, 0.7108743, 
    0.710321, 0.7058374, 0.7103833, 0.6688027, 0.6676859, 0.6638409, 
    0.6668458, 0.6613927, 0.6644333, 0.6661956, 0.6730922, 0.6746284, 
    0.6760606, 0.6789091, 0.6826057, 0.6892048, 0.6950704, 0.7005307, 
    0.7001271, 0.7002691, 0.7015024, 0.6984575, 0.7020053, 0.7026053, 
    0.7010396, 0.710247, 0.7075859, 0.7103093, 0.7085733, 0.6680484, 
    0.6699321, 0.6689128, 0.6708325, 0.6694789, 0.6755454, 0.6773884, 
    0.6861679, 0.6825325, 0.6883391, 0.683117, 0.6840357, 0.6885313, 
    0.6833967, 0.6947443, 0.6870038, 0.7015504, 0.6936398, 0.7020535, 
    0.7005069, 0.703072, 0.7053893, 0.7083312, 0.713842, 0.7125562, 
    0.7172273, 0.672762, 0.6752465, 0.6750265, 0.6776467, 0.6795995, 
    0.6838763, 0.6908692, 0.6882198, 0.6931019, 0.6940922, 0.6866817, 
    0.6912096, 0.6769205, 0.6791831, 0.6778337, 0.6729575, 0.6888287, 
    0.6805774, 0.6960008, 0.6913906, 0.7050577, 0.69818, 0.711851, 0.7179045, 
    0.7237219, 0.7306815, 0.6766108, 0.6749127, 0.6779597, 0.6822283, 
    0.6862438, 0.6916698, 0.6922304, 0.6932604, 0.6959449, 0.6982217, 
    0.6935872, 0.6987953, 0.6797112, 0.6895558, 0.6742736, 0.6787933, 
    0.6819748, 0.6805746, 0.6879184, 0.6896765, 0.6969327, 0.6931587, 
    0.7163987, 0.7058818, 0.7360995, 0.7273188, 0.6743218, 0.6766047, 
    0.6846905, 0.6808156, 0.6920354, 0.6948648, 0.6971852, 0.7001796, 
    0.7005044, 0.7022954, 0.6993665, 0.702179, 0.6916814, 0.6963252, 
    0.6837546, 0.6867649, 0.685376, 0.6838604, 0.6885635, 0.6936597, 
    0.6937689, 0.6954229, 0.7001367, 0.6920817, 0.7177866, 0.7016412, 
    0.6791143, 0.6836007, 0.6842464, 0.6824967, 0.6945799, 0.6901437, 
    0.7022516, 0.6989285, 0.7043934, 0.7016648, 0.7012656, 0.6978035, 
    0.6956691, 0.6903458, 0.6860851, 0.6827497, 0.6835218, 0.6871974, 
    0.6939742, 0.7005342, 0.6990844, 0.7039744, 0.6912072, 0.6964923, 
    0.6944383, 0.6998248, 0.6881498, 0.6980637, 0.6856694, 0.686735, 
    0.6900563, 0.6968548, 0.6983797, 0.7000182, 0.6990059, 0.6941482, 
    0.6933598, 0.689975, 0.6890477, 0.6865026, 0.6844125, 0.6863217, 
    0.6883404, 0.6941499, 0.6994876, 0.7054225, 0.7068936, 0.7140281, 
    0.7082077, 0.7178792, 0.7096372, 0.7240614, 0.6986477, 0.709397, 
    0.6902081, 0.6922148, 0.6958807, 0.7044679, 0.6997992, 0.7052665, 
    0.6933289, 0.6873254, 0.6857913, 0.6829515, 0.6858565, 0.6856191, 
    0.6884239, 0.6875196, 0.6943448, 0.6906587, 0.7012558, 0.7052227, 
    0.7167343, 0.7240329, 0.731664, 0.7351019, 0.7361569, 0.7365991,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 XSMRPOOL =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 XSMRPOOL_RECOVER =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZBOT =
  5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 
    5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5 ;

 ZWT =
  8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 8.801882, 
    8.801882, 8.801882 ;

 ZWT_CH4_UNSAT =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ZWT_PERCH =
  3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 3.801882, 
    3.801882, 3.801882 ;

 o2_decomp_depth_unsat =
  3.463412e-11, 3.47895e-11, 3.475921e-11, 3.488463e-11, 3.481502e-11, 
    3.489708e-11, 3.466544e-11, 3.479539e-11, 3.471238e-11, 3.464781e-11, 
    3.512799e-11, 3.488993e-11, 3.537605e-11, 3.522373e-11, 3.560661e-11, 
    3.53522e-11, 3.565795e-11, 3.559924e-11, 3.577601e-11, 3.572528e-11, 
    3.595148e-11, 3.57993e-11, 3.606896e-11, 3.591509e-11, 3.593907e-11, 
    3.579409e-11, 3.493813e-11, 3.509859e-11, 3.492854e-11, 3.495142e-11, 
    3.494112e-11, 3.481627e-11, 3.475338e-11, 3.462195e-11, 3.464575e-11, 
    3.474228e-11, 3.496143e-11, 3.488695e-11, 3.507467e-11, 3.507044e-11, 
    3.52797e-11, 3.518527e-11, 3.553768e-11, 3.543735e-11, 3.572736e-11, 
    3.565429e-11, 3.572384e-11, 3.570269e-11, 3.5724e-11, 3.561695e-11, 
    3.566272e-11, 3.556859e-11, 3.520339e-11, 3.531077e-11, 3.499057e-11, 
    3.479832e-11, 3.467096e-11, 3.458068e-11, 3.459335e-11, 3.461768e-11, 
    3.474276e-11, 3.486054e-11, 3.495039e-11, 3.501047e-11, 3.506971e-11, 
    3.524922e-11, 3.534444e-11, 3.555784e-11, 3.551933e-11, 3.558454e-11, 
    3.564699e-11, 3.575179e-11, 3.573451e-11, 3.578066e-11, 3.558265e-11, 
    3.571417e-11, 3.549706e-11, 3.555638e-11, 3.5086e-11, 3.490721e-11, 
    3.483112e-11, 3.476468e-11, 3.460313e-11, 3.471463e-11, 3.467061e-11, 
    3.477523e-11, 3.484175e-11, 3.480879e-11, 3.501207e-11, 3.493292e-11, 
    3.535002e-11, 3.517017e-11, 3.563974e-11, 3.552715e-11, 3.566663e-11, 
    3.559543e-11, 3.571737e-11, 3.560756e-11, 3.57978e-11, 3.583927e-11, 
    3.581084e-11, 3.591982e-11, 3.560123e-11, 3.572343e-11, 3.480808e-11, 
    3.481345e-11, 3.483842e-11, 3.472842e-11, 3.472169e-11, 3.462105e-11, 
    3.471052e-11, 3.474865e-11, 3.484552e-11, 3.490279e-11, 3.495728e-11, 
    3.50773e-11, 3.521138e-11, 3.539921e-11, 3.553439e-11, 3.562504e-11, 
    3.556941e-11, 3.561845e-11, 3.556354e-11, 3.553777e-11, 3.58236e-11, 
    3.566299e-11, 3.590403e-11, 3.589069e-11, 3.578145e-11, 3.589208e-11, 
    3.481715e-11, 3.478622e-11, 3.467901e-11, 3.476282e-11, 3.461003e-11, 
    3.469549e-11, 3.474458e-11, 3.493447e-11, 3.497625e-11, 3.501499e-11, 
    3.509153e-11, 3.518981e-11, 3.536248e-11, 3.551291e-11, 3.565047e-11, 
    3.564033e-11, 3.564386e-11, 3.567453e-11, 3.559838e-11, 3.568696e-11, 
    3.570177e-11, 3.566289e-11, 3.588879e-11, 3.58242e-11, 3.589025e-11, 
    3.584813e-11, 3.479621e-11, 3.484812e-11, 3.481998e-11, 3.48728e-11, 
    3.483549e-11, 3.500106e-11, 3.505069e-11, 3.528346e-11, 3.518786e-11, 
    3.534004e-11, 3.520325e-11, 3.522745e-11, 3.534478e-11, 3.521054e-11, 
    3.550444e-11, 3.530495e-11, 3.567568e-11, 3.547609e-11, 3.568811e-11, 
    3.564956e-11, 3.571327e-11, 3.577039e-11, 3.584223e-11, 3.597499e-11, 
    3.594416e-11, 3.605531e-11, 3.492561e-11, 3.499302e-11, 3.49871e-11, 
    3.505772e-11, 3.510995e-11, 3.522342e-11, 3.540552e-11, 3.533694e-11, 
    3.546275e-11, 3.548802e-11, 3.529677e-11, 3.541407e-11, 3.503783e-11, 
    3.509843e-11, 3.506232e-11, 3.493033e-11, 3.535235e-11, 3.513548e-11, 
    3.553616e-11, 3.541843e-11, 3.576213e-11, 3.559102e-11, 3.592721e-11, 
    3.607113e-11, 3.620686e-11, 3.636543e-11, 3.502986e-11, 3.498394e-11, 
    3.506606e-11, 3.517978e-11, 3.528542e-11, 3.542606e-11, 3.544043e-11, 
    3.546673e-11, 3.553502e-11, 3.55925e-11, 3.547493e-11, 3.560681e-11, 
    3.511237e-11, 3.537119e-11, 3.496606e-11, 3.508784e-11, 3.517255e-11, 
    3.51354e-11, 3.532863e-11, 3.537415e-11, 3.555949e-11, 3.546365e-11, 
    3.603544e-11, 3.578211e-11, 3.648639e-11, 3.628916e-11, 3.496786e-11, 
    3.502956e-11, 3.524464e-11, 3.514225e-11, 3.543537e-11, 3.550764e-11, 
    3.556636e-11, 3.564152e-11, 3.564959e-11, 3.569415e-11, 3.562105e-11, 
    3.569121e-11, 3.542594e-11, 3.554439e-11, 3.521966e-11, 3.529852e-11, 
    3.526221e-11, 3.522232e-11, 3.534524e-11, 3.547633e-11, 3.547915e-11, 
    3.552115e-11, 3.563958e-11, 3.543585e-11, 3.60679e-11, 3.567699e-11, 
    3.509689e-11, 3.521586e-11, 3.52329e-11, 3.518677e-11, 3.550028e-11, 
    3.538655e-11, 3.569307e-11, 3.56101e-11, 3.574595e-11, 3.56784e-11, 
    3.566838e-11, 3.55817e-11, 3.552765e-11, 3.539145e-11, 3.528067e-11, 
    3.519302e-11, 3.521331e-11, 3.530965e-11, 3.548426e-11, 3.564982e-11, 
    3.561347e-11, 3.573513e-11, 3.541329e-11, 3.55481e-11, 3.549587e-11, 
    3.563189e-11, 3.533495e-11, 3.558825e-11, 3.527022e-11, 3.529802e-11, 
    3.538419e-11, 3.555778e-11, 3.559623e-11, 3.563728e-11, 3.561189e-11, 
    3.5489e-11, 3.546886e-11, 3.538186e-11, 3.535778e-11, 3.529162e-11, 
    3.523675e-11, 3.528679e-11, 3.533927e-11, 3.548878e-11, 3.562357e-11, 
    3.577072e-11, 3.580678e-11, 3.597881e-11, 3.583859e-11, 3.606987e-11, 
    3.5873e-11, 3.621397e-11, 3.560293e-11, 3.586815e-11, 3.538814e-11, 
    3.543972e-11, 3.553307e-11, 3.574759e-11, 3.563172e-11, 3.576722e-11, 
    3.546805e-11, 3.5313e-11, 3.527297e-11, 3.519828e-11, 3.52746e-11, 
    3.52684e-11, 3.53415e-11, 3.531793e-11, 3.549363e-11, 3.53992e-11, 
    3.56676e-11, 3.576571e-11, 3.604319e-11, 3.621351e-11, 3.638728e-11, 
    3.646396e-11, 3.648732e-11, 3.649705e-11,
  1.775765e-11, 1.789211e-11, 1.786595e-11, 1.797461e-11, 1.791431e-11, 
    1.79855e-11, 1.778489e-11, 1.789745e-11, 1.782557e-11, 1.776975e-11, 
    1.818614e-11, 1.797947e-11, 1.840188e-11, 1.826937e-11, 1.860296e-11, 
    1.838122e-11, 1.86478e-11, 1.859658e-11, 1.875096e-11, 1.870669e-11, 
    1.890459e-11, 1.877141e-11, 1.900753e-11, 1.887277e-11, 1.889382e-11, 
    1.876702e-11, 1.802101e-11, 1.816035e-11, 1.801276e-11, 1.803261e-11, 
    1.802371e-11, 1.791555e-11, 1.786111e-11, 1.774741e-11, 1.776804e-11, 
    1.785157e-11, 1.804153e-11, 1.797698e-11, 1.813989e-11, 1.81362e-11, 
    1.831817e-11, 1.823604e-11, 1.854292e-11, 1.845552e-11, 1.870854e-11, 
    1.864478e-11, 1.870554e-11, 1.868711e-11, 1.870578e-11, 1.861231e-11, 
    1.865233e-11, 1.857017e-11, 1.825141e-11, 1.834487e-11, 1.806664e-11, 
    1.790006e-11, 1.778982e-11, 1.771172e-11, 1.772275e-11, 1.774379e-11, 
    1.785206e-11, 1.795411e-11, 1.803202e-11, 1.80842e-11, 1.813567e-11, 
    1.829173e-11, 1.83746e-11, 1.85606e-11, 1.852701e-11, 1.858395e-11, 
    1.863844e-11, 1.873003e-11, 1.871495e-11, 1.875534e-11, 1.858247e-11, 
    1.869728e-11, 1.850788e-11, 1.855961e-11, 1.814958e-11, 1.799439e-11, 
    1.79285e-11, 1.787097e-11, 1.773123e-11, 1.782769e-11, 1.778964e-11, 
    1.788023e-11, 1.793787e-11, 1.790935e-11, 1.808563e-11, 1.801702e-11, 
    1.837952e-11, 1.822305e-11, 1.863209e-11, 1.853391e-11, 1.865565e-11, 
    1.85935e-11, 1.870003e-11, 1.860414e-11, 1.877038e-11, 1.880664e-11, 
    1.878186e-11, 1.887716e-11, 1.859883e-11, 1.870552e-11, 1.790855e-11, 
    1.79132e-11, 1.793487e-11, 1.783968e-11, 1.783386e-11, 1.774684e-11, 
    1.782428e-11, 1.785728e-11, 1.794122e-11, 1.799091e-11, 1.803821e-11, 
    1.814237e-11, 1.825894e-11, 1.842245e-11, 1.854026e-11, 1.861939e-11, 
    1.857086e-11, 1.86137e-11, 1.856581e-11, 1.854338e-11, 1.879305e-11, 
    1.86527e-11, 1.886344e-11, 1.885176e-11, 1.875629e-11, 1.885308e-11, 
    1.791647e-11, 1.788972e-11, 1.779694e-11, 1.786953e-11, 1.773737e-11, 
    1.781129e-11, 1.785384e-11, 1.801843e-11, 1.805469e-11, 1.808831e-11, 
    1.81548e-11, 1.824024e-11, 1.839049e-11, 1.852161e-11, 1.864162e-11, 
    1.863282e-11, 1.863592e-11, 1.866275e-11, 1.859629e-11, 1.867367e-11, 
    1.868666e-11, 1.865269e-11, 1.88502e-11, 1.879369e-11, 1.885151e-11, 
    1.881472e-11, 1.789841e-11, 1.794344e-11, 1.79191e-11, 1.796487e-11, 
    1.793262e-11, 1.807619e-11, 1.811932e-11, 1.832168e-11, 1.823855e-11, 
    1.837094e-11, 1.825199e-11, 1.827304e-11, 1.837522e-11, 1.825842e-11, 
    1.851435e-11, 1.834066e-11, 1.86638e-11, 1.848978e-11, 1.867472e-11, 
    1.86411e-11, 1.869678e-11, 1.874669e-11, 1.880957e-11, 1.892575e-11, 
    1.889883e-11, 1.899616e-11, 1.801065e-11, 1.806919e-11, 1.806406e-11, 
    1.81254e-11, 1.817081e-11, 1.826941e-11, 1.842794e-11, 1.836828e-11, 
    1.847789e-11, 1.849992e-11, 1.833342e-11, 1.843557e-11, 1.810842e-11, 
    1.816111e-11, 1.812975e-11, 1.801526e-11, 1.838199e-11, 1.819343e-11, 
    1.854221e-11, 1.843964e-11, 1.873957e-11, 1.859017e-11, 1.888401e-11, 
    1.901008e-11, 1.91291e-11, 1.926843e-11, 1.810119e-11, 1.806138e-11, 
    1.813271e-11, 1.823152e-11, 1.832345e-11, 1.844589e-11, 1.845844e-11, 
    1.848141e-11, 1.854099e-11, 1.859113e-11, 1.848866e-11, 1.860371e-11, 
    1.81733e-11, 1.83984e-11, 1.804632e-11, 1.815205e-11, 1.82257e-11, 
    1.81934e-11, 1.836147e-11, 1.840116e-11, 1.856275e-11, 1.847916e-11, 
    1.897892e-11, 1.875721e-11, 1.937482e-11, 1.920149e-11, 1.804747e-11, 
    1.810106e-11, 1.828801e-11, 1.819898e-11, 1.845408e-11, 1.851707e-11, 
    1.856835e-11, 1.863394e-11, 1.864104e-11, 1.867996e-11, 1.861621e-11, 
    1.867744e-11, 1.844615e-11, 1.854938e-11, 1.826663e-11, 1.833529e-11, 
    1.83037e-11, 1.826906e-11, 1.837605e-11, 1.849027e-11, 1.849274e-11, 
    1.852942e-11, 1.863285e-11, 1.845512e-11, 1.900754e-11, 1.866562e-11, 
    1.815957e-11, 1.826304e-11, 1.827788e-11, 1.823775e-11, 1.851075e-11, 
    1.841165e-11, 1.867901e-11, 1.860662e-11, 1.872529e-11, 1.866629e-11, 
    1.865761e-11, 1.858194e-11, 1.853488e-11, 1.841619e-11, 1.831983e-11, 
    1.824357e-11, 1.82613e-11, 1.83451e-11, 1.849727e-11, 1.864167e-11, 
    1.861e-11, 1.871626e-11, 1.843554e-11, 1.855305e-11, 1.850759e-11, 
    1.862621e-11, 1.836668e-11, 1.858751e-11, 1.831039e-11, 1.833463e-11, 
    1.840969e-11, 1.856101e-11, 1.859459e-11, 1.863042e-11, 1.860832e-11, 
    1.850115e-11, 1.848362e-11, 1.840787e-11, 1.838696e-11, 1.832935e-11, 
    1.828169e-11, 1.832523e-11, 1.837098e-11, 1.85012e-11, 1.861883e-11, 
    1.87474e-11, 1.877892e-11, 1.892956e-11, 1.880686e-11, 1.900945e-11, 
    1.883709e-11, 1.913584e-11, 1.860038e-11, 1.883209e-11, 1.841312e-11, 
    1.84581e-11, 1.853952e-11, 1.872683e-11, 1.862566e-11, 1.874402e-11, 
    1.848294e-11, 1.834798e-11, 1.831316e-11, 1.82482e-11, 1.831465e-11, 
    1.830924e-11, 1.83729e-11, 1.835244e-11, 1.850553e-11, 1.842324e-11, 
    1.865738e-11, 1.874309e-11, 1.898594e-11, 1.913535e-11, 1.928792e-11, 
    1.93554e-11, 1.937596e-11, 1.938455e-11,
  1.677681e-11, 1.692557e-11, 1.689661e-11, 1.701692e-11, 1.695014e-11, 
    1.702898e-11, 1.680693e-11, 1.693149e-11, 1.685193e-11, 1.679019e-11, 
    1.725139e-11, 1.702229e-11, 1.749082e-11, 1.734369e-11, 1.771432e-11, 
    1.746788e-11, 1.77642e-11, 1.770721e-11, 1.7879e-11, 1.782971e-11, 
    1.805015e-11, 1.790176e-11, 1.816489e-11, 1.801468e-11, 1.803814e-11, 
    1.789687e-11, 1.706831e-11, 1.722279e-11, 1.705917e-11, 1.708116e-11, 
    1.70713e-11, 1.695151e-11, 1.689128e-11, 1.676547e-11, 1.678829e-11, 
    1.688071e-11, 1.709105e-11, 1.701954e-11, 1.720005e-11, 1.719597e-11, 
    1.739786e-11, 1.730671e-11, 1.764754e-11, 1.755039e-11, 1.783177e-11, 
    1.776083e-11, 1.782843e-11, 1.780792e-11, 1.78287e-11, 1.77247e-11, 
    1.776923e-11, 1.767784e-11, 1.732376e-11, 1.74275e-11, 1.711887e-11, 
    1.693439e-11, 1.681238e-11, 1.672602e-11, 1.673822e-11, 1.676148e-11, 
    1.688125e-11, 1.69942e-11, 1.70805e-11, 1.713832e-11, 1.719538e-11, 
    1.736854e-11, 1.746053e-11, 1.766721e-11, 1.762985e-11, 1.769317e-11, 
    1.775378e-11, 1.78557e-11, 1.783891e-11, 1.788387e-11, 1.769151e-11, 
    1.781925e-11, 1.760858e-11, 1.766609e-11, 1.721085e-11, 1.703882e-11, 
    1.696587e-11, 1.690218e-11, 1.67476e-11, 1.685428e-11, 1.681219e-11, 
    1.691241e-11, 1.697622e-11, 1.694465e-11, 1.71399e-11, 1.706388e-11, 
    1.746599e-11, 1.72923e-11, 1.77467e-11, 1.763752e-11, 1.777292e-11, 
    1.770377e-11, 1.782231e-11, 1.771561e-11, 1.790062e-11, 1.794101e-11, 
    1.79134e-11, 1.801955e-11, 1.770971e-11, 1.782842e-11, 1.694376e-11, 
    1.694891e-11, 1.69729e-11, 1.686755e-11, 1.686111e-11, 1.676485e-11, 
    1.68505e-11, 1.688702e-11, 1.697992e-11, 1.703497e-11, 1.708736e-11, 
    1.720281e-11, 1.733213e-11, 1.751366e-11, 1.764458e-11, 1.773257e-11, 
    1.76786e-11, 1.772625e-11, 1.767299e-11, 1.764805e-11, 1.792587e-11, 
    1.776964e-11, 1.800427e-11, 1.799126e-11, 1.788494e-11, 1.799272e-11, 
    1.695252e-11, 1.692291e-11, 1.682026e-11, 1.690057e-11, 1.675438e-11, 
    1.683614e-11, 1.688322e-11, 1.706545e-11, 1.710562e-11, 1.714288e-11, 
    1.721659e-11, 1.731137e-11, 1.747817e-11, 1.762386e-11, 1.775731e-11, 
    1.774752e-11, 1.775096e-11, 1.778082e-11, 1.770689e-11, 1.779297e-11, 
    1.780743e-11, 1.776963e-11, 1.798951e-11, 1.792658e-11, 1.799098e-11, 
    1.794999e-11, 1.693254e-11, 1.698239e-11, 1.695544e-11, 1.700613e-11, 
    1.697041e-11, 1.712946e-11, 1.717728e-11, 1.740176e-11, 1.73095e-11, 
    1.745645e-11, 1.73244e-11, 1.734777e-11, 1.746123e-11, 1.733153e-11, 
    1.76158e-11, 1.742284e-11, 1.778198e-11, 1.75885e-11, 1.779413e-11, 
    1.775673e-11, 1.781869e-11, 1.787424e-11, 1.794426e-11, 1.807372e-11, 
    1.804371e-11, 1.815221e-11, 1.705683e-11, 1.71217e-11, 1.7116e-11, 
    1.718399e-11, 1.723435e-11, 1.734373e-11, 1.751976e-11, 1.745348e-11, 
    1.757526e-11, 1.759974e-11, 1.741478e-11, 1.752823e-11, 1.716518e-11, 
    1.722361e-11, 1.718882e-11, 1.706194e-11, 1.746873e-11, 1.725945e-11, 
    1.764675e-11, 1.753275e-11, 1.786632e-11, 1.770009e-11, 1.802719e-11, 
    1.816776e-11, 1.830052e-11, 1.845612e-11, 1.715716e-11, 1.711303e-11, 
    1.719209e-11, 1.730171e-11, 1.740371e-11, 1.75397e-11, 1.755364e-11, 
    1.757917e-11, 1.764539e-11, 1.770114e-11, 1.758724e-11, 1.771513e-11, 
    1.723715e-11, 1.748695e-11, 1.709635e-11, 1.721356e-11, 1.729524e-11, 
    1.72594e-11, 1.744592e-11, 1.749e-11, 1.76696e-11, 1.757667e-11, 
    1.813301e-11, 1.788597e-11, 1.857499e-11, 1.838135e-11, 1.709762e-11, 
    1.715701e-11, 1.736439e-11, 1.726559e-11, 1.75488e-11, 1.76188e-11, 
    1.767581e-11, 1.774877e-11, 1.775667e-11, 1.779997e-11, 1.772903e-11, 
    1.779717e-11, 1.753999e-11, 1.765472e-11, 1.734064e-11, 1.741686e-11, 
    1.738178e-11, 1.734333e-11, 1.746212e-11, 1.758902e-11, 1.759176e-11, 
    1.763253e-11, 1.774762e-11, 1.754995e-11, 1.816497e-11, 1.778407e-11, 
    1.722188e-11, 1.733668e-11, 1.735313e-11, 1.73086e-11, 1.761178e-11, 
    1.750167e-11, 1.779891e-11, 1.771837e-11, 1.785042e-11, 1.778475e-11, 
    1.77751e-11, 1.769093e-11, 1.76386e-11, 1.75067e-11, 1.73997e-11, 
    1.731505e-11, 1.733472e-11, 1.742776e-11, 1.75968e-11, 1.775737e-11, 
    1.772214e-11, 1.784037e-11, 1.75282e-11, 1.76588e-11, 1.760827e-11, 
    1.774017e-11, 1.745172e-11, 1.769717e-11, 1.738921e-11, 1.741612e-11, 
    1.749948e-11, 1.766767e-11, 1.770499e-11, 1.774485e-11, 1.772026e-11, 
    1.760111e-11, 1.758163e-11, 1.749746e-11, 1.747424e-11, 1.741026e-11, 
    1.735736e-11, 1.740569e-11, 1.74565e-11, 1.760117e-11, 1.773196e-11, 
    1.787503e-11, 1.791013e-11, 1.807799e-11, 1.794127e-11, 1.816709e-11, 
    1.797499e-11, 1.830809e-11, 1.771146e-11, 1.796938e-11, 1.750329e-11, 
    1.755326e-11, 1.764377e-11, 1.785216e-11, 1.773955e-11, 1.787128e-11, 
    1.758087e-11, 1.743096e-11, 1.739229e-11, 1.732019e-11, 1.739394e-11, 
    1.738793e-11, 1.745861e-11, 1.743589e-11, 1.760598e-11, 1.751453e-11, 
    1.777485e-11, 1.787024e-11, 1.814082e-11, 1.830751e-11, 1.847787e-11, 
    1.855328e-11, 1.857626e-11, 1.858587e-11,
  1.72212e-11, 1.738502e-11, 1.735312e-11, 1.748567e-11, 1.741208e-11, 
    1.749897e-11, 1.725435e-11, 1.739153e-11, 1.73039e-11, 1.723592e-11, 
    1.774431e-11, 1.74916e-11, 1.80087e-11, 1.784616e-11, 1.825583e-11, 
    1.798336e-11, 1.831101e-11, 1.824795e-11, 1.843809e-11, 1.838352e-11, 
    1.862775e-11, 1.84633e-11, 1.875497e-11, 1.858841e-11, 1.861442e-11, 
    1.845789e-11, 1.754232e-11, 1.771275e-11, 1.753225e-11, 1.755649e-11, 
    1.754561e-11, 1.74136e-11, 1.734725e-11, 1.720871e-11, 1.723383e-11, 
    1.73356e-11, 1.75674e-11, 1.748855e-11, 1.768762e-11, 1.768311e-11, 
    1.790598e-11, 1.780533e-11, 1.818194e-11, 1.807452e-11, 1.83858e-11, 
    1.830727e-11, 1.83821e-11, 1.83594e-11, 1.83824e-11, 1.82673e-11, 
    1.831657e-11, 1.821545e-11, 1.782415e-11, 1.793872e-11, 1.759807e-11, 
    1.739475e-11, 1.726036e-11, 1.716529e-11, 1.717872e-11, 1.720432e-11, 
    1.733619e-11, 1.746063e-11, 1.755576e-11, 1.761952e-11, 1.768246e-11, 
    1.787362e-11, 1.797522e-11, 1.82037e-11, 1.816237e-11, 1.823242e-11, 
    1.829947e-11, 1.84123e-11, 1.83937e-11, 1.844349e-11, 1.823057e-11, 
    1.837195e-11, 1.813885e-11, 1.820246e-11, 1.769957e-11, 1.750981e-11, 
    1.742943e-11, 1.735924e-11, 1.718904e-11, 1.730649e-11, 1.726014e-11, 
    1.737051e-11, 1.744081e-11, 1.740603e-11, 1.762127e-11, 1.753744e-11, 
    1.798125e-11, 1.778943e-11, 1.829164e-11, 1.817085e-11, 1.832065e-11, 
    1.824414e-11, 1.837533e-11, 1.825724e-11, 1.846204e-11, 1.850678e-11, 
    1.84762e-11, 1.859381e-11, 1.82507e-11, 1.83821e-11, 1.740505e-11, 
    1.741072e-11, 1.743716e-11, 1.73211e-11, 1.731402e-11, 1.720802e-11, 
    1.730232e-11, 1.734255e-11, 1.744489e-11, 1.750556e-11, 1.756333e-11, 
    1.769066e-11, 1.78334e-11, 1.803393e-11, 1.817867e-11, 1.8276e-11, 
    1.821629e-11, 1.8269e-11, 1.821008e-11, 1.81825e-11, 1.849001e-11, 
    1.831703e-11, 1.857687e-11, 1.856245e-11, 1.844468e-11, 1.856407e-11, 
    1.741471e-11, 1.738208e-11, 1.726903e-11, 1.735747e-11, 1.71965e-11, 
    1.728651e-11, 1.733837e-11, 1.753918e-11, 1.758346e-11, 1.762455e-11, 
    1.770586e-11, 1.781047e-11, 1.79947e-11, 1.815575e-11, 1.830337e-11, 
    1.829254e-11, 1.829635e-11, 1.83294e-11, 1.824759e-11, 1.834285e-11, 
    1.835886e-11, 1.831701e-11, 1.856052e-11, 1.849079e-11, 1.856214e-11, 
    1.851673e-11, 1.739268e-11, 1.744761e-11, 1.741792e-11, 1.747378e-11, 
    1.743442e-11, 1.760976e-11, 1.76625e-11, 1.79103e-11, 1.780841e-11, 
    1.797071e-11, 1.782486e-11, 1.785066e-11, 1.797601e-11, 1.783273e-11, 
    1.814685e-11, 1.793359e-11, 1.833068e-11, 1.811667e-11, 1.834414e-11, 
    1.830273e-11, 1.837131e-11, 1.843283e-11, 1.851038e-11, 1.865386e-11, 
    1.862059e-11, 1.874089e-11, 1.752966e-11, 1.76012e-11, 1.75949e-11, 
    1.76699e-11, 1.772547e-11, 1.78462e-11, 1.804067e-11, 1.796742e-11, 
    1.8102e-11, 1.812908e-11, 1.792466e-11, 1.805003e-11, 1.764915e-11, 
    1.771362e-11, 1.767523e-11, 1.75353e-11, 1.798428e-11, 1.775317e-11, 
    1.818106e-11, 1.805502e-11, 1.842405e-11, 1.824007e-11, 1.860228e-11, 
    1.875816e-11, 1.890546e-11, 1.907827e-11, 1.76403e-11, 1.759163e-11, 
    1.767883e-11, 1.779982e-11, 1.791244e-11, 1.80627e-11, 1.807811e-11, 
    1.810634e-11, 1.817956e-11, 1.824123e-11, 1.811526e-11, 1.82567e-11, 
    1.772858e-11, 1.800441e-11, 1.757324e-11, 1.770254e-11, 1.779268e-11, 
    1.775311e-11, 1.795906e-11, 1.800777e-11, 1.820634e-11, 1.810356e-11, 
    1.871962e-11, 1.844584e-11, 1.921037e-11, 1.899521e-11, 1.757464e-11, 
    1.764014e-11, 1.786902e-11, 1.775994e-11, 1.807275e-11, 1.815015e-11, 
    1.82132e-11, 1.829394e-11, 1.830266e-11, 1.835059e-11, 1.827209e-11, 
    1.834749e-11, 1.806302e-11, 1.818988e-11, 1.784279e-11, 1.792697e-11, 
    1.788822e-11, 1.784576e-11, 1.797696e-11, 1.811724e-11, 1.812025e-11, 
    1.816535e-11, 1.82927e-11, 1.807403e-11, 1.875509e-11, 1.833304e-11, 
    1.77117e-11, 1.783843e-11, 1.785658e-11, 1.780741e-11, 1.814239e-11, 
    1.802066e-11, 1.834943e-11, 1.826029e-11, 1.840645e-11, 1.833375e-11, 
    1.832307e-11, 1.822992e-11, 1.817205e-11, 1.802624e-11, 1.790801e-11, 
    1.781454e-11, 1.783625e-11, 1.793901e-11, 1.812584e-11, 1.830345e-11, 
    1.826448e-11, 1.839532e-11, 1.804998e-11, 1.81944e-11, 1.813852e-11, 
    1.828441e-11, 1.796548e-11, 1.823688e-11, 1.789642e-11, 1.792614e-11, 
    1.801825e-11, 1.820421e-11, 1.824549e-11, 1.82896e-11, 1.826238e-11, 
    1.81306e-11, 1.810905e-11, 1.801601e-11, 1.799036e-11, 1.791967e-11, 
    1.786125e-11, 1.791462e-11, 1.797076e-11, 1.813065e-11, 1.827533e-11, 
    1.843371e-11, 1.847257e-11, 1.865862e-11, 1.850709e-11, 1.875745e-11, 
    1.854448e-11, 1.89139e-11, 1.825268e-11, 1.853825e-11, 1.802245e-11, 
    1.807768e-11, 1.817778e-11, 1.840839e-11, 1.828372e-11, 1.842956e-11, 
    1.810821e-11, 1.794255e-11, 1.789982e-11, 1.782021e-11, 1.790164e-11, 
    1.789501e-11, 1.797309e-11, 1.794798e-11, 1.813598e-11, 1.803488e-11, 
    1.832279e-11, 1.842841e-11, 1.872826e-11, 1.891323e-11, 1.910242e-11, 
    1.918623e-11, 1.921177e-11, 1.922246e-11,
  1.879542e-11, 1.897096e-11, 1.893676e-11, 1.907888e-11, 1.899996e-11, 
    1.909314e-11, 1.883093e-11, 1.897795e-11, 1.888402e-11, 1.881118e-11, 
    1.935645e-11, 1.908524e-11, 1.964049e-11, 1.94658e-11, 1.990635e-11, 
    1.961326e-11, 1.996576e-11, 1.989786e-11, 2.010262e-11, 2.004384e-11, 
    2.030709e-11, 2.012979e-11, 2.044433e-11, 2.026466e-11, 2.029271e-11, 
    2.012395e-11, 1.913963e-11, 1.932256e-11, 1.912883e-11, 1.915484e-11, 
    1.914316e-11, 1.900159e-11, 1.893048e-11, 1.878204e-11, 1.880894e-11, 
    1.891799e-11, 1.916655e-11, 1.908196e-11, 1.929554e-11, 1.929071e-11, 
    1.953008e-11, 1.942194e-11, 1.982682e-11, 1.971125e-11, 2.004629e-11, 
    1.996172e-11, 2.004231e-11, 2.001785e-11, 2.004263e-11, 1.991869e-11, 
    1.997174e-11, 1.986288e-11, 1.944216e-11, 1.956527e-11, 1.919945e-11, 
    1.898141e-11, 1.883736e-11, 1.873554e-11, 1.874991e-11, 1.877734e-11, 
    1.891863e-11, 1.905202e-11, 1.915404e-11, 1.922246e-11, 1.929001e-11, 
    1.949533e-11, 1.960451e-11, 1.985024e-11, 1.980576e-11, 1.988115e-11, 
    1.995332e-11, 2.007484e-11, 2.005481e-11, 2.010845e-11, 1.987915e-11, 
    2.003138e-11, 1.978045e-11, 1.98489e-11, 1.930842e-11, 1.910476e-11, 
    1.901859e-11, 1.894333e-11, 1.876097e-11, 1.888679e-11, 1.883714e-11, 
    1.89554e-11, 1.903077e-11, 1.899347e-11, 1.922433e-11, 1.913439e-11, 
    1.961099e-11, 1.940487e-11, 1.994489e-11, 1.981488e-11, 1.997613e-11, 
    1.989375e-11, 2.003502e-11, 1.990785e-11, 2.012844e-11, 2.017666e-11, 
    2.01437e-11, 2.027047e-11, 1.990082e-11, 2.004231e-11, 1.899243e-11, 
    1.89985e-11, 1.902684e-11, 1.890245e-11, 1.889486e-11, 1.87813e-11, 
    1.888232e-11, 1.892544e-11, 1.903514e-11, 1.91002e-11, 1.916217e-11, 
    1.929882e-11, 1.94521e-11, 1.966762e-11, 1.98233e-11, 1.992805e-11, 
    1.986378e-11, 1.992052e-11, 1.98571e-11, 1.982741e-11, 2.015858e-11, 
    1.997223e-11, 2.025221e-11, 2.023666e-11, 2.010973e-11, 2.023841e-11, 
    1.900278e-11, 1.89678e-11, 1.884665e-11, 1.894142e-11, 1.876896e-11, 
    1.886538e-11, 1.892096e-11, 1.913627e-11, 1.918376e-11, 1.922786e-11, 
    1.931513e-11, 1.942746e-11, 1.962544e-11, 1.979864e-11, 1.995752e-11, 
    1.994586e-11, 1.994996e-11, 1.998555e-11, 1.989747e-11, 2.000003e-11, 
    2.001728e-11, 1.997221e-11, 2.023457e-11, 2.015941e-11, 2.023633e-11, 
    2.018737e-11, 1.897916e-11, 1.903806e-11, 1.900622e-11, 1.906612e-11, 
    1.902391e-11, 1.9212e-11, 1.92686e-11, 1.953473e-11, 1.942525e-11, 
    1.959965e-11, 1.944292e-11, 1.947064e-11, 1.960536e-11, 1.945137e-11, 
    1.978907e-11, 1.955976e-11, 1.998693e-11, 1.975662e-11, 2.000142e-11, 
    1.995683e-11, 2.003068e-11, 2.009696e-11, 2.018052e-11, 2.033524e-11, 
    2.029935e-11, 2.042913e-11, 1.912605e-11, 1.92028e-11, 1.919604e-11, 
    1.927653e-11, 1.933618e-11, 1.946584e-11, 1.967486e-11, 1.959611e-11, 
    1.974081e-11, 1.976994e-11, 1.955014e-11, 1.968493e-11, 1.925427e-11, 
    1.932348e-11, 1.928225e-11, 1.91321e-11, 1.961424e-11, 1.936594e-11, 
    1.982588e-11, 1.969029e-11, 2.00875e-11, 1.988939e-11, 2.027961e-11, 
    2.044779e-11, 2.060679e-11, 2.079355e-11, 1.924476e-11, 1.919253e-11, 
    1.928611e-11, 1.941603e-11, 1.953702e-11, 1.969855e-11, 1.971512e-11, 
    1.974548e-11, 1.982425e-11, 1.989062e-11, 1.975509e-11, 1.990728e-11, 
    1.933956e-11, 1.963588e-11, 1.91728e-11, 1.931158e-11, 1.940836e-11, 
    1.936586e-11, 1.958711e-11, 1.963948e-11, 1.985308e-11, 1.974249e-11, 
    2.040621e-11, 2.011098e-11, 2.093641e-11, 2.070378e-11, 1.91743e-11, 
    1.924458e-11, 1.949036e-11, 1.93732e-11, 1.970936e-11, 1.979262e-11, 
    1.986045e-11, 1.994737e-11, 1.995676e-11, 2.000838e-11, 1.992384e-11, 
    2.000503e-11, 1.969889e-11, 1.983536e-11, 1.946217e-11, 1.955263e-11, 
    1.951098e-11, 1.946537e-11, 1.960636e-11, 1.975722e-11, 1.976044e-11, 
    1.980897e-11, 1.994608e-11, 1.971073e-11, 2.044451e-11, 1.998951e-11, 
    1.932139e-11, 1.945751e-11, 1.947699e-11, 1.942417e-11, 1.978426e-11, 
    1.965335e-11, 2.000712e-11, 1.991114e-11, 2.006853e-11, 1.999023e-11, 
    1.997873e-11, 1.987845e-11, 1.981618e-11, 1.965934e-11, 1.953226e-11, 
    1.943183e-11, 1.945515e-11, 1.956557e-11, 1.976647e-11, 1.995761e-11, 
    1.991565e-11, 2.005654e-11, 1.968487e-11, 1.984023e-11, 1.97801e-11, 
    1.993711e-11, 1.959402e-11, 1.988598e-11, 1.951979e-11, 1.955174e-11, 
    1.965075e-11, 1.98508e-11, 1.989521e-11, 1.99427e-11, 1.991339e-11, 
    1.977158e-11, 1.97484e-11, 1.964834e-11, 1.962077e-11, 1.954478e-11, 
    1.9482e-11, 1.953936e-11, 1.95997e-11, 1.977164e-11, 1.992734e-11, 
    2.009791e-11, 2.013978e-11, 2.03404e-11, 2.0177e-11, 2.044706e-11, 
    2.021734e-11, 2.061595e-11, 1.990297e-11, 2.021059e-11, 1.965526e-11, 
    1.971466e-11, 1.982235e-11, 2.007064e-11, 1.993637e-11, 2.009345e-11, 
    1.97475e-11, 1.956939e-11, 1.952345e-11, 1.943793e-11, 1.952541e-11, 
    1.951828e-11, 1.960219e-11, 1.957521e-11, 1.977736e-11, 1.966862e-11, 
    1.997844e-11, 2.00922e-11, 2.041551e-11, 2.06152e-11, 2.081964e-11, 
    2.091028e-11, 2.093791e-11, 2.094947e-11,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
